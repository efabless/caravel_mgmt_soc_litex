VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mgmt_core_wrapper
  CLASS BLOCK ;
  FOREIGN mgmt_core_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2620.000 BY 800.000 ;
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 134.280 11.000 137.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 549.000 134.280 601.000 137.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 2589.000 134.280 2614.180 137.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 264.280 11.000 267.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 549.000 264.280 601.000 267.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 2589.000 264.280 2614.180 267.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 394.280 11.000 397.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 549.000 394.280 601.000 397.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 2589.000 394.280 2614.180 397.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 524.280 11.000 527.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 549.000 524.280 601.000 527.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 2589.000 524.280 2614.180 527.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 654.280 11.000 657.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 549.000 654.280 601.000 657.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 2589.000 654.280 2614.180 657.480 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 69.280 11.000 72.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 549.000 69.280 601.000 72.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 2589.000 69.280 2614.180 72.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 199.280 11.000 202.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 549.000 199.280 601.000 202.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 2589.000 199.280 2614.180 202.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 329.280 11.000 332.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 549.000 329.280 601.000 332.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 2589.000 329.280 2614.180 332.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 459.280 11.000 462.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 549.000 459.280 601.000 462.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 2589.000 459.280 2614.180 462.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 589.280 11.000 592.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 549.000 589.280 601.000 592.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 2589.000 589.280 2614.180 592.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 719.280 11.000 722.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 549.000 719.280 601.000 722.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 2589.000 719.280 2614.180 722.480 ;
    END
  END VPWR
  PIN core_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1473.930 -2.000 1474.210 4.000 ;
    END
  END core_clk
  PIN core_rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.370 -2.000 491.650 4.000 ;
    END
  END core_rstn
  PIN debug_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 314.200 2622.000 314.800 ;
    END
  END debug_in
  PIN debug_mode
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 321.680 2622.000 322.280 ;
    END
  END debug_mode
  PIN debug_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 329.160 2622.000 329.760 ;
    END
  END debug_oeb
  PIN debug_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 336.640 2622.000 337.240 ;
    END
  END debug_out
  PIN flash_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 706.560 2622.000 707.160 ;
    END
  END flash_clk
  PIN flash_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 699.080 2622.000 699.680 ;
    END
  END flash_csb
  PIN flash_io0_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 714.040 2622.000 714.640 ;
    END
  END flash_io0_di
  PIN flash_io0_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 721.520 2622.000 722.120 ;
    END
  END flash_io0_do
  PIN flash_io0_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 729.000 2622.000 729.600 ;
    END
  END flash_io0_oeb
  PIN flash_io1_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 736.480 2622.000 737.080 ;
    END
  END flash_io1_di
  PIN flash_io1_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 743.280 2622.000 743.880 ;
    END
  END flash_io1_do
  PIN flash_io1_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 750.760 2622.000 751.360 ;
    END
  END flash_io1_oeb
  PIN flash_io2_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 758.240 2622.000 758.840 ;
    END
  END flash_io2_di
  PIN flash_io2_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 765.720 2622.000 766.320 ;
    END
  END flash_io2_do
  PIN flash_io2_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 773.200 2622.000 773.800 ;
    END
  END flash_io2_oeb
  PIN flash_io3_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 780.680 2622.000 781.280 ;
    END
  END flash_io3_di
  PIN flash_io3_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 788.160 2622.000 788.760 ;
    END
  END flash_io3_do
  PIN flash_io3_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 795.640 2622.000 796.240 ;
    END
  END flash_io3_oeb
  PIN gpio_in_pad
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 -2.000 164.130 4.000 ;
    END
  END gpio_in_pad
  PIN gpio_inenb_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.890 -2.000 819.170 4.000 ;
    END
  END gpio_inenb_pad
  PIN gpio_mode0_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1146.410 -2.000 1146.690 4.000 ;
    END
  END gpio_mode0_pad
  PIN gpio_mode1_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1801.450 -2.000 1801.730 4.000 ;
    END
  END gpio_mode1_pad
  PIN gpio_out_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2128.970 -2.000 2129.250 4.000 ;
    END
  END gpio_out_pad
  PIN gpio_outenb_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2456.490 -2.000 2456.770 4.000 ;
    END
  END gpio_outenb_pad
  PIN hk_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 447.480 2622.000 448.080 ;
    END
  END hk_ack_i
  PIN hk_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2617.490 796.000 2617.770 802.000 ;
    END
  END hk_cyc_o
  PIN hk_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 462.440 2622.000 463.040 ;
    END
  END hk_dat_i[0]
  PIN hk_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 536.560 2622.000 537.160 ;
    END
  END hk_dat_i[10]
  PIN hk_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 543.360 2622.000 543.960 ;
    END
  END hk_dat_i[11]
  PIN hk_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 550.840 2622.000 551.440 ;
    END
  END hk_dat_i[12]
  PIN hk_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 558.320 2622.000 558.920 ;
    END
  END hk_dat_i[13]
  PIN hk_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 565.800 2622.000 566.400 ;
    END
  END hk_dat_i[14]
  PIN hk_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 573.280 2622.000 573.880 ;
    END
  END hk_dat_i[15]
  PIN hk_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 580.760 2622.000 581.360 ;
    END
  END hk_dat_i[16]
  PIN hk_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 588.240 2622.000 588.840 ;
    END
  END hk_dat_i[17]
  PIN hk_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 595.720 2622.000 596.320 ;
    END
  END hk_dat_i[18]
  PIN hk_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 603.200 2622.000 603.800 ;
    END
  END hk_dat_i[19]
  PIN hk_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 469.920 2622.000 470.520 ;
    END
  END hk_dat_i[1]
  PIN hk_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 610.000 2622.000 610.600 ;
    END
  END hk_dat_i[20]
  PIN hk_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 617.480 2622.000 618.080 ;
    END
  END hk_dat_i[21]
  PIN hk_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 624.960 2622.000 625.560 ;
    END
  END hk_dat_i[22]
  PIN hk_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 632.440 2622.000 633.040 ;
    END
  END hk_dat_i[23]
  PIN hk_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 639.920 2622.000 640.520 ;
    END
  END hk_dat_i[24]
  PIN hk_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 647.400 2622.000 648.000 ;
    END
  END hk_dat_i[25]
  PIN hk_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 654.880 2622.000 655.480 ;
    END
  END hk_dat_i[26]
  PIN hk_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 662.360 2622.000 662.960 ;
    END
  END hk_dat_i[27]
  PIN hk_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 669.840 2622.000 670.440 ;
    END
  END hk_dat_i[28]
  PIN hk_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 676.640 2622.000 677.240 ;
    END
  END hk_dat_i[29]
  PIN hk_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 476.720 2622.000 477.320 ;
    END
  END hk_dat_i[2]
  PIN hk_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 684.120 2622.000 684.720 ;
    END
  END hk_dat_i[30]
  PIN hk_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 691.600 2622.000 692.200 ;
    END
  END hk_dat_i[31]
  PIN hk_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 484.200 2622.000 484.800 ;
    END
  END hk_dat_i[3]
  PIN hk_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 491.680 2622.000 492.280 ;
    END
  END hk_dat_i[4]
  PIN hk_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 499.160 2622.000 499.760 ;
    END
  END hk_dat_i[5]
  PIN hk_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 506.640 2622.000 507.240 ;
    END
  END hk_dat_i[6]
  PIN hk_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 514.120 2622.000 514.720 ;
    END
  END hk_dat_i[7]
  PIN hk_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 521.600 2622.000 522.200 ;
    END
  END hk_dat_i[8]
  PIN hk_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 529.080 2622.000 529.680 ;
    END
  END hk_dat_i[9]
  PIN hk_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 454.960 2622.000 455.560 ;
    END
  END hk_stb_o
  PIN irq[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2605.070 796.000 2605.350 802.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2609.210 796.000 2609.490 802.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2613.350 796.000 2613.630 802.000 ;
    END
  END irq[2]
  PIN irq[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 365.880 2622.000 366.480 ;
    END
  END irq[3]
  PIN irq[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 358.400 2622.000 359.000 ;
    END
  END irq[4]
  PIN irq[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 350.920 2622.000 351.520 ;
    END
  END irq[5]
  PIN la_iena[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 796.000 2.210 802.000 ;
    END
  END la_iena[0]
  PIN la_iena[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1681.390 796.000 1681.670 802.000 ;
    END
  END la_iena[100]
  PIN la_iena[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1697.950 796.000 1698.230 802.000 ;
    END
  END la_iena[101]
  PIN la_iena[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1714.970 796.000 1715.250 802.000 ;
    END
  END la_iena[102]
  PIN la_iena[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1731.530 796.000 1731.810 802.000 ;
    END
  END la_iena[103]
  PIN la_iena[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1748.550 796.000 1748.830 802.000 ;
    END
  END la_iena[104]
  PIN la_iena[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1765.110 796.000 1765.390 802.000 ;
    END
  END la_iena[105]
  PIN la_iena[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1782.130 796.000 1782.410 802.000 ;
    END
  END la_iena[106]
  PIN la_iena[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1798.690 796.000 1798.970 802.000 ;
    END
  END la_iena[107]
  PIN la_iena[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1815.710 796.000 1815.990 802.000 ;
    END
  END la_iena[108]
  PIN la_iena[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1832.270 796.000 1832.550 802.000 ;
    END
  END la_iena[109]
  PIN la_iena[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 796.000 170.110 802.000 ;
    END
  END la_iena[10]
  PIN la_iena[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1849.290 796.000 1849.570 802.000 ;
    END
  END la_iena[110]
  PIN la_iena[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1865.850 796.000 1866.130 802.000 ;
    END
  END la_iena[111]
  PIN la_iena[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1882.870 796.000 1883.150 802.000 ;
    END
  END la_iena[112]
  PIN la_iena[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1899.430 796.000 1899.710 802.000 ;
    END
  END la_iena[113]
  PIN la_iena[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1916.450 796.000 1916.730 802.000 ;
    END
  END la_iena[114]
  PIN la_iena[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1933.010 796.000 1933.290 802.000 ;
    END
  END la_iena[115]
  PIN la_iena[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1950.030 796.000 1950.310 802.000 ;
    END
  END la_iena[116]
  PIN la_iena[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1967.050 796.000 1967.330 802.000 ;
    END
  END la_iena[117]
  PIN la_iena[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1983.610 796.000 1983.890 802.000 ;
    END
  END la_iena[118]
  PIN la_iena[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2000.630 796.000 2000.910 802.000 ;
    END
  END la_iena[119]
  PIN la_iena[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 796.000 186.670 802.000 ;
    END
  END la_iena[11]
  PIN la_iena[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2017.190 796.000 2017.470 802.000 ;
    END
  END la_iena[120]
  PIN la_iena[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2034.210 796.000 2034.490 802.000 ;
    END
  END la_iena[121]
  PIN la_iena[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2050.770 796.000 2051.050 802.000 ;
    END
  END la_iena[122]
  PIN la_iena[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2067.790 796.000 2068.070 802.000 ;
    END
  END la_iena[123]
  PIN la_iena[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2084.350 796.000 2084.630 802.000 ;
    END
  END la_iena[124]
  PIN la_iena[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2101.370 796.000 2101.650 802.000 ;
    END
  END la_iena[125]
  PIN la_iena[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2117.930 796.000 2118.210 802.000 ;
    END
  END la_iena[126]
  PIN la_iena[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2134.950 796.000 2135.230 802.000 ;
    END
  END la_iena[127]
  PIN la_iena[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 796.000 203.690 802.000 ;
    END
  END la_iena[12]
  PIN la_iena[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 796.000 220.250 802.000 ;
    END
  END la_iena[13]
  PIN la_iena[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 796.000 237.270 802.000 ;
    END
  END la_iena[14]
  PIN la_iena[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 796.000 253.830 802.000 ;
    END
  END la_iena[15]
  PIN la_iena[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 796.000 270.850 802.000 ;
    END
  END la_iena[16]
  PIN la_iena[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 796.000 287.410 802.000 ;
    END
  END la_iena[17]
  PIN la_iena[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.150 796.000 304.430 802.000 ;
    END
  END la_iena[18]
  PIN la_iena[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.710 796.000 320.990 802.000 ;
    END
  END la_iena[19]
  PIN la_iena[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 796.000 18.770 802.000 ;
    END
  END la_iena[1]
  PIN la_iena[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 796.000 338.010 802.000 ;
    END
  END la_iena[20]
  PIN la_iena[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 796.000 354.570 802.000 ;
    END
  END la_iena[21]
  PIN la_iena[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 796.000 371.590 802.000 ;
    END
  END la_iena[22]
  PIN la_iena[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 796.000 388.150 802.000 ;
    END
  END la_iena[23]
  PIN la_iena[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 796.000 405.170 802.000 ;
    END
  END la_iena[24]
  PIN la_iena[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.450 796.000 421.730 802.000 ;
    END
  END la_iena[25]
  PIN la_iena[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.470 796.000 438.750 802.000 ;
    END
  END la_iena[26]
  PIN la_iena[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.030 796.000 455.310 802.000 ;
    END
  END la_iena[27]
  PIN la_iena[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.050 796.000 472.330 802.000 ;
    END
  END la_iena[28]
  PIN la_iena[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 796.000 488.890 802.000 ;
    END
  END la_iena[29]
  PIN la_iena[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 796.000 35.790 802.000 ;
    END
  END la_iena[2]
  PIN la_iena[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 796.000 505.910 802.000 ;
    END
  END la_iena[30]
  PIN la_iena[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 796.000 522.470 802.000 ;
    END
  END la_iena[31]
  PIN la_iena[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 796.000 539.490 802.000 ;
    END
  END la_iena[32]
  PIN la_iena[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.770 796.000 556.050 802.000 ;
    END
  END la_iena[33]
  PIN la_iena[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.790 796.000 573.070 802.000 ;
    END
  END la_iena[34]
  PIN la_iena[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 796.000 589.630 802.000 ;
    END
  END la_iena[35]
  PIN la_iena[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.370 796.000 606.650 802.000 ;
    END
  END la_iena[36]
  PIN la_iena[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.930 796.000 623.210 802.000 ;
    END
  END la_iena[37]
  PIN la_iena[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.950 796.000 640.230 802.000 ;
    END
  END la_iena[38]
  PIN la_iena[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 796.000 657.250 802.000 ;
    END
  END la_iena[39]
  PIN la_iena[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 796.000 52.350 802.000 ;
    END
  END la_iena[3]
  PIN la_iena[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.530 796.000 673.810 802.000 ;
    END
  END la_iena[40]
  PIN la_iena[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.550 796.000 690.830 802.000 ;
    END
  END la_iena[41]
  PIN la_iena[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.110 796.000 707.390 802.000 ;
    END
  END la_iena[42]
  PIN la_iena[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.130 796.000 724.410 802.000 ;
    END
  END la_iena[43]
  PIN la_iena[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 796.000 740.970 802.000 ;
    END
  END la_iena[44]
  PIN la_iena[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.710 796.000 757.990 802.000 ;
    END
  END la_iena[45]
  PIN la_iena[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.270 796.000 774.550 802.000 ;
    END
  END la_iena[46]
  PIN la_iena[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.290 796.000 791.570 802.000 ;
    END
  END la_iena[47]
  PIN la_iena[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.850 796.000 808.130 802.000 ;
    END
  END la_iena[48]
  PIN la_iena[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.870 796.000 825.150 802.000 ;
    END
  END la_iena[49]
  PIN la_iena[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 796.000 69.370 802.000 ;
    END
  END la_iena[4]
  PIN la_iena[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.430 796.000 841.710 802.000 ;
    END
  END la_iena[50]
  PIN la_iena[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.450 796.000 858.730 802.000 ;
    END
  END la_iena[51]
  PIN la_iena[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.010 796.000 875.290 802.000 ;
    END
  END la_iena[52]
  PIN la_iena[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.030 796.000 892.310 802.000 ;
    END
  END la_iena[53]
  PIN la_iena[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.590 796.000 908.870 802.000 ;
    END
  END la_iena[54]
  PIN la_iena[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 925.610 796.000 925.890 802.000 ;
    END
  END la_iena[55]
  PIN la_iena[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.170 796.000 942.450 802.000 ;
    END
  END la_iena[56]
  PIN la_iena[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.190 796.000 959.470 802.000 ;
    END
  END la_iena[57]
  PIN la_iena[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.750 796.000 976.030 802.000 ;
    END
  END la_iena[58]
  PIN la_iena[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 992.770 796.000 993.050 802.000 ;
    END
  END la_iena[59]
  PIN la_iena[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 796.000 85.930 802.000 ;
    END
  END la_iena[5]
  PIN la_iena[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.330 796.000 1009.610 802.000 ;
    END
  END la_iena[60]
  PIN la_iena[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1026.350 796.000 1026.630 802.000 ;
    END
  END la_iena[61]
  PIN la_iena[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.910 796.000 1043.190 802.000 ;
    END
  END la_iena[62]
  PIN la_iena[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.930 796.000 1060.210 802.000 ;
    END
  END la_iena[63]
  PIN la_iena[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.490 796.000 1076.770 802.000 ;
    END
  END la_iena[64]
  PIN la_iena[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1093.510 796.000 1093.790 802.000 ;
    END
  END la_iena[65]
  PIN la_iena[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.070 796.000 1110.350 802.000 ;
    END
  END la_iena[66]
  PIN la_iena[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.090 796.000 1127.370 802.000 ;
    END
  END la_iena[67]
  PIN la_iena[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.650 796.000 1143.930 802.000 ;
    END
  END la_iena[68]
  PIN la_iena[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.670 796.000 1160.950 802.000 ;
    END
  END la_iena[69]
  PIN la_iena[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 796.000 102.950 802.000 ;
    END
  END la_iena[6]
  PIN la_iena[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1177.230 796.000 1177.510 802.000 ;
    END
  END la_iena[70]
  PIN la_iena[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.250 796.000 1194.530 802.000 ;
    END
  END la_iena[71]
  PIN la_iena[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1210.810 796.000 1211.090 802.000 ;
    END
  END la_iena[72]
  PIN la_iena[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.830 796.000 1228.110 802.000 ;
    END
  END la_iena[73]
  PIN la_iena[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1244.390 796.000 1244.670 802.000 ;
    END
  END la_iena[74]
  PIN la_iena[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1261.410 796.000 1261.690 802.000 ;
    END
  END la_iena[75]
  PIN la_iena[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1277.970 796.000 1278.250 802.000 ;
    END
  END la_iena[76]
  PIN la_iena[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.990 796.000 1295.270 802.000 ;
    END
  END la_iena[77]
  PIN la_iena[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1312.010 796.000 1312.290 802.000 ;
    END
  END la_iena[78]
  PIN la_iena[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1328.570 796.000 1328.850 802.000 ;
    END
  END la_iena[79]
  PIN la_iena[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 796.000 119.510 802.000 ;
    END
  END la_iena[7]
  PIN la_iena[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1345.590 796.000 1345.870 802.000 ;
    END
  END la_iena[80]
  PIN la_iena[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.150 796.000 1362.430 802.000 ;
    END
  END la_iena[81]
  PIN la_iena[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1379.170 796.000 1379.450 802.000 ;
    END
  END la_iena[82]
  PIN la_iena[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1395.730 796.000 1396.010 802.000 ;
    END
  END la_iena[83]
  PIN la_iena[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1412.750 796.000 1413.030 802.000 ;
    END
  END la_iena[84]
  PIN la_iena[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.310 796.000 1429.590 802.000 ;
    END
  END la_iena[85]
  PIN la_iena[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1446.330 796.000 1446.610 802.000 ;
    END
  END la_iena[86]
  PIN la_iena[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.890 796.000 1463.170 802.000 ;
    END
  END la_iena[87]
  PIN la_iena[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1479.910 796.000 1480.190 802.000 ;
    END
  END la_iena[88]
  PIN la_iena[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1496.470 796.000 1496.750 802.000 ;
    END
  END la_iena[89]
  PIN la_iena[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 796.000 136.530 802.000 ;
    END
  END la_iena[8]
  PIN la_iena[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.490 796.000 1513.770 802.000 ;
    END
  END la_iena[90]
  PIN la_iena[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1530.050 796.000 1530.330 802.000 ;
    END
  END la_iena[91]
  PIN la_iena[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1547.070 796.000 1547.350 802.000 ;
    END
  END la_iena[92]
  PIN la_iena[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1563.630 796.000 1563.910 802.000 ;
    END
  END la_iena[93]
  PIN la_iena[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.650 796.000 1580.930 802.000 ;
    END
  END la_iena[94]
  PIN la_iena[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.210 796.000 1597.490 802.000 ;
    END
  END la_iena[95]
  PIN la_iena[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1614.230 796.000 1614.510 802.000 ;
    END
  END la_iena[96]
  PIN la_iena[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1630.790 796.000 1631.070 802.000 ;
    END
  END la_iena[97]
  PIN la_iena[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1647.810 796.000 1648.090 802.000 ;
    END
  END la_iena[98]
  PIN la_iena[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1664.370 796.000 1664.650 802.000 ;
    END
  END la_iena[99]
  PIN la_iena[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 796.000 153.090 802.000 ;
    END
  END la_iena[9]
  PIN la_input[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 796.000 6.350 802.000 ;
    END
  END la_input[0]
  PIN la_input[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1685.530 796.000 1685.810 802.000 ;
    END
  END la_input[100]
  PIN la_input[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1702.090 796.000 1702.370 802.000 ;
    END
  END la_input[101]
  PIN la_input[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1719.110 796.000 1719.390 802.000 ;
    END
  END la_input[102]
  PIN la_input[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1735.670 796.000 1735.950 802.000 ;
    END
  END la_input[103]
  PIN la_input[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1752.690 796.000 1752.970 802.000 ;
    END
  END la_input[104]
  PIN la_input[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1769.250 796.000 1769.530 802.000 ;
    END
  END la_input[105]
  PIN la_input[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1786.270 796.000 1786.550 802.000 ;
    END
  END la_input[106]
  PIN la_input[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1803.290 796.000 1803.570 802.000 ;
    END
  END la_input[107]
  PIN la_input[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1819.850 796.000 1820.130 802.000 ;
    END
  END la_input[108]
  PIN la_input[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1836.870 796.000 1837.150 802.000 ;
    END
  END la_input[109]
  PIN la_input[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 796.000 174.250 802.000 ;
    END
  END la_input[10]
  PIN la_input[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1853.430 796.000 1853.710 802.000 ;
    END
  END la_input[110]
  PIN la_input[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1870.450 796.000 1870.730 802.000 ;
    END
  END la_input[111]
  PIN la_input[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1887.010 796.000 1887.290 802.000 ;
    END
  END la_input[112]
  PIN la_input[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1904.030 796.000 1904.310 802.000 ;
    END
  END la_input[113]
  PIN la_input[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1920.590 796.000 1920.870 802.000 ;
    END
  END la_input[114]
  PIN la_input[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1937.610 796.000 1937.890 802.000 ;
    END
  END la_input[115]
  PIN la_input[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1954.170 796.000 1954.450 802.000 ;
    END
  END la_input[116]
  PIN la_input[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1971.190 796.000 1971.470 802.000 ;
    END
  END la_input[117]
  PIN la_input[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1987.750 796.000 1988.030 802.000 ;
    END
  END la_input[118]
  PIN la_input[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2004.770 796.000 2005.050 802.000 ;
    END
  END la_input[119]
  PIN la_input[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 796.000 190.810 802.000 ;
    END
  END la_input[11]
  PIN la_input[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2021.330 796.000 2021.610 802.000 ;
    END
  END la_input[120]
  PIN la_input[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2038.350 796.000 2038.630 802.000 ;
    END
  END la_input[121]
  PIN la_input[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2054.910 796.000 2055.190 802.000 ;
    END
  END la_input[122]
  PIN la_input[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2071.930 796.000 2072.210 802.000 ;
    END
  END la_input[123]
  PIN la_input[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2088.490 796.000 2088.770 802.000 ;
    END
  END la_input[124]
  PIN la_input[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2105.510 796.000 2105.790 802.000 ;
    END
  END la_input[125]
  PIN la_input[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2122.070 796.000 2122.350 802.000 ;
    END
  END la_input[126]
  PIN la_input[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2139.090 796.000 2139.370 802.000 ;
    END
  END la_input[127]
  PIN la_input[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 796.000 207.830 802.000 ;
    END
  END la_input[12]
  PIN la_input[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 796.000 224.390 802.000 ;
    END
  END la_input[13]
  PIN la_input[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.130 796.000 241.410 802.000 ;
    END
  END la_input[14]
  PIN la_input[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 796.000 257.970 802.000 ;
    END
  END la_input[15]
  PIN la_input[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 796.000 274.990 802.000 ;
    END
  END la_input[16]
  PIN la_input[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 796.000 291.550 802.000 ;
    END
  END la_input[17]
  PIN la_input[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 796.000 308.570 802.000 ;
    END
  END la_input[18]
  PIN la_input[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 796.000 325.130 802.000 ;
    END
  END la_input[19]
  PIN la_input[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 796.000 22.910 802.000 ;
    END
  END la_input[1]
  PIN la_input[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 796.000 342.150 802.000 ;
    END
  END la_input[20]
  PIN la_input[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 796.000 358.710 802.000 ;
    END
  END la_input[21]
  PIN la_input[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.450 796.000 375.730 802.000 ;
    END
  END la_input[22]
  PIN la_input[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 796.000 392.290 802.000 ;
    END
  END la_input[23]
  PIN la_input[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 796.000 409.310 802.000 ;
    END
  END la_input[24]
  PIN la_input[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 796.000 425.870 802.000 ;
    END
  END la_input[25]
  PIN la_input[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.610 796.000 442.890 802.000 ;
    END
  END la_input[26]
  PIN la_input[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.170 796.000 459.450 802.000 ;
    END
  END la_input[27]
  PIN la_input[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.190 796.000 476.470 802.000 ;
    END
  END la_input[28]
  PIN la_input[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.210 796.000 493.490 802.000 ;
    END
  END la_input[29]
  PIN la_input[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 796.000 39.930 802.000 ;
    END
  END la_input[2]
  PIN la_input[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 796.000 510.050 802.000 ;
    END
  END la_input[30]
  PIN la_input[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.790 796.000 527.070 802.000 ;
    END
  END la_input[31]
  PIN la_input[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.350 796.000 543.630 802.000 ;
    END
  END la_input[32]
  PIN la_input[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 796.000 560.650 802.000 ;
    END
  END la_input[33]
  PIN la_input[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.930 796.000 577.210 802.000 ;
    END
  END la_input[34]
  PIN la_input[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.950 796.000 594.230 802.000 ;
    END
  END la_input[35]
  PIN la_input[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.510 796.000 610.790 802.000 ;
    END
  END la_input[36]
  PIN la_input[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.530 796.000 627.810 802.000 ;
    END
  END la_input[37]
  PIN la_input[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 796.000 644.370 802.000 ;
    END
  END la_input[38]
  PIN la_input[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.110 796.000 661.390 802.000 ;
    END
  END la_input[39]
  PIN la_input[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 796.000 56.490 802.000 ;
    END
  END la_input[3]
  PIN la_input[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.670 796.000 677.950 802.000 ;
    END
  END la_input[40]
  PIN la_input[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.690 796.000 694.970 802.000 ;
    END
  END la_input[41]
  PIN la_input[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.250 796.000 711.530 802.000 ;
    END
  END la_input[42]
  PIN la_input[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.270 796.000 728.550 802.000 ;
    END
  END la_input[43]
  PIN la_input[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.830 796.000 745.110 802.000 ;
    END
  END la_input[44]
  PIN la_input[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.850 796.000 762.130 802.000 ;
    END
  END la_input[45]
  PIN la_input[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.410 796.000 778.690 802.000 ;
    END
  END la_input[46]
  PIN la_input[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.430 796.000 795.710 802.000 ;
    END
  END la_input[47]
  PIN la_input[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.990 796.000 812.270 802.000 ;
    END
  END la_input[48]
  PIN la_input[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.010 796.000 829.290 802.000 ;
    END
  END la_input[49]
  PIN la_input[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 796.000 73.510 802.000 ;
    END
  END la_input[4]
  PIN la_input[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.570 796.000 845.850 802.000 ;
    END
  END la_input[50]
  PIN la_input[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.590 796.000 862.870 802.000 ;
    END
  END la_input[51]
  PIN la_input[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 796.000 879.430 802.000 ;
    END
  END la_input[52]
  PIN la_input[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 896.170 796.000 896.450 802.000 ;
    END
  END la_input[53]
  PIN la_input[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.730 796.000 913.010 802.000 ;
    END
  END la_input[54]
  PIN la_input[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.750 796.000 930.030 802.000 ;
    END
  END la_input[55]
  PIN la_input[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.310 796.000 946.590 802.000 ;
    END
  END la_input[56]
  PIN la_input[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.330 796.000 963.610 802.000 ;
    END
  END la_input[57]
  PIN la_input[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.890 796.000 980.170 802.000 ;
    END
  END la_input[58]
  PIN la_input[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 996.910 796.000 997.190 802.000 ;
    END
  END la_input[59]
  PIN la_input[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 796.000 90.070 802.000 ;
    END
  END la_input[5]
  PIN la_input[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.470 796.000 1013.750 802.000 ;
    END
  END la_input[60]
  PIN la_input[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.490 796.000 1030.770 802.000 ;
    END
  END la_input[61]
  PIN la_input[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.050 796.000 1047.330 802.000 ;
    END
  END la_input[62]
  PIN la_input[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.070 796.000 1064.350 802.000 ;
    END
  END la_input[63]
  PIN la_input[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1080.630 796.000 1080.910 802.000 ;
    END
  END la_input[64]
  PIN la_input[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1097.650 796.000 1097.930 802.000 ;
    END
  END la_input[65]
  PIN la_input[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.210 796.000 1114.490 802.000 ;
    END
  END la_input[66]
  PIN la_input[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.230 796.000 1131.510 802.000 ;
    END
  END la_input[67]
  PIN la_input[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1148.250 796.000 1148.530 802.000 ;
    END
  END la_input[68]
  PIN la_input[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1164.810 796.000 1165.090 802.000 ;
    END
  END la_input[69]
  PIN la_input[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 796.000 107.090 802.000 ;
    END
  END la_input[6]
  PIN la_input[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1181.830 796.000 1182.110 802.000 ;
    END
  END la_input[70]
  PIN la_input[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1198.390 796.000 1198.670 802.000 ;
    END
  END la_input[71]
  PIN la_input[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1215.410 796.000 1215.690 802.000 ;
    END
  END la_input[72]
  PIN la_input[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.970 796.000 1232.250 802.000 ;
    END
  END la_input[73]
  PIN la_input[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1248.990 796.000 1249.270 802.000 ;
    END
  END la_input[74]
  PIN la_input[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1265.550 796.000 1265.830 802.000 ;
    END
  END la_input[75]
  PIN la_input[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1282.570 796.000 1282.850 802.000 ;
    END
  END la_input[76]
  PIN la_input[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1299.130 796.000 1299.410 802.000 ;
    END
  END la_input[77]
  PIN la_input[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1316.150 796.000 1316.430 802.000 ;
    END
  END la_input[78]
  PIN la_input[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.710 796.000 1332.990 802.000 ;
    END
  END la_input[79]
  PIN la_input[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 796.000 123.650 802.000 ;
    END
  END la_input[7]
  PIN la_input[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.730 796.000 1350.010 802.000 ;
    END
  END la_input[80]
  PIN la_input[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1366.290 796.000 1366.570 802.000 ;
    END
  END la_input[81]
  PIN la_input[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1383.310 796.000 1383.590 802.000 ;
    END
  END la_input[82]
  PIN la_input[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1399.870 796.000 1400.150 802.000 ;
    END
  END la_input[83]
  PIN la_input[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1416.890 796.000 1417.170 802.000 ;
    END
  END la_input[84]
  PIN la_input[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1433.450 796.000 1433.730 802.000 ;
    END
  END la_input[85]
  PIN la_input[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1450.470 796.000 1450.750 802.000 ;
    END
  END la_input[86]
  PIN la_input[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1467.030 796.000 1467.310 802.000 ;
    END
  END la_input[87]
  PIN la_input[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.050 796.000 1484.330 802.000 ;
    END
  END la_input[88]
  PIN la_input[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.610 796.000 1500.890 802.000 ;
    END
  END la_input[89]
  PIN la_input[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 796.000 140.670 802.000 ;
    END
  END la_input[8]
  PIN la_input[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1517.630 796.000 1517.910 802.000 ;
    END
  END la_input[90]
  PIN la_input[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1534.190 796.000 1534.470 802.000 ;
    END
  END la_input[91]
  PIN la_input[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1551.210 796.000 1551.490 802.000 ;
    END
  END la_input[92]
  PIN la_input[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1567.770 796.000 1568.050 802.000 ;
    END
  END la_input[93]
  PIN la_input[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.790 796.000 1585.070 802.000 ;
    END
  END la_input[94]
  PIN la_input[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1601.350 796.000 1601.630 802.000 ;
    END
  END la_input[95]
  PIN la_input[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1618.370 796.000 1618.650 802.000 ;
    END
  END la_input[96]
  PIN la_input[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1634.930 796.000 1635.210 802.000 ;
    END
  END la_input[97]
  PIN la_input[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.950 796.000 1652.230 802.000 ;
    END
  END la_input[98]
  PIN la_input[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1668.510 796.000 1668.790 802.000 ;
    END
  END la_input[99]
  PIN la_input[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 796.000 157.230 802.000 ;
    END
  END la_input[9]
  PIN la_oenb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 796.000 10.490 802.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1689.670 796.000 1689.950 802.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1706.690 796.000 1706.970 802.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1723.250 796.000 1723.530 802.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1740.270 796.000 1740.550 802.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1756.830 796.000 1757.110 802.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1773.850 796.000 1774.130 802.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1790.410 796.000 1790.690 802.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1807.430 796.000 1807.710 802.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1823.990 796.000 1824.270 802.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1841.010 796.000 1841.290 802.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 796.000 178.390 802.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1857.570 796.000 1857.850 802.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1874.590 796.000 1874.870 802.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1891.150 796.000 1891.430 802.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1908.170 796.000 1908.450 802.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1924.730 796.000 1925.010 802.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.750 796.000 1942.030 802.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1958.310 796.000 1958.590 802.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1975.330 796.000 1975.610 802.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1991.890 796.000 1992.170 802.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2008.910 796.000 2009.190 802.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 796.000 194.950 802.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2025.470 796.000 2025.750 802.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2042.490 796.000 2042.770 802.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2059.050 796.000 2059.330 802.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2076.070 796.000 2076.350 802.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2092.630 796.000 2092.910 802.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2109.650 796.000 2109.930 802.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2126.210 796.000 2126.490 802.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2143.230 796.000 2143.510 802.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 796.000 211.970 802.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 796.000 228.530 802.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 796.000 245.550 802.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 796.000 262.110 802.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 796.000 279.130 802.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 796.000 295.690 802.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 796.000 312.710 802.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.450 796.000 329.730 802.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 796.000 27.050 802.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.010 796.000 346.290 802.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.030 796.000 363.310 802.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 796.000 379.870 802.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.610 796.000 396.890 802.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.170 796.000 413.450 802.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 796.000 430.470 802.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.750 796.000 447.030 802.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 796.000 464.050 802.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.330 796.000 480.610 802.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.350 796.000 497.630 802.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 796.000 44.070 802.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.910 796.000 514.190 802.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.930 796.000 531.210 802.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 796.000 547.770 802.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.510 796.000 564.790 802.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.070 796.000 581.350 802.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.090 796.000 598.370 802.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.650 796.000 614.930 802.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.670 796.000 631.950 802.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.230 796.000 648.510 802.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.250 796.000 665.530 802.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 796.000 60.630 802.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.810 796.000 682.090 802.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.830 796.000 699.110 802.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.390 796.000 715.670 802.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.410 796.000 732.690 802.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.970 796.000 749.250 802.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.990 796.000 766.270 802.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 796.000 782.830 802.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.570 796.000 799.850 802.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.130 796.000 816.410 802.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.150 796.000 833.430 802.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 796.000 77.650 802.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.710 796.000 849.990 802.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.730 796.000 867.010 802.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.290 796.000 883.570 802.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.310 796.000 900.590 802.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.870 796.000 917.150 802.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.890 796.000 934.170 802.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 950.450 796.000 950.730 802.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.470 796.000 967.750 802.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.490 796.000 984.770 802.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.050 796.000 1001.330 802.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 796.000 94.210 802.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.070 796.000 1018.350 802.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1034.630 796.000 1034.910 802.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.650 796.000 1051.930 802.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1068.210 796.000 1068.490 802.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.230 796.000 1085.510 802.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1101.790 796.000 1102.070 802.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1118.810 796.000 1119.090 802.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1135.370 796.000 1135.650 802.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.390 796.000 1152.670 802.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.950 796.000 1169.230 802.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 796.000 111.230 802.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.970 796.000 1186.250 802.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.530 796.000 1202.810 802.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1219.550 796.000 1219.830 802.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1236.110 796.000 1236.390 802.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1253.130 796.000 1253.410 802.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1269.690 796.000 1269.970 802.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1286.710 796.000 1286.990 802.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1303.270 796.000 1303.550 802.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.290 796.000 1320.570 802.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1336.850 796.000 1337.130 802.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 796.000 127.790 802.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1353.870 796.000 1354.150 802.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1370.430 796.000 1370.710 802.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1387.450 796.000 1387.730 802.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1404.010 796.000 1404.290 802.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.030 796.000 1421.310 802.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1437.590 796.000 1437.870 802.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1454.610 796.000 1454.890 802.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.170 796.000 1471.450 802.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1488.190 796.000 1488.470 802.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1504.750 796.000 1505.030 802.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 796.000 144.810 802.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.770 796.000 1522.050 802.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1538.330 796.000 1538.610 802.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1555.350 796.000 1555.630 802.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1571.910 796.000 1572.190 802.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1588.930 796.000 1589.210 802.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1605.490 796.000 1605.770 802.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1622.510 796.000 1622.790 802.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.530 796.000 1639.810 802.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1656.090 796.000 1656.370 802.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1673.110 796.000 1673.390 802.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 796.000 161.370 802.000 ;
    END
  END la_oenb[9]
  PIN la_output[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 796.000 14.630 802.000 ;
    END
  END la_output[0]
  PIN la_output[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.810 796.000 1694.090 802.000 ;
    END
  END la_output[100]
  PIN la_output[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1710.830 796.000 1711.110 802.000 ;
    END
  END la_output[101]
  PIN la_output[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1727.390 796.000 1727.670 802.000 ;
    END
  END la_output[102]
  PIN la_output[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1744.410 796.000 1744.690 802.000 ;
    END
  END la_output[103]
  PIN la_output[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1760.970 796.000 1761.250 802.000 ;
    END
  END la_output[104]
  PIN la_output[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1777.990 796.000 1778.270 802.000 ;
    END
  END la_output[105]
  PIN la_output[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1794.550 796.000 1794.830 802.000 ;
    END
  END la_output[106]
  PIN la_output[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1811.570 796.000 1811.850 802.000 ;
    END
  END la_output[107]
  PIN la_output[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1828.130 796.000 1828.410 802.000 ;
    END
  END la_output[108]
  PIN la_output[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1845.150 796.000 1845.430 802.000 ;
    END
  END la_output[109]
  PIN la_output[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 796.000 182.530 802.000 ;
    END
  END la_output[10]
  PIN la_output[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1861.710 796.000 1861.990 802.000 ;
    END
  END la_output[110]
  PIN la_output[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1878.730 796.000 1879.010 802.000 ;
    END
  END la_output[111]
  PIN la_output[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1895.290 796.000 1895.570 802.000 ;
    END
  END la_output[112]
  PIN la_output[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1912.310 796.000 1912.590 802.000 ;
    END
  END la_output[113]
  PIN la_output[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1928.870 796.000 1929.150 802.000 ;
    END
  END la_output[114]
  PIN la_output[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1945.890 796.000 1946.170 802.000 ;
    END
  END la_output[115]
  PIN la_output[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1962.450 796.000 1962.730 802.000 ;
    END
  END la_output[116]
  PIN la_output[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1979.470 796.000 1979.750 802.000 ;
    END
  END la_output[117]
  PIN la_output[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1996.030 796.000 1996.310 802.000 ;
    END
  END la_output[118]
  PIN la_output[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2013.050 796.000 2013.330 802.000 ;
    END
  END la_output[119]
  PIN la_output[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.270 796.000 199.550 802.000 ;
    END
  END la_output[11]
  PIN la_output[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2029.610 796.000 2029.890 802.000 ;
    END
  END la_output[120]
  PIN la_output[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2046.630 796.000 2046.910 802.000 ;
    END
  END la_output[121]
  PIN la_output[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2063.190 796.000 2063.470 802.000 ;
    END
  END la_output[122]
  PIN la_output[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2080.210 796.000 2080.490 802.000 ;
    END
  END la_output[123]
  PIN la_output[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2096.770 796.000 2097.050 802.000 ;
    END
  END la_output[124]
  PIN la_output[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2113.790 796.000 2114.070 802.000 ;
    END
  END la_output[125]
  PIN la_output[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2130.810 796.000 2131.090 802.000 ;
    END
  END la_output[126]
  PIN la_output[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2147.370 796.000 2147.650 802.000 ;
    END
  END la_output[127]
  PIN la_output[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 796.000 216.110 802.000 ;
    END
  END la_output[12]
  PIN la_output[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 796.000 233.130 802.000 ;
    END
  END la_output[13]
  PIN la_output[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 796.000 249.690 802.000 ;
    END
  END la_output[14]
  PIN la_output[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 796.000 266.710 802.000 ;
    END
  END la_output[15]
  PIN la_output[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 796.000 283.270 802.000 ;
    END
  END la_output[16]
  PIN la_output[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 796.000 300.290 802.000 ;
    END
  END la_output[17]
  PIN la_output[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 796.000 316.850 802.000 ;
    END
  END la_output[18]
  PIN la_output[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 796.000 333.870 802.000 ;
    END
  END la_output[19]
  PIN la_output[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 796.000 31.190 802.000 ;
    END
  END la_output[1]
  PIN la_output[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 796.000 350.430 802.000 ;
    END
  END la_output[20]
  PIN la_output[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 796.000 367.450 802.000 ;
    END
  END la_output[21]
  PIN la_output[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.730 796.000 384.010 802.000 ;
    END
  END la_output[22]
  PIN la_output[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.750 796.000 401.030 802.000 ;
    END
  END la_output[23]
  PIN la_output[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.310 796.000 417.590 802.000 ;
    END
  END la_output[24]
  PIN la_output[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.330 796.000 434.610 802.000 ;
    END
  END la_output[25]
  PIN la_output[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 796.000 451.170 802.000 ;
    END
  END la_output[26]
  PIN la_output[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.910 796.000 468.190 802.000 ;
    END
  END la_output[27]
  PIN la_output[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.470 796.000 484.750 802.000 ;
    END
  END la_output[28]
  PIN la_output[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.490 796.000 501.770 802.000 ;
    END
  END la_output[29]
  PIN la_output[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 796.000 48.210 802.000 ;
    END
  END la_output[2]
  PIN la_output[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.050 796.000 518.330 802.000 ;
    END
  END la_output[30]
  PIN la_output[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.070 796.000 535.350 802.000 ;
    END
  END la_output[31]
  PIN la_output[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.630 796.000 551.910 802.000 ;
    END
  END la_output[32]
  PIN la_output[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.650 796.000 568.930 802.000 ;
    END
  END la_output[33]
  PIN la_output[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 796.000 585.490 802.000 ;
    END
  END la_output[34]
  PIN la_output[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 796.000 602.510 802.000 ;
    END
  END la_output[35]
  PIN la_output[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.790 796.000 619.070 802.000 ;
    END
  END la_output[36]
  PIN la_output[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.810 796.000 636.090 802.000 ;
    END
  END la_output[37]
  PIN la_output[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.370 796.000 652.650 802.000 ;
    END
  END la_output[38]
  PIN la_output[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.390 796.000 669.670 802.000 ;
    END
  END la_output[39]
  PIN la_output[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 796.000 64.770 802.000 ;
    END
  END la_output[3]
  PIN la_output[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 796.000 686.230 802.000 ;
    END
  END la_output[40]
  PIN la_output[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.970 796.000 703.250 802.000 ;
    END
  END la_output[41]
  PIN la_output[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.530 796.000 719.810 802.000 ;
    END
  END la_output[42]
  PIN la_output[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.550 796.000 736.830 802.000 ;
    END
  END la_output[43]
  PIN la_output[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.110 796.000 753.390 802.000 ;
    END
  END la_output[44]
  PIN la_output[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.130 796.000 770.410 802.000 ;
    END
  END la_output[45]
  PIN la_output[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.690 796.000 786.970 802.000 ;
    END
  END la_output[46]
  PIN la_output[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.710 796.000 803.990 802.000 ;
    END
  END la_output[47]
  PIN la_output[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.730 796.000 821.010 802.000 ;
    END
  END la_output[48]
  PIN la_output[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 796.000 837.570 802.000 ;
    END
  END la_output[49]
  PIN la_output[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 796.000 81.790 802.000 ;
    END
  END la_output[4]
  PIN la_output[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.310 796.000 854.590 802.000 ;
    END
  END la_output[50]
  PIN la_output[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.870 796.000 871.150 802.000 ;
    END
  END la_output[51]
  PIN la_output[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.890 796.000 888.170 802.000 ;
    END
  END la_output[52]
  PIN la_output[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.450 796.000 904.730 802.000 ;
    END
  END la_output[53]
  PIN la_output[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.470 796.000 921.750 802.000 ;
    END
  END la_output[54]
  PIN la_output[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.030 796.000 938.310 802.000 ;
    END
  END la_output[55]
  PIN la_output[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.050 796.000 955.330 802.000 ;
    END
  END la_output[56]
  PIN la_output[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.610 796.000 971.890 802.000 ;
    END
  END la_output[57]
  PIN la_output[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.630 796.000 988.910 802.000 ;
    END
  END la_output[58]
  PIN la_output[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1005.190 796.000 1005.470 802.000 ;
    END
  END la_output[59]
  PIN la_output[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 796.000 98.350 802.000 ;
    END
  END la_output[5]
  PIN la_output[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1022.210 796.000 1022.490 802.000 ;
    END
  END la_output[60]
  PIN la_output[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1038.770 796.000 1039.050 802.000 ;
    END
  END la_output[61]
  PIN la_output[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1055.790 796.000 1056.070 802.000 ;
    END
  END la_output[62]
  PIN la_output[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 796.000 1072.630 802.000 ;
    END
  END la_output[63]
  PIN la_output[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1089.370 796.000 1089.650 802.000 ;
    END
  END la_output[64]
  PIN la_output[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1105.930 796.000 1106.210 802.000 ;
    END
  END la_output[65]
  PIN la_output[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1122.950 796.000 1123.230 802.000 ;
    END
  END la_output[66]
  PIN la_output[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.510 796.000 1139.790 802.000 ;
    END
  END la_output[67]
  PIN la_output[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.530 796.000 1156.810 802.000 ;
    END
  END la_output[68]
  PIN la_output[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1173.090 796.000 1173.370 802.000 ;
    END
  END la_output[69]
  PIN la_output[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 796.000 115.370 802.000 ;
    END
  END la_output[6]
  PIN la_output[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1190.110 796.000 1190.390 802.000 ;
    END
  END la_output[70]
  PIN la_output[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1206.670 796.000 1206.950 802.000 ;
    END
  END la_output[71]
  PIN la_output[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1223.690 796.000 1223.970 802.000 ;
    END
  END la_output[72]
  PIN la_output[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1240.250 796.000 1240.530 802.000 ;
    END
  END la_output[73]
  PIN la_output[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.270 796.000 1257.550 802.000 ;
    END
  END la_output[74]
  PIN la_output[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.830 796.000 1274.110 802.000 ;
    END
  END la_output[75]
  PIN la_output[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1290.850 796.000 1291.130 802.000 ;
    END
  END la_output[76]
  PIN la_output[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1307.410 796.000 1307.690 802.000 ;
    END
  END la_output[77]
  PIN la_output[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1324.430 796.000 1324.710 802.000 ;
    END
  END la_output[78]
  PIN la_output[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.990 796.000 1341.270 802.000 ;
    END
  END la_output[79]
  PIN la_output[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 796.000 131.930 802.000 ;
    END
  END la_output[7]
  PIN la_output[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.010 796.000 1358.290 802.000 ;
    END
  END la_output[80]
  PIN la_output[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1374.570 796.000 1374.850 802.000 ;
    END
  END la_output[81]
  PIN la_output[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.590 796.000 1391.870 802.000 ;
    END
  END la_output[82]
  PIN la_output[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1408.150 796.000 1408.430 802.000 ;
    END
  END la_output[83]
  PIN la_output[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1425.170 796.000 1425.450 802.000 ;
    END
  END la_output[84]
  PIN la_output[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1441.730 796.000 1442.010 802.000 ;
    END
  END la_output[85]
  PIN la_output[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1458.750 796.000 1459.030 802.000 ;
    END
  END la_output[86]
  PIN la_output[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1475.770 796.000 1476.050 802.000 ;
    END
  END la_output[87]
  PIN la_output[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.330 796.000 1492.610 802.000 ;
    END
  END la_output[88]
  PIN la_output[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1509.350 796.000 1509.630 802.000 ;
    END
  END la_output[89]
  PIN la_output[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 796.000 148.950 802.000 ;
    END
  END la_output[8]
  PIN la_output[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1525.910 796.000 1526.190 802.000 ;
    END
  END la_output[90]
  PIN la_output[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.930 796.000 1543.210 802.000 ;
    END
  END la_output[91]
  PIN la_output[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1559.490 796.000 1559.770 802.000 ;
    END
  END la_output[92]
  PIN la_output[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1576.510 796.000 1576.790 802.000 ;
    END
  END la_output[93]
  PIN la_output[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1593.070 796.000 1593.350 802.000 ;
    END
  END la_output[94]
  PIN la_output[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.090 796.000 1610.370 802.000 ;
    END
  END la_output[95]
  PIN la_output[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1626.650 796.000 1626.930 802.000 ;
    END
  END la_output[96]
  PIN la_output[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1643.670 796.000 1643.950 802.000 ;
    END
  END la_output[97]
  PIN la_output[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1660.230 796.000 1660.510 802.000 ;
    END
  END la_output[98]
  PIN la_output[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1677.250 796.000 1677.530 802.000 ;
    END
  END la_output[99]
  PIN la_output[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 796.000 165.970 802.000 ;
    END
  END la_output[9]
  PIN mprj_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2151.510 796.000 2151.790 802.000 ;
    END
  END mprj_ack_i
  PIN mprj_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2172.670 796.000 2172.950 802.000 ;
    END
  END mprj_adr_o[0]
  PIN mprj_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2315.270 796.000 2315.550 802.000 ;
    END
  END mprj_adr_o[10]
  PIN mprj_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2328.150 796.000 2328.430 802.000 ;
    END
  END mprj_adr_o[11]
  PIN mprj_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2340.570 796.000 2340.850 802.000 ;
    END
  END mprj_adr_o[12]
  PIN mprj_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2352.990 796.000 2353.270 802.000 ;
    END
  END mprj_adr_o[13]
  PIN mprj_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2365.870 796.000 2366.150 802.000 ;
    END
  END mprj_adr_o[14]
  PIN mprj_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2378.290 796.000 2378.570 802.000 ;
    END
  END mprj_adr_o[15]
  PIN mprj_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2390.710 796.000 2390.990 802.000 ;
    END
  END mprj_adr_o[16]
  PIN mprj_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2403.590 796.000 2403.870 802.000 ;
    END
  END mprj_adr_o[17]
  PIN mprj_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2416.010 796.000 2416.290 802.000 ;
    END
  END mprj_adr_o[18]
  PIN mprj_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2428.890 796.000 2429.170 802.000 ;
    END
  END mprj_adr_o[19]
  PIN mprj_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2189.230 796.000 2189.510 802.000 ;
    END
  END mprj_adr_o[1]
  PIN mprj_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2441.310 796.000 2441.590 802.000 ;
    END
  END mprj_adr_o[20]
  PIN mprj_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2453.730 796.000 2454.010 802.000 ;
    END
  END mprj_adr_o[21]
  PIN mprj_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2466.610 796.000 2466.890 802.000 ;
    END
  END mprj_adr_o[22]
  PIN mprj_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2479.030 796.000 2479.310 802.000 ;
    END
  END mprj_adr_o[23]
  PIN mprj_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2491.910 796.000 2492.190 802.000 ;
    END
  END mprj_adr_o[24]
  PIN mprj_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2504.330 796.000 2504.610 802.000 ;
    END
  END mprj_adr_o[25]
  PIN mprj_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2516.750 796.000 2517.030 802.000 ;
    END
  END mprj_adr_o[26]
  PIN mprj_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2529.630 796.000 2529.910 802.000 ;
    END
  END mprj_adr_o[27]
  PIN mprj_adr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2542.050 796.000 2542.330 802.000 ;
    END
  END mprj_adr_o[28]
  PIN mprj_adr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2554.470 796.000 2554.750 802.000 ;
    END
  END mprj_adr_o[29]
  PIN mprj_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2206.250 796.000 2206.530 802.000 ;
    END
  END mprj_adr_o[2]
  PIN mprj_adr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2567.350 796.000 2567.630 802.000 ;
    END
  END mprj_adr_o[30]
  PIN mprj_adr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2579.770 796.000 2580.050 802.000 ;
    END
  END mprj_adr_o[31]
  PIN mprj_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2222.810 796.000 2223.090 802.000 ;
    END
  END mprj_adr_o[3]
  PIN mprj_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2239.830 796.000 2240.110 802.000 ;
    END
  END mprj_adr_o[4]
  PIN mprj_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2252.250 796.000 2252.530 802.000 ;
    END
  END mprj_adr_o[5]
  PIN mprj_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2265.130 796.000 2265.410 802.000 ;
    END
  END mprj_adr_o[6]
  PIN mprj_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2277.550 796.000 2277.830 802.000 ;
    END
  END mprj_adr_o[7]
  PIN mprj_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2289.970 796.000 2290.250 802.000 ;
    END
  END mprj_adr_o[8]
  PIN mprj_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2302.850 796.000 2303.130 802.000 ;
    END
  END mprj_adr_o[9]
  PIN mprj_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2155.650 796.000 2155.930 802.000 ;
    END
  END mprj_cyc_o
  PIN mprj_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2176.810 796.000 2177.090 802.000 ;
    END
  END mprj_dat_i[0]
  PIN mprj_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2319.410 796.000 2319.690 802.000 ;
    END
  END mprj_dat_i[10]
  PIN mprj_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2332.290 796.000 2332.570 802.000 ;
    END
  END mprj_dat_i[11]
  PIN mprj_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2344.710 796.000 2344.990 802.000 ;
    END
  END mprj_dat_i[12]
  PIN mprj_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2357.130 796.000 2357.410 802.000 ;
    END
  END mprj_dat_i[13]
  PIN mprj_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2370.010 796.000 2370.290 802.000 ;
    END
  END mprj_dat_i[14]
  PIN mprj_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2382.430 796.000 2382.710 802.000 ;
    END
  END mprj_dat_i[15]
  PIN mprj_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2395.310 796.000 2395.590 802.000 ;
    END
  END mprj_dat_i[16]
  PIN mprj_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2407.730 796.000 2408.010 802.000 ;
    END
  END mprj_dat_i[17]
  PIN mprj_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2420.150 796.000 2420.430 802.000 ;
    END
  END mprj_dat_i[18]
  PIN mprj_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2433.030 796.000 2433.310 802.000 ;
    END
  END mprj_dat_i[19]
  PIN mprj_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2193.370 796.000 2193.650 802.000 ;
    END
  END mprj_dat_i[1]
  PIN mprj_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2445.450 796.000 2445.730 802.000 ;
    END
  END mprj_dat_i[20]
  PIN mprj_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2458.330 796.000 2458.610 802.000 ;
    END
  END mprj_dat_i[21]
  PIN mprj_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2470.750 796.000 2471.030 802.000 ;
    END
  END mprj_dat_i[22]
  PIN mprj_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2483.170 796.000 2483.450 802.000 ;
    END
  END mprj_dat_i[23]
  PIN mprj_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2496.050 796.000 2496.330 802.000 ;
    END
  END mprj_dat_i[24]
  PIN mprj_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2508.470 796.000 2508.750 802.000 ;
    END
  END mprj_dat_i[25]
  PIN mprj_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2520.890 796.000 2521.170 802.000 ;
    END
  END mprj_dat_i[26]
  PIN mprj_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2533.770 796.000 2534.050 802.000 ;
    END
  END mprj_dat_i[27]
  PIN mprj_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2546.190 796.000 2546.470 802.000 ;
    END
  END mprj_dat_i[28]
  PIN mprj_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2559.070 796.000 2559.350 802.000 ;
    END
  END mprj_dat_i[29]
  PIN mprj_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2210.390 796.000 2210.670 802.000 ;
    END
  END mprj_dat_i[2]
  PIN mprj_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2571.490 796.000 2571.770 802.000 ;
    END
  END mprj_dat_i[30]
  PIN mprj_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2583.910 796.000 2584.190 802.000 ;
    END
  END mprj_dat_i[31]
  PIN mprj_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2226.950 796.000 2227.230 802.000 ;
    END
  END mprj_dat_i[3]
  PIN mprj_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2243.970 796.000 2244.250 802.000 ;
    END
  END mprj_dat_i[4]
  PIN mprj_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2256.390 796.000 2256.670 802.000 ;
    END
  END mprj_dat_i[5]
  PIN mprj_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2269.270 796.000 2269.550 802.000 ;
    END
  END mprj_dat_i[6]
  PIN mprj_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2281.690 796.000 2281.970 802.000 ;
    END
  END mprj_dat_i[7]
  PIN mprj_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2294.570 796.000 2294.850 802.000 ;
    END
  END mprj_dat_i[8]
  PIN mprj_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2306.990 796.000 2307.270 802.000 ;
    END
  END mprj_dat_i[9]
  PIN mprj_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2180.950 796.000 2181.230 802.000 ;
    END
  END mprj_dat_o[0]
  PIN mprj_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2323.550 796.000 2323.830 802.000 ;
    END
  END mprj_dat_o[10]
  PIN mprj_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2336.430 796.000 2336.710 802.000 ;
    END
  END mprj_dat_o[11]
  PIN mprj_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2348.850 796.000 2349.130 802.000 ;
    END
  END mprj_dat_o[12]
  PIN mprj_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2361.730 796.000 2362.010 802.000 ;
    END
  END mprj_dat_o[13]
  PIN mprj_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2374.150 796.000 2374.430 802.000 ;
    END
  END mprj_dat_o[14]
  PIN mprj_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2386.570 796.000 2386.850 802.000 ;
    END
  END mprj_dat_o[15]
  PIN mprj_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2399.450 796.000 2399.730 802.000 ;
    END
  END mprj_dat_o[16]
  PIN mprj_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2411.870 796.000 2412.150 802.000 ;
    END
  END mprj_dat_o[17]
  PIN mprj_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2424.290 796.000 2424.570 802.000 ;
    END
  END mprj_dat_o[18]
  PIN mprj_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2437.170 796.000 2437.450 802.000 ;
    END
  END mprj_dat_o[19]
  PIN mprj_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2197.970 796.000 2198.250 802.000 ;
    END
  END mprj_dat_o[1]
  PIN mprj_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2449.590 796.000 2449.870 802.000 ;
    END
  END mprj_dat_o[20]
  PIN mprj_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2462.470 796.000 2462.750 802.000 ;
    END
  END mprj_dat_o[21]
  PIN mprj_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2474.890 796.000 2475.170 802.000 ;
    END
  END mprj_dat_o[22]
  PIN mprj_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2487.310 796.000 2487.590 802.000 ;
    END
  END mprj_dat_o[23]
  PIN mprj_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2500.190 796.000 2500.470 802.000 ;
    END
  END mprj_dat_o[24]
  PIN mprj_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2512.610 796.000 2512.890 802.000 ;
    END
  END mprj_dat_o[25]
  PIN mprj_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2525.490 796.000 2525.770 802.000 ;
    END
  END mprj_dat_o[26]
  PIN mprj_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2537.910 796.000 2538.190 802.000 ;
    END
  END mprj_dat_o[27]
  PIN mprj_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2550.330 796.000 2550.610 802.000 ;
    END
  END mprj_dat_o[28]
  PIN mprj_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2563.210 796.000 2563.490 802.000 ;
    END
  END mprj_dat_o[29]
  PIN mprj_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2214.530 796.000 2214.810 802.000 ;
    END
  END mprj_dat_o[2]
  PIN mprj_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2575.630 796.000 2575.910 802.000 ;
    END
  END mprj_dat_o[30]
  PIN mprj_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2588.050 796.000 2588.330 802.000 ;
    END
  END mprj_dat_o[31]
  PIN mprj_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2231.550 796.000 2231.830 802.000 ;
    END
  END mprj_dat_o[3]
  PIN mprj_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2248.110 796.000 2248.390 802.000 ;
    END
  END mprj_dat_o[4]
  PIN mprj_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2260.530 796.000 2260.810 802.000 ;
    END
  END mprj_dat_o[5]
  PIN mprj_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2273.410 796.000 2273.690 802.000 ;
    END
  END mprj_dat_o[6]
  PIN mprj_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2285.830 796.000 2286.110 802.000 ;
    END
  END mprj_dat_o[7]
  PIN mprj_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2298.710 796.000 2298.990 802.000 ;
    END
  END mprj_dat_o[8]
  PIN mprj_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2311.130 796.000 2311.410 802.000 ;
    END
  END mprj_dat_o[9]
  PIN mprj_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2185.090 796.000 2185.370 802.000 ;
    END
  END mprj_sel_o[0]
  PIN mprj_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2202.110 796.000 2202.390 802.000 ;
    END
  END mprj_sel_o[1]
  PIN mprj_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.670 796.000 2218.950 802.000 ;
    END
  END mprj_sel_o[2]
  PIN mprj_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2235.690 796.000 2235.970 802.000 ;
    END
  END mprj_sel_o[3]
  PIN mprj_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2159.790 796.000 2160.070 802.000 ;
    END
  END mprj_stb_o
  PIN mprj_wb_iena
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2164.390 796.000 2164.670 802.000 ;
    END
  END mprj_wb_iena
  PIN mprj_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2168.530 796.000 2168.810 802.000 ;
    END
  END mprj_we_o
  PIN qspi_enabled
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 440.000 2622.000 440.600 ;
    END
  END qspi_enabled
  PIN ser_rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 410.080 2622.000 410.680 ;
    END
  END ser_rx
  PIN ser_tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 417.560 2622.000 418.160 ;
    END
  END ser_tx
  PIN spi_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 395.800 2622.000 396.400 ;
    END
  END spi_csb
  PIN spi_enabled
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 425.040 2622.000 425.640 ;
    END
  END spi_enabled
  PIN spi_sck
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 388.320 2622.000 388.920 ;
    END
  END spi_sck
  PIN spi_sdi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 403.280 2622.000 403.880 ;
    END
  END spi_sdi
  PIN spi_sdo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 380.840 2622.000 381.440 ;
    END
  END spi_sdo
  PIN spi_sdoenb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 373.360 2622.000 373.960 ;
    END
  END spi_sdoenb
  PIN sram_ro_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 10.240 2622.000 10.840 ;
    END
  END sram_ro_addr[0]
  PIN sram_ro_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 17.720 2622.000 18.320 ;
    END
  END sram_ro_addr[1]
  PIN sram_ro_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 25.200 2622.000 25.800 ;
    END
  END sram_ro_addr[2]
  PIN sram_ro_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 32.680 2622.000 33.280 ;
    END
  END sram_ro_addr[3]
  PIN sram_ro_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 40.160 2622.000 40.760 ;
    END
  END sram_ro_addr[4]
  PIN sram_ro_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 47.640 2622.000 48.240 ;
    END
  END sram_ro_addr[5]
  PIN sram_ro_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 55.120 2622.000 55.720 ;
    END
  END sram_ro_addr[6]
  PIN sram_ro_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 62.600 2622.000 63.200 ;
    END
  END sram_ro_addr[7]
  PIN sram_ro_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 70.080 2622.000 70.680 ;
    END
  END sram_ro_clk
  PIN sram_ro_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 3.440 2622.000 4.040 ;
    END
  END sram_ro_csb
  PIN sram_ro_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 76.880 2622.000 77.480 ;
    END
  END sram_ro_data[0]
  PIN sram_ro_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 151.000 2622.000 151.600 ;
    END
  END sram_ro_data[10]
  PIN sram_ro_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 158.480 2622.000 159.080 ;
    END
  END sram_ro_data[11]
  PIN sram_ro_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 165.960 2622.000 166.560 ;
    END
  END sram_ro_data[12]
  PIN sram_ro_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 173.440 2622.000 174.040 ;
    END
  END sram_ro_data[13]
  PIN sram_ro_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 180.920 2622.000 181.520 ;
    END
  END sram_ro_data[14]
  PIN sram_ro_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 188.400 2622.000 189.000 ;
    END
  END sram_ro_data[15]
  PIN sram_ro_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 195.880 2622.000 196.480 ;
    END
  END sram_ro_data[16]
  PIN sram_ro_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 203.360 2622.000 203.960 ;
    END
  END sram_ro_data[17]
  PIN sram_ro_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 210.160 2622.000 210.760 ;
    END
  END sram_ro_data[18]
  PIN sram_ro_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 217.640 2622.000 218.240 ;
    END
  END sram_ro_data[19]
  PIN sram_ro_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 84.360 2622.000 84.960 ;
    END
  END sram_ro_data[1]
  PIN sram_ro_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 225.120 2622.000 225.720 ;
    END
  END sram_ro_data[20]
  PIN sram_ro_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 232.600 2622.000 233.200 ;
    END
  END sram_ro_data[21]
  PIN sram_ro_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 240.080 2622.000 240.680 ;
    END
  END sram_ro_data[22]
  PIN sram_ro_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 247.560 2622.000 248.160 ;
    END
  END sram_ro_data[23]
  PIN sram_ro_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 255.040 2622.000 255.640 ;
    END
  END sram_ro_data[24]
  PIN sram_ro_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 262.520 2622.000 263.120 ;
    END
  END sram_ro_data[25]
  PIN sram_ro_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 270.000 2622.000 270.600 ;
    END
  END sram_ro_data[26]
  PIN sram_ro_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 276.800 2622.000 277.400 ;
    END
  END sram_ro_data[27]
  PIN sram_ro_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 284.280 2622.000 284.880 ;
    END
  END sram_ro_data[28]
  PIN sram_ro_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 291.760 2622.000 292.360 ;
    END
  END sram_ro_data[29]
  PIN sram_ro_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 91.840 2622.000 92.440 ;
    END
  END sram_ro_data[2]
  PIN sram_ro_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 299.240 2622.000 299.840 ;
    END
  END sram_ro_data[30]
  PIN sram_ro_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 306.720 2622.000 307.320 ;
    END
  END sram_ro_data[31]
  PIN sram_ro_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 99.320 2622.000 99.920 ;
    END
  END sram_ro_data[3]
  PIN sram_ro_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 106.800 2622.000 107.400 ;
    END
  END sram_ro_data[4]
  PIN sram_ro_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 114.280 2622.000 114.880 ;
    END
  END sram_ro_data[5]
  PIN sram_ro_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 121.760 2622.000 122.360 ;
    END
  END sram_ro_data[6]
  PIN sram_ro_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 129.240 2622.000 129.840 ;
    END
  END sram_ro_data[7]
  PIN sram_ro_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 136.720 2622.000 137.320 ;
    END
  END sram_ro_data[8]
  PIN sram_ro_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 143.520 2622.000 144.120 ;
    END
  END sram_ro_data[9]
  PIN trap
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 343.440 2622.000 344.040 ;
    END
  END trap
  PIN uart_enabled
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 432.520 2622.000 433.120 ;
    END
  END uart_enabled
  PIN user_irq_ena[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2592.650 796.000 2592.930 802.000 ;
    END
  END user_irq_ena[0]
  PIN user_irq_ena[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2596.790 796.000 2597.070 802.000 ;
    END
  END user_irq_ena[1]
  PIN user_irq_ena[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2600.930 796.000 2601.210 802.000 ;
    END
  END user_irq_ena[2]
  OBS
      LAYER li1 ;
        RECT 14.345 20.795 2584.500 739.045 ;
      LAYER met1 ;
        RECT 1.910 1.740 2617.790 792.840 ;
      LAYER met2 ;
        RECT 2.490 795.720 5.790 796.690 ;
        RECT 6.630 795.720 9.930 796.690 ;
        RECT 10.770 795.720 14.070 796.690 ;
        RECT 14.910 795.720 18.210 796.690 ;
        RECT 19.050 795.720 22.350 796.690 ;
        RECT 23.190 795.720 26.490 796.690 ;
        RECT 27.330 795.720 30.630 796.690 ;
        RECT 31.470 795.720 35.230 796.690 ;
        RECT 36.070 795.720 39.370 796.690 ;
        RECT 40.210 795.720 43.510 796.690 ;
        RECT 44.350 795.720 47.650 796.690 ;
        RECT 48.490 795.720 51.790 796.690 ;
        RECT 52.630 795.720 55.930 796.690 ;
        RECT 56.770 795.720 60.070 796.690 ;
        RECT 60.910 795.720 64.210 796.690 ;
        RECT 65.050 795.720 68.810 796.690 ;
        RECT 69.650 795.720 72.950 796.690 ;
        RECT 73.790 795.720 77.090 796.690 ;
        RECT 77.930 795.720 81.230 796.690 ;
        RECT 82.070 795.720 85.370 796.690 ;
        RECT 86.210 795.720 89.510 796.690 ;
        RECT 90.350 795.720 93.650 796.690 ;
        RECT 94.490 795.720 97.790 796.690 ;
        RECT 98.630 795.720 102.390 796.690 ;
        RECT 103.230 795.720 106.530 796.690 ;
        RECT 107.370 795.720 110.670 796.690 ;
        RECT 111.510 795.720 114.810 796.690 ;
        RECT 115.650 795.720 118.950 796.690 ;
        RECT 119.790 795.720 123.090 796.690 ;
        RECT 123.930 795.720 127.230 796.690 ;
        RECT 128.070 795.720 131.370 796.690 ;
        RECT 132.210 795.720 135.970 796.690 ;
        RECT 136.810 795.720 140.110 796.690 ;
        RECT 140.950 795.720 144.250 796.690 ;
        RECT 145.090 795.720 148.390 796.690 ;
        RECT 149.230 795.720 152.530 796.690 ;
        RECT 153.370 795.720 156.670 796.690 ;
        RECT 157.510 795.720 160.810 796.690 ;
        RECT 161.650 795.720 165.410 796.690 ;
        RECT 166.250 795.720 169.550 796.690 ;
        RECT 170.390 795.720 173.690 796.690 ;
        RECT 174.530 795.720 177.830 796.690 ;
        RECT 178.670 795.720 181.970 796.690 ;
        RECT 182.810 795.720 186.110 796.690 ;
        RECT 186.950 795.720 190.250 796.690 ;
        RECT 191.090 795.720 194.390 796.690 ;
        RECT 195.230 795.720 198.990 796.690 ;
        RECT 199.830 795.720 203.130 796.690 ;
        RECT 203.970 795.720 207.270 796.690 ;
        RECT 208.110 795.720 211.410 796.690 ;
        RECT 212.250 795.720 215.550 796.690 ;
        RECT 216.390 795.720 219.690 796.690 ;
        RECT 220.530 795.720 223.830 796.690 ;
        RECT 224.670 795.720 227.970 796.690 ;
        RECT 228.810 795.720 232.570 796.690 ;
        RECT 233.410 795.720 236.710 796.690 ;
        RECT 237.550 795.720 240.850 796.690 ;
        RECT 241.690 795.720 244.990 796.690 ;
        RECT 245.830 795.720 249.130 796.690 ;
        RECT 249.970 795.720 253.270 796.690 ;
        RECT 254.110 795.720 257.410 796.690 ;
        RECT 258.250 795.720 261.550 796.690 ;
        RECT 262.390 795.720 266.150 796.690 ;
        RECT 266.990 795.720 270.290 796.690 ;
        RECT 271.130 795.720 274.430 796.690 ;
        RECT 275.270 795.720 278.570 796.690 ;
        RECT 279.410 795.720 282.710 796.690 ;
        RECT 283.550 795.720 286.850 796.690 ;
        RECT 287.690 795.720 290.990 796.690 ;
        RECT 291.830 795.720 295.130 796.690 ;
        RECT 295.970 795.720 299.730 796.690 ;
        RECT 300.570 795.720 303.870 796.690 ;
        RECT 304.710 795.720 308.010 796.690 ;
        RECT 308.850 795.720 312.150 796.690 ;
        RECT 312.990 795.720 316.290 796.690 ;
        RECT 317.130 795.720 320.430 796.690 ;
        RECT 321.270 795.720 324.570 796.690 ;
        RECT 325.410 795.720 329.170 796.690 ;
        RECT 330.010 795.720 333.310 796.690 ;
        RECT 334.150 795.720 337.450 796.690 ;
        RECT 338.290 795.720 341.590 796.690 ;
        RECT 342.430 795.720 345.730 796.690 ;
        RECT 346.570 795.720 349.870 796.690 ;
        RECT 350.710 795.720 354.010 796.690 ;
        RECT 354.850 795.720 358.150 796.690 ;
        RECT 358.990 795.720 362.750 796.690 ;
        RECT 363.590 795.720 366.890 796.690 ;
        RECT 367.730 795.720 371.030 796.690 ;
        RECT 371.870 795.720 375.170 796.690 ;
        RECT 376.010 795.720 379.310 796.690 ;
        RECT 380.150 795.720 383.450 796.690 ;
        RECT 384.290 795.720 387.590 796.690 ;
        RECT 388.430 795.720 391.730 796.690 ;
        RECT 392.570 795.720 396.330 796.690 ;
        RECT 397.170 795.720 400.470 796.690 ;
        RECT 401.310 795.720 404.610 796.690 ;
        RECT 405.450 795.720 408.750 796.690 ;
        RECT 409.590 795.720 412.890 796.690 ;
        RECT 413.730 795.720 417.030 796.690 ;
        RECT 417.870 795.720 421.170 796.690 ;
        RECT 422.010 795.720 425.310 796.690 ;
        RECT 426.150 795.720 429.910 796.690 ;
        RECT 430.750 795.720 434.050 796.690 ;
        RECT 434.890 795.720 438.190 796.690 ;
        RECT 439.030 795.720 442.330 796.690 ;
        RECT 443.170 795.720 446.470 796.690 ;
        RECT 447.310 795.720 450.610 796.690 ;
        RECT 451.450 795.720 454.750 796.690 ;
        RECT 455.590 795.720 458.890 796.690 ;
        RECT 459.730 795.720 463.490 796.690 ;
        RECT 464.330 795.720 467.630 796.690 ;
        RECT 468.470 795.720 471.770 796.690 ;
        RECT 472.610 795.720 475.910 796.690 ;
        RECT 476.750 795.720 480.050 796.690 ;
        RECT 480.890 795.720 484.190 796.690 ;
        RECT 485.030 795.720 488.330 796.690 ;
        RECT 489.170 795.720 492.930 796.690 ;
        RECT 493.770 795.720 497.070 796.690 ;
        RECT 497.910 795.720 501.210 796.690 ;
        RECT 502.050 795.720 505.350 796.690 ;
        RECT 506.190 795.720 509.490 796.690 ;
        RECT 510.330 795.720 513.630 796.690 ;
        RECT 514.470 795.720 517.770 796.690 ;
        RECT 518.610 795.720 521.910 796.690 ;
        RECT 522.750 795.720 526.510 796.690 ;
        RECT 527.350 795.720 530.650 796.690 ;
        RECT 531.490 795.720 534.790 796.690 ;
        RECT 535.630 795.720 538.930 796.690 ;
        RECT 539.770 795.720 543.070 796.690 ;
        RECT 543.910 795.720 547.210 796.690 ;
        RECT 548.050 795.720 551.350 796.690 ;
        RECT 552.190 795.720 555.490 796.690 ;
        RECT 556.330 795.720 560.090 796.690 ;
        RECT 560.930 795.720 564.230 796.690 ;
        RECT 565.070 795.720 568.370 796.690 ;
        RECT 569.210 795.720 572.510 796.690 ;
        RECT 573.350 795.720 576.650 796.690 ;
        RECT 577.490 795.720 580.790 796.690 ;
        RECT 581.630 795.720 584.930 796.690 ;
        RECT 585.770 795.720 589.070 796.690 ;
        RECT 589.910 795.720 593.670 796.690 ;
        RECT 594.510 795.720 597.810 796.690 ;
        RECT 598.650 795.720 601.950 796.690 ;
        RECT 602.790 795.720 606.090 796.690 ;
        RECT 606.930 795.720 610.230 796.690 ;
        RECT 611.070 795.720 614.370 796.690 ;
        RECT 615.210 795.720 618.510 796.690 ;
        RECT 619.350 795.720 622.650 796.690 ;
        RECT 623.490 795.720 627.250 796.690 ;
        RECT 628.090 795.720 631.390 796.690 ;
        RECT 632.230 795.720 635.530 796.690 ;
        RECT 636.370 795.720 639.670 796.690 ;
        RECT 640.510 795.720 643.810 796.690 ;
        RECT 644.650 795.720 647.950 796.690 ;
        RECT 648.790 795.720 652.090 796.690 ;
        RECT 652.930 795.720 656.690 796.690 ;
        RECT 657.530 795.720 660.830 796.690 ;
        RECT 661.670 795.720 664.970 796.690 ;
        RECT 665.810 795.720 669.110 796.690 ;
        RECT 669.950 795.720 673.250 796.690 ;
        RECT 674.090 795.720 677.390 796.690 ;
        RECT 678.230 795.720 681.530 796.690 ;
        RECT 682.370 795.720 685.670 796.690 ;
        RECT 686.510 795.720 690.270 796.690 ;
        RECT 691.110 795.720 694.410 796.690 ;
        RECT 695.250 795.720 698.550 796.690 ;
        RECT 699.390 795.720 702.690 796.690 ;
        RECT 703.530 795.720 706.830 796.690 ;
        RECT 707.670 795.720 710.970 796.690 ;
        RECT 711.810 795.720 715.110 796.690 ;
        RECT 715.950 795.720 719.250 796.690 ;
        RECT 720.090 795.720 723.850 796.690 ;
        RECT 724.690 795.720 727.990 796.690 ;
        RECT 728.830 795.720 732.130 796.690 ;
        RECT 732.970 795.720 736.270 796.690 ;
        RECT 737.110 795.720 740.410 796.690 ;
        RECT 741.250 795.720 744.550 796.690 ;
        RECT 745.390 795.720 748.690 796.690 ;
        RECT 749.530 795.720 752.830 796.690 ;
        RECT 753.670 795.720 757.430 796.690 ;
        RECT 758.270 795.720 761.570 796.690 ;
        RECT 762.410 795.720 765.710 796.690 ;
        RECT 766.550 795.720 769.850 796.690 ;
        RECT 770.690 795.720 773.990 796.690 ;
        RECT 774.830 795.720 778.130 796.690 ;
        RECT 778.970 795.720 782.270 796.690 ;
        RECT 783.110 795.720 786.410 796.690 ;
        RECT 787.250 795.720 791.010 796.690 ;
        RECT 791.850 795.720 795.150 796.690 ;
        RECT 795.990 795.720 799.290 796.690 ;
        RECT 800.130 795.720 803.430 796.690 ;
        RECT 804.270 795.720 807.570 796.690 ;
        RECT 808.410 795.720 811.710 796.690 ;
        RECT 812.550 795.720 815.850 796.690 ;
        RECT 816.690 795.720 820.450 796.690 ;
        RECT 821.290 795.720 824.590 796.690 ;
        RECT 825.430 795.720 828.730 796.690 ;
        RECT 829.570 795.720 832.870 796.690 ;
        RECT 833.710 795.720 837.010 796.690 ;
        RECT 837.850 795.720 841.150 796.690 ;
        RECT 841.990 795.720 845.290 796.690 ;
        RECT 846.130 795.720 849.430 796.690 ;
        RECT 850.270 795.720 854.030 796.690 ;
        RECT 854.870 795.720 858.170 796.690 ;
        RECT 859.010 795.720 862.310 796.690 ;
        RECT 863.150 795.720 866.450 796.690 ;
        RECT 867.290 795.720 870.590 796.690 ;
        RECT 871.430 795.720 874.730 796.690 ;
        RECT 875.570 795.720 878.870 796.690 ;
        RECT 879.710 795.720 883.010 796.690 ;
        RECT 883.850 795.720 887.610 796.690 ;
        RECT 888.450 795.720 891.750 796.690 ;
        RECT 892.590 795.720 895.890 796.690 ;
        RECT 896.730 795.720 900.030 796.690 ;
        RECT 900.870 795.720 904.170 796.690 ;
        RECT 905.010 795.720 908.310 796.690 ;
        RECT 909.150 795.720 912.450 796.690 ;
        RECT 913.290 795.720 916.590 796.690 ;
        RECT 917.430 795.720 921.190 796.690 ;
        RECT 922.030 795.720 925.330 796.690 ;
        RECT 926.170 795.720 929.470 796.690 ;
        RECT 930.310 795.720 933.610 796.690 ;
        RECT 934.450 795.720 937.750 796.690 ;
        RECT 938.590 795.720 941.890 796.690 ;
        RECT 942.730 795.720 946.030 796.690 ;
        RECT 946.870 795.720 950.170 796.690 ;
        RECT 951.010 795.720 954.770 796.690 ;
        RECT 955.610 795.720 958.910 796.690 ;
        RECT 959.750 795.720 963.050 796.690 ;
        RECT 963.890 795.720 967.190 796.690 ;
        RECT 968.030 795.720 971.330 796.690 ;
        RECT 972.170 795.720 975.470 796.690 ;
        RECT 976.310 795.720 979.610 796.690 ;
        RECT 980.450 795.720 984.210 796.690 ;
        RECT 985.050 795.720 988.350 796.690 ;
        RECT 989.190 795.720 992.490 796.690 ;
        RECT 993.330 795.720 996.630 796.690 ;
        RECT 997.470 795.720 1000.770 796.690 ;
        RECT 1001.610 795.720 1004.910 796.690 ;
        RECT 1005.750 795.720 1009.050 796.690 ;
        RECT 1009.890 795.720 1013.190 796.690 ;
        RECT 1014.030 795.720 1017.790 796.690 ;
        RECT 1018.630 795.720 1021.930 796.690 ;
        RECT 1022.770 795.720 1026.070 796.690 ;
        RECT 1026.910 795.720 1030.210 796.690 ;
        RECT 1031.050 795.720 1034.350 796.690 ;
        RECT 1035.190 795.720 1038.490 796.690 ;
        RECT 1039.330 795.720 1042.630 796.690 ;
        RECT 1043.470 795.720 1046.770 796.690 ;
        RECT 1047.610 795.720 1051.370 796.690 ;
        RECT 1052.210 795.720 1055.510 796.690 ;
        RECT 1056.350 795.720 1059.650 796.690 ;
        RECT 1060.490 795.720 1063.790 796.690 ;
        RECT 1064.630 795.720 1067.930 796.690 ;
        RECT 1068.770 795.720 1072.070 796.690 ;
        RECT 1072.910 795.720 1076.210 796.690 ;
        RECT 1077.050 795.720 1080.350 796.690 ;
        RECT 1081.190 795.720 1084.950 796.690 ;
        RECT 1085.790 795.720 1089.090 796.690 ;
        RECT 1089.930 795.720 1093.230 796.690 ;
        RECT 1094.070 795.720 1097.370 796.690 ;
        RECT 1098.210 795.720 1101.510 796.690 ;
        RECT 1102.350 795.720 1105.650 796.690 ;
        RECT 1106.490 795.720 1109.790 796.690 ;
        RECT 1110.630 795.720 1113.930 796.690 ;
        RECT 1114.770 795.720 1118.530 796.690 ;
        RECT 1119.370 795.720 1122.670 796.690 ;
        RECT 1123.510 795.720 1126.810 796.690 ;
        RECT 1127.650 795.720 1130.950 796.690 ;
        RECT 1131.790 795.720 1135.090 796.690 ;
        RECT 1135.930 795.720 1139.230 796.690 ;
        RECT 1140.070 795.720 1143.370 796.690 ;
        RECT 1144.210 795.720 1147.970 796.690 ;
        RECT 1148.810 795.720 1152.110 796.690 ;
        RECT 1152.950 795.720 1156.250 796.690 ;
        RECT 1157.090 795.720 1160.390 796.690 ;
        RECT 1161.230 795.720 1164.530 796.690 ;
        RECT 1165.370 795.720 1168.670 796.690 ;
        RECT 1169.510 795.720 1172.810 796.690 ;
        RECT 1173.650 795.720 1176.950 796.690 ;
        RECT 1177.790 795.720 1181.550 796.690 ;
        RECT 1182.390 795.720 1185.690 796.690 ;
        RECT 1186.530 795.720 1189.830 796.690 ;
        RECT 1190.670 795.720 1193.970 796.690 ;
        RECT 1194.810 795.720 1198.110 796.690 ;
        RECT 1198.950 795.720 1202.250 796.690 ;
        RECT 1203.090 795.720 1206.390 796.690 ;
        RECT 1207.230 795.720 1210.530 796.690 ;
        RECT 1211.370 795.720 1215.130 796.690 ;
        RECT 1215.970 795.720 1219.270 796.690 ;
        RECT 1220.110 795.720 1223.410 796.690 ;
        RECT 1224.250 795.720 1227.550 796.690 ;
        RECT 1228.390 795.720 1231.690 796.690 ;
        RECT 1232.530 795.720 1235.830 796.690 ;
        RECT 1236.670 795.720 1239.970 796.690 ;
        RECT 1240.810 795.720 1244.110 796.690 ;
        RECT 1244.950 795.720 1248.710 796.690 ;
        RECT 1249.550 795.720 1252.850 796.690 ;
        RECT 1253.690 795.720 1256.990 796.690 ;
        RECT 1257.830 795.720 1261.130 796.690 ;
        RECT 1261.970 795.720 1265.270 796.690 ;
        RECT 1266.110 795.720 1269.410 796.690 ;
        RECT 1270.250 795.720 1273.550 796.690 ;
        RECT 1274.390 795.720 1277.690 796.690 ;
        RECT 1278.530 795.720 1282.290 796.690 ;
        RECT 1283.130 795.720 1286.430 796.690 ;
        RECT 1287.270 795.720 1290.570 796.690 ;
        RECT 1291.410 795.720 1294.710 796.690 ;
        RECT 1295.550 795.720 1298.850 796.690 ;
        RECT 1299.690 795.720 1302.990 796.690 ;
        RECT 1303.830 795.720 1307.130 796.690 ;
        RECT 1307.970 795.720 1311.730 796.690 ;
        RECT 1312.570 795.720 1315.870 796.690 ;
        RECT 1316.710 795.720 1320.010 796.690 ;
        RECT 1320.850 795.720 1324.150 796.690 ;
        RECT 1324.990 795.720 1328.290 796.690 ;
        RECT 1329.130 795.720 1332.430 796.690 ;
        RECT 1333.270 795.720 1336.570 796.690 ;
        RECT 1337.410 795.720 1340.710 796.690 ;
        RECT 1341.550 795.720 1345.310 796.690 ;
        RECT 1346.150 795.720 1349.450 796.690 ;
        RECT 1350.290 795.720 1353.590 796.690 ;
        RECT 1354.430 795.720 1357.730 796.690 ;
        RECT 1358.570 795.720 1361.870 796.690 ;
        RECT 1362.710 795.720 1366.010 796.690 ;
        RECT 1366.850 795.720 1370.150 796.690 ;
        RECT 1370.990 795.720 1374.290 796.690 ;
        RECT 1375.130 795.720 1378.890 796.690 ;
        RECT 1379.730 795.720 1383.030 796.690 ;
        RECT 1383.870 795.720 1387.170 796.690 ;
        RECT 1388.010 795.720 1391.310 796.690 ;
        RECT 1392.150 795.720 1395.450 796.690 ;
        RECT 1396.290 795.720 1399.590 796.690 ;
        RECT 1400.430 795.720 1403.730 796.690 ;
        RECT 1404.570 795.720 1407.870 796.690 ;
        RECT 1408.710 795.720 1412.470 796.690 ;
        RECT 1413.310 795.720 1416.610 796.690 ;
        RECT 1417.450 795.720 1420.750 796.690 ;
        RECT 1421.590 795.720 1424.890 796.690 ;
        RECT 1425.730 795.720 1429.030 796.690 ;
        RECT 1429.870 795.720 1433.170 796.690 ;
        RECT 1434.010 795.720 1437.310 796.690 ;
        RECT 1438.150 795.720 1441.450 796.690 ;
        RECT 1442.290 795.720 1446.050 796.690 ;
        RECT 1446.890 795.720 1450.190 796.690 ;
        RECT 1451.030 795.720 1454.330 796.690 ;
        RECT 1455.170 795.720 1458.470 796.690 ;
        RECT 1459.310 795.720 1462.610 796.690 ;
        RECT 1463.450 795.720 1466.750 796.690 ;
        RECT 1467.590 795.720 1470.890 796.690 ;
        RECT 1471.730 795.720 1475.490 796.690 ;
        RECT 1476.330 795.720 1479.630 796.690 ;
        RECT 1480.470 795.720 1483.770 796.690 ;
        RECT 1484.610 795.720 1487.910 796.690 ;
        RECT 1488.750 795.720 1492.050 796.690 ;
        RECT 1492.890 795.720 1496.190 796.690 ;
        RECT 1497.030 795.720 1500.330 796.690 ;
        RECT 1501.170 795.720 1504.470 796.690 ;
        RECT 1505.310 795.720 1509.070 796.690 ;
        RECT 1509.910 795.720 1513.210 796.690 ;
        RECT 1514.050 795.720 1517.350 796.690 ;
        RECT 1518.190 795.720 1521.490 796.690 ;
        RECT 1522.330 795.720 1525.630 796.690 ;
        RECT 1526.470 795.720 1529.770 796.690 ;
        RECT 1530.610 795.720 1533.910 796.690 ;
        RECT 1534.750 795.720 1538.050 796.690 ;
        RECT 1538.890 795.720 1542.650 796.690 ;
        RECT 1543.490 795.720 1546.790 796.690 ;
        RECT 1547.630 795.720 1550.930 796.690 ;
        RECT 1551.770 795.720 1555.070 796.690 ;
        RECT 1555.910 795.720 1559.210 796.690 ;
        RECT 1560.050 795.720 1563.350 796.690 ;
        RECT 1564.190 795.720 1567.490 796.690 ;
        RECT 1568.330 795.720 1571.630 796.690 ;
        RECT 1572.470 795.720 1576.230 796.690 ;
        RECT 1577.070 795.720 1580.370 796.690 ;
        RECT 1581.210 795.720 1584.510 796.690 ;
        RECT 1585.350 795.720 1588.650 796.690 ;
        RECT 1589.490 795.720 1592.790 796.690 ;
        RECT 1593.630 795.720 1596.930 796.690 ;
        RECT 1597.770 795.720 1601.070 796.690 ;
        RECT 1601.910 795.720 1605.210 796.690 ;
        RECT 1606.050 795.720 1609.810 796.690 ;
        RECT 1610.650 795.720 1613.950 796.690 ;
        RECT 1614.790 795.720 1618.090 796.690 ;
        RECT 1618.930 795.720 1622.230 796.690 ;
        RECT 1623.070 795.720 1626.370 796.690 ;
        RECT 1627.210 795.720 1630.510 796.690 ;
        RECT 1631.350 795.720 1634.650 796.690 ;
        RECT 1635.490 795.720 1639.250 796.690 ;
        RECT 1640.090 795.720 1643.390 796.690 ;
        RECT 1644.230 795.720 1647.530 796.690 ;
        RECT 1648.370 795.720 1651.670 796.690 ;
        RECT 1652.510 795.720 1655.810 796.690 ;
        RECT 1656.650 795.720 1659.950 796.690 ;
        RECT 1660.790 795.720 1664.090 796.690 ;
        RECT 1664.930 795.720 1668.230 796.690 ;
        RECT 1669.070 795.720 1672.830 796.690 ;
        RECT 1673.670 795.720 1676.970 796.690 ;
        RECT 1677.810 795.720 1681.110 796.690 ;
        RECT 1681.950 795.720 1685.250 796.690 ;
        RECT 1686.090 795.720 1689.390 796.690 ;
        RECT 1690.230 795.720 1693.530 796.690 ;
        RECT 1694.370 795.720 1697.670 796.690 ;
        RECT 1698.510 795.720 1701.810 796.690 ;
        RECT 1702.650 795.720 1706.410 796.690 ;
        RECT 1707.250 795.720 1710.550 796.690 ;
        RECT 1711.390 795.720 1714.690 796.690 ;
        RECT 1715.530 795.720 1718.830 796.690 ;
        RECT 1719.670 795.720 1722.970 796.690 ;
        RECT 1723.810 795.720 1727.110 796.690 ;
        RECT 1727.950 795.720 1731.250 796.690 ;
        RECT 1732.090 795.720 1735.390 796.690 ;
        RECT 1736.230 795.720 1739.990 796.690 ;
        RECT 1740.830 795.720 1744.130 796.690 ;
        RECT 1744.970 795.720 1748.270 796.690 ;
        RECT 1749.110 795.720 1752.410 796.690 ;
        RECT 1753.250 795.720 1756.550 796.690 ;
        RECT 1757.390 795.720 1760.690 796.690 ;
        RECT 1761.530 795.720 1764.830 796.690 ;
        RECT 1765.670 795.720 1768.970 796.690 ;
        RECT 1769.810 795.720 1773.570 796.690 ;
        RECT 1774.410 795.720 1777.710 796.690 ;
        RECT 1778.550 795.720 1781.850 796.690 ;
        RECT 1782.690 795.720 1785.990 796.690 ;
        RECT 1786.830 795.720 1790.130 796.690 ;
        RECT 1790.970 795.720 1794.270 796.690 ;
        RECT 1795.110 795.720 1798.410 796.690 ;
        RECT 1799.250 795.720 1803.010 796.690 ;
        RECT 1803.850 795.720 1807.150 796.690 ;
        RECT 1807.990 795.720 1811.290 796.690 ;
        RECT 1812.130 795.720 1815.430 796.690 ;
        RECT 1816.270 795.720 1819.570 796.690 ;
        RECT 1820.410 795.720 1823.710 796.690 ;
        RECT 1824.550 795.720 1827.850 796.690 ;
        RECT 1828.690 795.720 1831.990 796.690 ;
        RECT 1832.830 795.720 1836.590 796.690 ;
        RECT 1837.430 795.720 1840.730 796.690 ;
        RECT 1841.570 795.720 1844.870 796.690 ;
        RECT 1845.710 795.720 1849.010 796.690 ;
        RECT 1849.850 795.720 1853.150 796.690 ;
        RECT 1853.990 795.720 1857.290 796.690 ;
        RECT 1858.130 795.720 1861.430 796.690 ;
        RECT 1862.270 795.720 1865.570 796.690 ;
        RECT 1866.410 795.720 1870.170 796.690 ;
        RECT 1871.010 795.720 1874.310 796.690 ;
        RECT 1875.150 795.720 1878.450 796.690 ;
        RECT 1879.290 795.720 1882.590 796.690 ;
        RECT 1883.430 795.720 1886.730 796.690 ;
        RECT 1887.570 795.720 1890.870 796.690 ;
        RECT 1891.710 795.720 1895.010 796.690 ;
        RECT 1895.850 795.720 1899.150 796.690 ;
        RECT 1899.990 795.720 1903.750 796.690 ;
        RECT 1904.590 795.720 1907.890 796.690 ;
        RECT 1908.730 795.720 1912.030 796.690 ;
        RECT 1912.870 795.720 1916.170 796.690 ;
        RECT 1917.010 795.720 1920.310 796.690 ;
        RECT 1921.150 795.720 1924.450 796.690 ;
        RECT 1925.290 795.720 1928.590 796.690 ;
        RECT 1929.430 795.720 1932.730 796.690 ;
        RECT 1933.570 795.720 1937.330 796.690 ;
        RECT 1938.170 795.720 1941.470 796.690 ;
        RECT 1942.310 795.720 1945.610 796.690 ;
        RECT 1946.450 795.720 1949.750 796.690 ;
        RECT 1950.590 795.720 1953.890 796.690 ;
        RECT 1954.730 795.720 1958.030 796.690 ;
        RECT 1958.870 795.720 1962.170 796.690 ;
        RECT 1963.010 795.720 1966.770 796.690 ;
        RECT 1967.610 795.720 1970.910 796.690 ;
        RECT 1971.750 795.720 1975.050 796.690 ;
        RECT 1975.890 795.720 1979.190 796.690 ;
        RECT 1980.030 795.720 1983.330 796.690 ;
        RECT 1984.170 795.720 1987.470 796.690 ;
        RECT 1988.310 795.720 1991.610 796.690 ;
        RECT 1992.450 795.720 1995.750 796.690 ;
        RECT 1996.590 795.720 2000.350 796.690 ;
        RECT 2001.190 795.720 2004.490 796.690 ;
        RECT 2005.330 795.720 2008.630 796.690 ;
        RECT 2009.470 795.720 2012.770 796.690 ;
        RECT 2013.610 795.720 2016.910 796.690 ;
        RECT 2017.750 795.720 2021.050 796.690 ;
        RECT 2021.890 795.720 2025.190 796.690 ;
        RECT 2026.030 795.720 2029.330 796.690 ;
        RECT 2030.170 795.720 2033.930 796.690 ;
        RECT 2034.770 795.720 2038.070 796.690 ;
        RECT 2038.910 795.720 2042.210 796.690 ;
        RECT 2043.050 795.720 2046.350 796.690 ;
        RECT 2047.190 795.720 2050.490 796.690 ;
        RECT 2051.330 795.720 2054.630 796.690 ;
        RECT 2055.470 795.720 2058.770 796.690 ;
        RECT 2059.610 795.720 2062.910 796.690 ;
        RECT 2063.750 795.720 2067.510 796.690 ;
        RECT 2068.350 795.720 2071.650 796.690 ;
        RECT 2072.490 795.720 2075.790 796.690 ;
        RECT 2076.630 795.720 2079.930 796.690 ;
        RECT 2080.770 795.720 2084.070 796.690 ;
        RECT 2084.910 795.720 2088.210 796.690 ;
        RECT 2089.050 795.720 2092.350 796.690 ;
        RECT 2093.190 795.720 2096.490 796.690 ;
        RECT 2097.330 795.720 2101.090 796.690 ;
        RECT 2101.930 795.720 2105.230 796.690 ;
        RECT 2106.070 795.720 2109.370 796.690 ;
        RECT 2110.210 795.720 2113.510 796.690 ;
        RECT 2114.350 795.720 2117.650 796.690 ;
        RECT 2118.490 795.720 2121.790 796.690 ;
        RECT 2122.630 795.720 2125.930 796.690 ;
        RECT 2126.770 795.720 2130.530 796.690 ;
        RECT 2131.370 795.720 2134.670 796.690 ;
        RECT 2135.510 795.720 2138.810 796.690 ;
        RECT 2139.650 795.720 2142.950 796.690 ;
        RECT 2143.790 795.720 2147.090 796.690 ;
        RECT 2147.930 795.720 2151.230 796.690 ;
        RECT 2152.070 795.720 2155.370 796.690 ;
        RECT 2156.210 795.720 2159.510 796.690 ;
        RECT 2160.350 795.720 2164.110 796.690 ;
        RECT 2164.950 795.720 2168.250 796.690 ;
        RECT 2169.090 795.720 2172.390 796.690 ;
        RECT 2173.230 795.720 2176.530 796.690 ;
        RECT 2177.370 795.720 2180.670 796.690 ;
        RECT 2181.510 795.720 2184.810 796.690 ;
        RECT 2185.650 795.720 2188.950 796.690 ;
        RECT 2189.790 795.720 2193.090 796.690 ;
        RECT 2193.930 795.720 2197.690 796.690 ;
        RECT 2198.530 795.720 2201.830 796.690 ;
        RECT 2202.670 795.720 2205.970 796.690 ;
        RECT 2206.810 795.720 2210.110 796.690 ;
        RECT 2210.950 795.720 2214.250 796.690 ;
        RECT 2215.090 795.720 2218.390 796.690 ;
        RECT 2219.230 795.720 2222.530 796.690 ;
        RECT 2223.370 795.720 2226.670 796.690 ;
        RECT 2227.510 795.720 2231.270 796.690 ;
        RECT 2232.110 795.720 2235.410 796.690 ;
        RECT 2236.250 795.720 2239.550 796.690 ;
        RECT 2240.390 795.720 2243.690 796.690 ;
        RECT 2244.530 795.720 2247.830 796.690 ;
        RECT 2248.670 795.720 2251.970 796.690 ;
        RECT 2252.810 795.720 2256.110 796.690 ;
        RECT 2256.950 795.720 2260.250 796.690 ;
        RECT 2261.090 795.720 2264.850 796.690 ;
        RECT 2265.690 795.720 2268.990 796.690 ;
        RECT 2269.830 795.720 2273.130 796.690 ;
        RECT 2273.970 795.720 2277.270 796.690 ;
        RECT 2278.110 795.720 2281.410 796.690 ;
        RECT 2282.250 795.720 2285.550 796.690 ;
        RECT 2286.390 795.720 2289.690 796.690 ;
        RECT 2290.530 795.720 2294.290 796.690 ;
        RECT 2295.130 795.720 2298.430 796.690 ;
        RECT 2299.270 795.720 2302.570 796.690 ;
        RECT 2303.410 795.720 2306.710 796.690 ;
        RECT 2307.550 795.720 2310.850 796.690 ;
        RECT 2311.690 795.720 2314.990 796.690 ;
        RECT 2315.830 795.720 2319.130 796.690 ;
        RECT 2319.970 795.720 2323.270 796.690 ;
        RECT 2324.110 795.720 2327.870 796.690 ;
        RECT 2328.710 795.720 2332.010 796.690 ;
        RECT 2332.850 795.720 2336.150 796.690 ;
        RECT 2336.990 795.720 2340.290 796.690 ;
        RECT 2341.130 795.720 2344.430 796.690 ;
        RECT 2345.270 795.720 2348.570 796.690 ;
        RECT 2349.410 795.720 2352.710 796.690 ;
        RECT 2353.550 795.720 2356.850 796.690 ;
        RECT 2357.690 795.720 2361.450 796.690 ;
        RECT 2362.290 795.720 2365.590 796.690 ;
        RECT 2366.430 795.720 2369.730 796.690 ;
        RECT 2370.570 795.720 2373.870 796.690 ;
        RECT 2374.710 795.720 2378.010 796.690 ;
        RECT 2378.850 795.720 2382.150 796.690 ;
        RECT 2382.990 795.720 2386.290 796.690 ;
        RECT 2387.130 795.720 2390.430 796.690 ;
        RECT 2391.270 795.720 2395.030 796.690 ;
        RECT 2395.870 795.720 2399.170 796.690 ;
        RECT 2400.010 795.720 2403.310 796.690 ;
        RECT 2404.150 795.720 2407.450 796.690 ;
        RECT 2408.290 795.720 2411.590 796.690 ;
        RECT 2412.430 795.720 2415.730 796.690 ;
        RECT 2416.570 795.720 2419.870 796.690 ;
        RECT 2420.710 795.720 2424.010 796.690 ;
        RECT 2424.850 795.720 2428.610 796.690 ;
        RECT 2429.450 795.720 2432.750 796.690 ;
        RECT 2433.590 795.720 2436.890 796.690 ;
        RECT 2437.730 795.720 2441.030 796.690 ;
        RECT 2441.870 795.720 2445.170 796.690 ;
        RECT 2446.010 795.720 2449.310 796.690 ;
        RECT 2450.150 795.720 2453.450 796.690 ;
        RECT 2454.290 795.720 2458.050 796.690 ;
        RECT 2458.890 795.720 2462.190 796.690 ;
        RECT 2463.030 795.720 2466.330 796.690 ;
        RECT 2467.170 795.720 2470.470 796.690 ;
        RECT 2471.310 795.720 2474.610 796.690 ;
        RECT 2475.450 795.720 2478.750 796.690 ;
        RECT 2479.590 795.720 2482.890 796.690 ;
        RECT 2483.730 795.720 2487.030 796.690 ;
        RECT 2487.870 795.720 2491.630 796.690 ;
        RECT 2492.470 795.720 2495.770 796.690 ;
        RECT 2496.610 795.720 2499.910 796.690 ;
        RECT 2500.750 795.720 2504.050 796.690 ;
        RECT 2504.890 795.720 2508.190 796.690 ;
        RECT 2509.030 795.720 2512.330 796.690 ;
        RECT 2513.170 795.720 2516.470 796.690 ;
        RECT 2517.310 795.720 2520.610 796.690 ;
        RECT 2521.450 795.720 2525.210 796.690 ;
        RECT 2526.050 795.720 2529.350 796.690 ;
        RECT 2530.190 795.720 2533.490 796.690 ;
        RECT 2534.330 795.720 2537.630 796.690 ;
        RECT 2538.470 795.720 2541.770 796.690 ;
        RECT 2542.610 795.720 2545.910 796.690 ;
        RECT 2546.750 795.720 2550.050 796.690 ;
        RECT 2550.890 795.720 2554.190 796.690 ;
        RECT 2555.030 795.720 2558.790 796.690 ;
        RECT 2559.630 795.720 2562.930 796.690 ;
        RECT 2563.770 795.720 2567.070 796.690 ;
        RECT 2567.910 795.720 2571.210 796.690 ;
        RECT 2572.050 795.720 2575.350 796.690 ;
        RECT 2576.190 795.720 2579.490 796.690 ;
        RECT 2580.330 795.720 2583.630 796.690 ;
        RECT 2584.470 795.720 2587.770 796.690 ;
        RECT 2588.610 795.720 2592.370 796.690 ;
        RECT 2593.210 795.720 2596.510 796.690 ;
        RECT 2597.350 795.720 2600.650 796.690 ;
        RECT 2601.490 795.720 2604.790 796.690 ;
        RECT 2605.630 795.720 2608.930 796.690 ;
        RECT 2609.770 795.720 2613.070 796.690 ;
        RECT 2613.910 795.720 2617.210 796.690 ;
        RECT 1.940 4.280 2617.760 795.720 ;
        RECT 1.940 1.710 163.570 4.280 ;
        RECT 164.410 1.710 491.090 4.280 ;
        RECT 491.930 1.710 818.610 4.280 ;
        RECT 819.450 1.710 1146.130 4.280 ;
        RECT 1146.970 1.710 1473.650 4.280 ;
        RECT 1474.490 1.710 1801.170 4.280 ;
        RECT 1802.010 1.710 2128.690 4.280 ;
        RECT 2129.530 1.710 2456.210 4.280 ;
        RECT 2457.050 1.710 2617.760 4.280 ;
      LAYER met3 ;
        RECT 10.185 795.240 2615.600 796.105 ;
        RECT 10.185 789.160 2616.000 795.240 ;
        RECT 10.185 787.760 2615.600 789.160 ;
        RECT 10.185 781.680 2616.000 787.760 ;
        RECT 10.185 780.280 2615.600 781.680 ;
        RECT 10.185 774.200 2616.000 780.280 ;
        RECT 10.185 772.800 2615.600 774.200 ;
        RECT 10.185 766.720 2616.000 772.800 ;
        RECT 10.185 765.320 2615.600 766.720 ;
        RECT 10.185 759.240 2616.000 765.320 ;
        RECT 10.185 757.840 2615.600 759.240 ;
        RECT 10.185 751.760 2616.000 757.840 ;
        RECT 10.185 750.360 2615.600 751.760 ;
        RECT 10.185 744.280 2616.000 750.360 ;
        RECT 10.185 742.880 2615.600 744.280 ;
        RECT 10.185 737.480 2616.000 742.880 ;
        RECT 10.185 736.080 2615.600 737.480 ;
        RECT 10.185 730.000 2616.000 736.080 ;
        RECT 10.185 728.600 2615.600 730.000 ;
        RECT 10.185 722.520 2616.000 728.600 ;
        RECT 10.185 721.120 2615.600 722.520 ;
        RECT 10.185 715.040 2616.000 721.120 ;
        RECT 10.185 713.640 2615.600 715.040 ;
        RECT 10.185 707.560 2616.000 713.640 ;
        RECT 10.185 706.160 2615.600 707.560 ;
        RECT 10.185 700.080 2616.000 706.160 ;
        RECT 10.185 698.680 2615.600 700.080 ;
        RECT 10.185 692.600 2616.000 698.680 ;
        RECT 10.185 691.200 2615.600 692.600 ;
        RECT 10.185 685.120 2616.000 691.200 ;
        RECT 10.185 683.720 2615.600 685.120 ;
        RECT 10.185 677.640 2616.000 683.720 ;
        RECT 10.185 676.240 2615.600 677.640 ;
        RECT 10.185 670.840 2616.000 676.240 ;
        RECT 10.185 669.440 2615.600 670.840 ;
        RECT 10.185 663.360 2616.000 669.440 ;
        RECT 10.185 661.960 2615.600 663.360 ;
        RECT 10.185 655.880 2616.000 661.960 ;
        RECT 10.185 654.480 2615.600 655.880 ;
        RECT 10.185 648.400 2616.000 654.480 ;
        RECT 10.185 647.000 2615.600 648.400 ;
        RECT 10.185 640.920 2616.000 647.000 ;
        RECT 10.185 639.520 2615.600 640.920 ;
        RECT 10.185 633.440 2616.000 639.520 ;
        RECT 10.185 632.040 2615.600 633.440 ;
        RECT 10.185 625.960 2616.000 632.040 ;
        RECT 10.185 624.560 2615.600 625.960 ;
        RECT 10.185 618.480 2616.000 624.560 ;
        RECT 10.185 617.080 2615.600 618.480 ;
        RECT 10.185 611.000 2616.000 617.080 ;
        RECT 10.185 609.600 2615.600 611.000 ;
        RECT 10.185 604.200 2616.000 609.600 ;
        RECT 10.185 602.800 2615.600 604.200 ;
        RECT 10.185 596.720 2616.000 602.800 ;
        RECT 10.185 595.320 2615.600 596.720 ;
        RECT 10.185 589.240 2616.000 595.320 ;
        RECT 10.185 587.840 2615.600 589.240 ;
        RECT 10.185 581.760 2616.000 587.840 ;
        RECT 10.185 580.360 2615.600 581.760 ;
        RECT 10.185 574.280 2616.000 580.360 ;
        RECT 10.185 572.880 2615.600 574.280 ;
        RECT 10.185 566.800 2616.000 572.880 ;
        RECT 10.185 565.400 2615.600 566.800 ;
        RECT 10.185 559.320 2616.000 565.400 ;
        RECT 10.185 557.920 2615.600 559.320 ;
        RECT 10.185 551.840 2616.000 557.920 ;
        RECT 10.185 550.440 2615.600 551.840 ;
        RECT 10.185 544.360 2616.000 550.440 ;
        RECT 10.185 542.960 2615.600 544.360 ;
        RECT 10.185 537.560 2616.000 542.960 ;
        RECT 10.185 536.160 2615.600 537.560 ;
        RECT 10.185 530.080 2616.000 536.160 ;
        RECT 10.185 528.680 2615.600 530.080 ;
        RECT 10.185 522.600 2616.000 528.680 ;
        RECT 10.185 521.200 2615.600 522.600 ;
        RECT 10.185 515.120 2616.000 521.200 ;
        RECT 10.185 513.720 2615.600 515.120 ;
        RECT 10.185 507.640 2616.000 513.720 ;
        RECT 10.185 506.240 2615.600 507.640 ;
        RECT 10.185 500.160 2616.000 506.240 ;
        RECT 10.185 498.760 2615.600 500.160 ;
        RECT 10.185 492.680 2616.000 498.760 ;
        RECT 10.185 491.280 2615.600 492.680 ;
        RECT 10.185 485.200 2616.000 491.280 ;
        RECT 10.185 483.800 2615.600 485.200 ;
        RECT 10.185 477.720 2616.000 483.800 ;
        RECT 10.185 476.320 2615.600 477.720 ;
        RECT 10.185 470.920 2616.000 476.320 ;
        RECT 10.185 469.520 2615.600 470.920 ;
        RECT 10.185 463.440 2616.000 469.520 ;
        RECT 10.185 462.040 2615.600 463.440 ;
        RECT 10.185 455.960 2616.000 462.040 ;
        RECT 10.185 454.560 2615.600 455.960 ;
        RECT 10.185 448.480 2616.000 454.560 ;
        RECT 10.185 447.080 2615.600 448.480 ;
        RECT 10.185 441.000 2616.000 447.080 ;
        RECT 10.185 439.600 2615.600 441.000 ;
        RECT 10.185 433.520 2616.000 439.600 ;
        RECT 10.185 432.120 2615.600 433.520 ;
        RECT 10.185 426.040 2616.000 432.120 ;
        RECT 10.185 424.640 2615.600 426.040 ;
        RECT 10.185 418.560 2616.000 424.640 ;
        RECT 10.185 417.160 2615.600 418.560 ;
        RECT 10.185 411.080 2616.000 417.160 ;
        RECT 10.185 409.680 2615.600 411.080 ;
        RECT 10.185 404.280 2616.000 409.680 ;
        RECT 10.185 402.880 2615.600 404.280 ;
        RECT 10.185 396.800 2616.000 402.880 ;
        RECT 10.185 395.400 2615.600 396.800 ;
        RECT 10.185 389.320 2616.000 395.400 ;
        RECT 10.185 387.920 2615.600 389.320 ;
        RECT 10.185 381.840 2616.000 387.920 ;
        RECT 10.185 380.440 2615.600 381.840 ;
        RECT 10.185 374.360 2616.000 380.440 ;
        RECT 10.185 372.960 2615.600 374.360 ;
        RECT 10.185 366.880 2616.000 372.960 ;
        RECT 10.185 365.480 2615.600 366.880 ;
        RECT 10.185 359.400 2616.000 365.480 ;
        RECT 10.185 358.000 2615.600 359.400 ;
        RECT 10.185 351.920 2616.000 358.000 ;
        RECT 10.185 350.520 2615.600 351.920 ;
        RECT 10.185 344.440 2616.000 350.520 ;
        RECT 10.185 343.040 2615.600 344.440 ;
        RECT 10.185 337.640 2616.000 343.040 ;
        RECT 10.185 336.240 2615.600 337.640 ;
        RECT 10.185 330.160 2616.000 336.240 ;
        RECT 10.185 328.760 2615.600 330.160 ;
        RECT 10.185 322.680 2616.000 328.760 ;
        RECT 10.185 321.280 2615.600 322.680 ;
        RECT 10.185 315.200 2616.000 321.280 ;
        RECT 10.185 313.800 2615.600 315.200 ;
        RECT 10.185 307.720 2616.000 313.800 ;
        RECT 10.185 306.320 2615.600 307.720 ;
        RECT 10.185 300.240 2616.000 306.320 ;
        RECT 10.185 298.840 2615.600 300.240 ;
        RECT 10.185 292.760 2616.000 298.840 ;
        RECT 10.185 291.360 2615.600 292.760 ;
        RECT 10.185 285.280 2616.000 291.360 ;
        RECT 10.185 283.880 2615.600 285.280 ;
        RECT 10.185 277.800 2616.000 283.880 ;
        RECT 10.185 276.400 2615.600 277.800 ;
        RECT 10.185 271.000 2616.000 276.400 ;
        RECT 10.185 269.600 2615.600 271.000 ;
        RECT 10.185 263.520 2616.000 269.600 ;
        RECT 10.185 262.120 2615.600 263.520 ;
        RECT 10.185 256.040 2616.000 262.120 ;
        RECT 10.185 254.640 2615.600 256.040 ;
        RECT 10.185 248.560 2616.000 254.640 ;
        RECT 10.185 247.160 2615.600 248.560 ;
        RECT 10.185 241.080 2616.000 247.160 ;
        RECT 10.185 239.680 2615.600 241.080 ;
        RECT 10.185 233.600 2616.000 239.680 ;
        RECT 10.185 232.200 2615.600 233.600 ;
        RECT 10.185 226.120 2616.000 232.200 ;
        RECT 10.185 224.720 2615.600 226.120 ;
        RECT 10.185 218.640 2616.000 224.720 ;
        RECT 10.185 217.240 2615.600 218.640 ;
        RECT 10.185 211.160 2616.000 217.240 ;
        RECT 10.185 209.760 2615.600 211.160 ;
        RECT 10.185 204.360 2616.000 209.760 ;
        RECT 10.185 202.960 2615.600 204.360 ;
        RECT 10.185 196.880 2616.000 202.960 ;
        RECT 10.185 195.480 2615.600 196.880 ;
        RECT 10.185 189.400 2616.000 195.480 ;
        RECT 10.185 188.000 2615.600 189.400 ;
        RECT 10.185 181.920 2616.000 188.000 ;
        RECT 10.185 180.520 2615.600 181.920 ;
        RECT 10.185 174.440 2616.000 180.520 ;
        RECT 10.185 173.040 2615.600 174.440 ;
        RECT 10.185 166.960 2616.000 173.040 ;
        RECT 10.185 165.560 2615.600 166.960 ;
        RECT 10.185 159.480 2616.000 165.560 ;
        RECT 10.185 158.080 2615.600 159.480 ;
        RECT 10.185 152.000 2616.000 158.080 ;
        RECT 10.185 150.600 2615.600 152.000 ;
        RECT 10.185 144.520 2616.000 150.600 ;
        RECT 10.185 143.120 2615.600 144.520 ;
        RECT 10.185 137.720 2616.000 143.120 ;
        RECT 10.185 136.320 2615.600 137.720 ;
        RECT 10.185 130.240 2616.000 136.320 ;
        RECT 10.185 128.840 2615.600 130.240 ;
        RECT 10.185 122.760 2616.000 128.840 ;
        RECT 10.185 121.360 2615.600 122.760 ;
        RECT 10.185 115.280 2616.000 121.360 ;
        RECT 10.185 113.880 2615.600 115.280 ;
        RECT 10.185 107.800 2616.000 113.880 ;
        RECT 10.185 106.400 2615.600 107.800 ;
        RECT 10.185 100.320 2616.000 106.400 ;
        RECT 10.185 98.920 2615.600 100.320 ;
        RECT 10.185 92.840 2616.000 98.920 ;
        RECT 10.185 91.440 2615.600 92.840 ;
        RECT 10.185 85.360 2616.000 91.440 ;
        RECT 10.185 83.960 2615.600 85.360 ;
        RECT 10.185 77.880 2616.000 83.960 ;
        RECT 10.185 76.480 2615.600 77.880 ;
        RECT 10.185 71.080 2616.000 76.480 ;
        RECT 10.185 69.680 2615.600 71.080 ;
        RECT 10.185 63.600 2616.000 69.680 ;
        RECT 10.185 62.200 2615.600 63.600 ;
        RECT 10.185 56.120 2616.000 62.200 ;
        RECT 10.185 54.720 2615.600 56.120 ;
        RECT 10.185 48.640 2616.000 54.720 ;
        RECT 10.185 47.240 2615.600 48.640 ;
        RECT 10.185 41.160 2616.000 47.240 ;
        RECT 10.185 39.760 2615.600 41.160 ;
        RECT 10.185 33.680 2616.000 39.760 ;
        RECT 10.185 32.280 2615.600 33.680 ;
        RECT 10.185 26.200 2616.000 32.280 ;
        RECT 10.185 24.800 2615.600 26.200 ;
        RECT 10.185 18.720 2616.000 24.800 ;
        RECT 10.185 17.320 2615.600 18.720 ;
        RECT 10.185 11.240 2616.000 17.320 ;
        RECT 10.185 9.840 2615.600 11.240 ;
        RECT 10.185 4.440 2616.000 9.840 ;
        RECT 10.185 3.575 2615.600 4.440 ;
      LAYER met4 ;
        RECT 5.020 10.780 2594.600 749.060 ;
      LAYER met5 ;
        RECT 5.020 724.080 2594.600 749.060 ;
        RECT 12.600 717.680 547.400 724.080 ;
        RECT 602.600 717.680 2587.400 724.080 ;
        RECT 5.020 659.080 2594.600 717.680 ;
        RECT 12.600 652.680 547.400 659.080 ;
        RECT 602.600 652.680 2587.400 659.080 ;
        RECT 5.020 594.080 2594.600 652.680 ;
        RECT 12.600 587.680 547.400 594.080 ;
        RECT 602.600 587.680 2587.400 594.080 ;
        RECT 5.020 529.080 2594.600 587.680 ;
        RECT 12.600 522.680 547.400 529.080 ;
        RECT 602.600 522.680 2587.400 529.080 ;
        RECT 5.020 464.080 2594.600 522.680 ;
        RECT 12.600 457.680 547.400 464.080 ;
        RECT 602.600 457.680 2587.400 464.080 ;
        RECT 5.020 399.080 2594.600 457.680 ;
        RECT 12.600 392.680 547.400 399.080 ;
        RECT 602.600 392.680 2587.400 399.080 ;
        RECT 5.020 334.080 2594.600 392.680 ;
        RECT 12.600 327.680 547.400 334.080 ;
        RECT 602.600 327.680 2587.400 334.080 ;
        RECT 5.020 269.080 2594.600 327.680 ;
        RECT 12.600 262.680 547.400 269.080 ;
        RECT 602.600 262.680 2587.400 269.080 ;
        RECT 5.020 204.080 2594.600 262.680 ;
        RECT 12.600 197.680 547.400 204.080 ;
        RECT 602.600 197.680 2587.400 204.080 ;
        RECT 5.020 139.080 2594.600 197.680 ;
        RECT 12.600 132.680 547.400 139.080 ;
        RECT 602.600 132.680 2587.400 139.080 ;
        RECT 5.020 74.080 2594.600 132.680 ;
        RECT 12.600 67.680 547.400 74.080 ;
        RECT 602.600 67.680 2587.400 74.080 ;
        RECT 5.020 10.780 2594.600 67.680 ;
  END
END mgmt_core_wrapper
END LIBRARY

