magic
tech sky130A
magscale 1 2
timestamp 1638169271
<< locali >>
rect 165997 156587 166031 157233
rect 166089 156587 166123 157029
rect 172713 156451 172747 157233
rect 173449 156519 173483 157165
rect 173817 156451 173851 157097
rect 175841 156383 175875 157301
rect 485145 157063 485179 157301
rect 180809 156247 180843 156349
rect 180809 156213 180993 156247
rect 183385 155907 183419 156213
rect 191481 156043 191515 156281
rect 197185 156111 197219 156281
rect 200037 155907 200071 156077
rect 212365 155975 212399 156757
rect 485237 156383 485271 157029
rect 214021 156009 214297 156043
rect 214021 155975 214055 156009
rect 108313 155023 108347 155873
rect 183385 155873 183477 155907
rect 185351 155873 185719 155907
rect 127633 155601 127943 155635
rect 127633 155431 127667 155601
rect 127909 155567 127943 155601
rect 125149 155227 125183 155397
rect 109877 154819 109911 154989
rect 127541 153867 127575 155193
rect 127633 154683 127667 155193
rect 127725 154683 127759 155533
rect 127817 155397 128001 155431
rect 127817 155363 127851 155397
rect 133337 155295 133371 155601
rect 133429 155431 133463 155601
rect 133521 155227 133555 155397
rect 133187 155193 133555 155227
rect 136833 155227 136867 155737
rect 137293 155431 137327 155805
rect 155359 155737 156003 155771
rect 137787 155465 138155 155499
rect 138121 155295 138155 155465
rect 146861 154887 146895 155465
rect 146953 155091 146987 155397
rect 148241 155091 148275 155737
rect 155969 155499 156003 155737
rect 156463 155465 156739 155499
rect 156613 154955 156647 155397
rect 156705 154955 156739 155465
rect 166273 155431 166307 155737
rect 172253 154751 172287 155737
rect 175933 154751 175967 155873
rect 182649 155023 182683 155601
rect 185501 154751 185535 155805
rect 185685 155567 185719 155873
rect 219633 155771 219667 155873
rect 248889 155873 249107 155907
rect 222427 155805 222577 155839
rect 185593 155023 185627 155533
rect 187065 154615 187099 154785
rect 187157 154615 187191 155601
rect 195287 155533 195379 155567
rect 195161 154683 195195 154989
rect 195253 154615 195287 154785
rect 195345 154683 195379 155533
rect 213837 154683 213871 155261
rect 229385 155159 229419 155805
rect 233341 155431 233375 155669
rect 233893 155499 233927 155737
rect 239137 155635 239171 155805
rect 241069 155159 241103 155805
rect 248889 155771 248923 155873
rect 243093 155091 243127 155669
rect 127633 153833 128553 153867
rect 127449 153799 127483 153833
rect 127633 153799 127667 153833
rect 127449 153765 127667 153799
rect 130025 153255 130059 153833
rect 137937 153255 137971 153969
rect 161673 153799 161707 154377
rect 243461 154343 243495 155125
rect 243553 155023 243587 155125
rect 243645 154887 243679 155601
rect 248981 155091 249015 155805
rect 249073 155771 249107 155873
rect 249073 155737 249165 155771
rect 262689 155635 262723 155873
rect 262873 155771 262907 155941
rect 249107 155601 249199 155635
rect 249165 155363 249199 155601
rect 249073 154887 249107 155329
rect 243553 154615 243587 154853
rect 245945 154615 245979 154785
rect 164801 154139 164835 154309
rect 187801 153663 187835 154309
rect 197277 153595 197311 153697
rect 243369 153663 243403 154309
rect 248705 153595 248739 154513
rect 248797 154343 248831 154853
rect 248889 154547 248923 154785
rect 252661 154615 252695 155329
rect 262781 155295 262815 155737
rect 262873 154955 262907 155329
rect 261159 154785 261309 154819
rect 261401 154751 261435 154921
rect 262965 154887 262999 155329
rect 263517 154887 263551 155193
rect 268393 155023 268427 155737
rect 269347 155125 269439 155159
rect 269313 154683 269347 154989
rect 269405 154955 269439 155125
rect 272441 155091 272475 155329
rect 269405 154921 269589 154955
rect 249073 153663 249107 154445
rect 272349 153663 272383 155057
rect 272533 154615 272567 155465
rect 272625 154887 272659 155397
rect 277593 155159 277627 155329
rect 277869 155091 277903 155873
rect 278053 155703 278087 155805
rect 280353 155567 280387 155873
rect 287805 155635 287839 155941
rect 280111 155533 280387 155567
rect 287897 155227 287931 155601
rect 272717 154887 272751 155057
rect 275109 154921 275293 154955
rect 275109 154887 275143 154921
rect 281089 154547 281123 154717
rect 282009 154207 282043 155057
rect 289369 154819 289403 155941
rect 296545 155873 296637 155907
rect 296545 155567 296579 155873
rect 296821 155771 296855 155941
rect 296637 155227 296671 155533
rect 293785 154819 293819 154989
rect 296729 154751 296763 155737
rect 407037 155703 407071 155873
rect 301513 155363 301547 155669
rect 297649 153799 297683 154717
rect 300593 154615 300627 155057
rect 301053 154683 301087 155329
rect 301605 155295 301639 155669
rect 301513 155261 301639 155295
rect 301513 155159 301547 155261
rect 307309 154819 307343 155669
rect 307401 154819 307435 155329
rect 417341 154887 417375 155737
rect 417433 154955 417467 155669
rect 425529 155635 425563 155805
rect 428231 155805 428565 155839
rect 426541 155635 426575 155805
rect 417065 154751 417099 154785
rect 417065 154717 417525 154751
rect 300593 154581 300869 154615
rect 130025 153221 130485 153255
rect 137937 153221 138213 153255
rect 166089 152949 166365 152983
rect 166089 152915 166123 152949
rect 149103 152881 149379 152915
rect 149345 152643 149379 152881
rect 578433 152507 578467 154581
rect 190929 152065 191113 152099
rect 190929 151963 190963 152065
rect 16313 150467 16347 151521
rect 43821 150535 43855 151929
rect 57529 151011 57563 151929
rect 60841 151079 60875 151929
rect 64429 151215 64463 151929
rect 67373 150603 67407 151929
rect 74549 150671 74583 151929
rect 78137 150739 78171 151929
rect 85037 150807 85071 151929
rect 91017 151283 91051 151929
rect 95157 150875 95191 151929
rect 105645 150943 105679 151929
rect 192033 151895 192067 151929
rect 192033 151861 192217 151895
rect 177221 151283 177255 151385
rect 107945 5389 108405 5423
rect 65993 4267 66027 4845
rect 86877 3995 86911 4981
rect 107945 4471 107979 5389
rect 108255 5321 108439 5355
rect 108221 4539 108255 5049
rect 108313 4811 108347 5049
rect 108405 4811 108439 5321
rect 168849 4675 168883 5117
rect 474473 4675 474507 5117
rect 518633 4675 518667 5049
rect 107945 3519 107979 3961
rect 114201 3519 114235 3961
rect 114477 3485 114753 3519
rect 114477 2907 114511 3485
rect 121653 2907 121687 3961
rect 125517 3519 125551 4029
rect 125609 3043 125643 3485
rect 126989 2839 127023 3077
rect 127265 2839 127299 3009
rect 127449 2907 127483 3009
rect 127633 2907 127667 4029
rect 165111 3825 165261 3859
rect 141801 3179 141835 3485
rect 156705 3247 156739 3621
rect 400873 3315 400907 3621
rect 417433 2839 417467 3281
rect 431969 3179 432003 3349
<< viali >>
rect 175841 157301 175875 157335
rect 165997 157233 166031 157267
rect 172713 157233 172747 157267
rect 165997 156553 166031 156587
rect 166089 157029 166123 157063
rect 166089 156553 166123 156587
rect 173449 157165 173483 157199
rect 173449 156485 173483 156519
rect 173817 157097 173851 157131
rect 172713 156417 172747 156451
rect 173817 156417 173851 156451
rect 485145 157301 485179 157335
rect 485145 157029 485179 157063
rect 485237 157029 485271 157063
rect 212365 156757 212399 156791
rect 175841 156349 175875 156383
rect 180809 156349 180843 156383
rect 191481 156281 191515 156315
rect 180993 156213 181027 156247
rect 183385 156213 183419 156247
rect 197185 156281 197219 156315
rect 197185 156077 197219 156111
rect 200037 156077 200071 156111
rect 191481 156009 191515 156043
rect 485237 156349 485271 156383
rect 212365 155941 212399 155975
rect 214297 156009 214331 156043
rect 214021 155941 214055 155975
rect 262873 155941 262907 155975
rect 108313 155873 108347 155907
rect 175933 155873 175967 155907
rect 183477 155873 183511 155907
rect 185317 155873 185351 155907
rect 200037 155873 200071 155907
rect 219633 155873 219667 155907
rect 137293 155805 137327 155839
rect 136833 155737 136867 155771
rect 125149 155397 125183 155431
rect 127633 155397 127667 155431
rect 127725 155533 127759 155567
rect 127909 155533 127943 155567
rect 133337 155601 133371 155635
rect 125149 155193 125183 155227
rect 127541 155193 127575 155227
rect 108313 154989 108347 155023
rect 109877 154989 109911 155023
rect 109877 154785 109911 154819
rect 127633 155193 127667 155227
rect 127633 154649 127667 154683
rect 128001 155397 128035 155431
rect 127817 155329 127851 155363
rect 133429 155601 133463 155635
rect 133429 155397 133463 155431
rect 133521 155397 133555 155431
rect 133337 155261 133371 155295
rect 133153 155193 133187 155227
rect 148241 155737 148275 155771
rect 155325 155737 155359 155771
rect 137753 155465 137787 155499
rect 137293 155397 137327 155431
rect 138121 155261 138155 155295
rect 146861 155465 146895 155499
rect 136833 155193 136867 155227
rect 146953 155397 146987 155431
rect 146953 155057 146987 155091
rect 166273 155737 166307 155771
rect 155969 155465 156003 155499
rect 156429 155465 156463 155499
rect 148241 155057 148275 155091
rect 156613 155397 156647 155431
rect 156613 154921 156647 154955
rect 166273 155397 166307 155431
rect 172253 155737 172287 155771
rect 156705 154921 156739 154955
rect 146861 154853 146895 154887
rect 172253 154717 172287 154751
rect 185501 155805 185535 155839
rect 182649 155601 182683 155635
rect 182649 154989 182683 155023
rect 175933 154717 175967 154751
rect 222393 155805 222427 155839
rect 222577 155805 222611 155839
rect 229385 155805 229419 155839
rect 219633 155737 219667 155771
rect 185593 155533 185627 155567
rect 185685 155533 185719 155567
rect 187157 155601 187191 155635
rect 185593 154989 185627 155023
rect 185501 154717 185535 154751
rect 187065 154785 187099 154819
rect 127725 154649 127759 154683
rect 187065 154581 187099 154615
rect 195253 155533 195287 155567
rect 195161 154989 195195 155023
rect 195161 154649 195195 154683
rect 195253 154785 195287 154819
rect 187157 154581 187191 154615
rect 195345 154649 195379 154683
rect 213837 155261 213871 155295
rect 239137 155805 239171 155839
rect 233893 155737 233927 155771
rect 233341 155669 233375 155703
rect 239137 155601 239171 155635
rect 241069 155805 241103 155839
rect 233893 155465 233927 155499
rect 233341 155397 233375 155431
rect 229385 155125 229419 155159
rect 248889 155737 248923 155771
rect 248981 155805 249015 155839
rect 241069 155125 241103 155159
rect 243093 155669 243127 155703
rect 243645 155601 243679 155635
rect 243093 155057 243127 155091
rect 243461 155125 243495 155159
rect 213837 154649 213871 154683
rect 195253 154581 195287 154615
rect 161673 154377 161707 154411
rect 137937 153969 137971 154003
rect 127449 153833 127483 153867
rect 127541 153833 127575 153867
rect 128553 153833 128587 153867
rect 130025 153833 130059 153867
rect 243553 155125 243587 155159
rect 243553 154989 243587 155023
rect 262689 155873 262723 155907
rect 249165 155737 249199 155771
rect 287805 155941 287839 155975
rect 277869 155873 277903 155907
rect 249073 155601 249107 155635
rect 262689 155601 262723 155635
rect 262781 155737 262815 155771
rect 262873 155737 262907 155771
rect 268393 155737 268427 155771
rect 248981 155057 249015 155091
rect 249073 155329 249107 155363
rect 249165 155329 249199 155363
rect 252661 155329 252695 155363
rect 243553 154853 243587 154887
rect 243645 154853 243679 154887
rect 248797 154853 248831 154887
rect 249073 154853 249107 154887
rect 243553 154581 243587 154615
rect 245945 154785 245979 154819
rect 245945 154581 245979 154615
rect 164801 154309 164835 154343
rect 164801 154105 164835 154139
rect 187801 154309 187835 154343
rect 161673 153765 161707 153799
rect 243369 154309 243403 154343
rect 243461 154309 243495 154343
rect 248705 154513 248739 154547
rect 187801 153629 187835 153663
rect 197277 153697 197311 153731
rect 243369 153629 243403 153663
rect 197277 153561 197311 153595
rect 248889 154785 248923 154819
rect 262781 155261 262815 155295
rect 262873 155329 262907 155363
rect 261401 154921 261435 154955
rect 262873 154921 262907 154955
rect 262965 155329 262999 155363
rect 261125 154785 261159 154819
rect 261309 154785 261343 154819
rect 262965 154853 262999 154887
rect 263517 155193 263551 155227
rect 272533 155465 272567 155499
rect 272441 155329 272475 155363
rect 269313 155125 269347 155159
rect 268393 154989 268427 155023
rect 269313 154989 269347 155023
rect 263517 154853 263551 154887
rect 261401 154717 261435 154751
rect 272349 155057 272383 155091
rect 272441 155057 272475 155091
rect 269589 154921 269623 154955
rect 269313 154649 269347 154683
rect 252661 154581 252695 154615
rect 248889 154513 248923 154547
rect 248797 154309 248831 154343
rect 249073 154445 249107 154479
rect 249073 153629 249107 153663
rect 272625 155397 272659 155431
rect 277593 155329 277627 155363
rect 277593 155125 277627 155159
rect 280353 155873 280387 155907
rect 278053 155805 278087 155839
rect 278053 155669 278087 155703
rect 289369 155941 289403 155975
rect 287805 155601 287839 155635
rect 287897 155601 287931 155635
rect 280077 155533 280111 155567
rect 287897 155193 287931 155227
rect 272625 154853 272659 154887
rect 272717 155057 272751 155091
rect 277869 155057 277903 155091
rect 282009 155057 282043 155091
rect 272717 154853 272751 154887
rect 275293 154921 275327 154955
rect 275109 154853 275143 154887
rect 272533 154581 272567 154615
rect 281089 154717 281123 154751
rect 281089 154513 281123 154547
rect 296821 155941 296855 155975
rect 296637 155873 296671 155907
rect 296729 155737 296763 155771
rect 296821 155737 296855 155771
rect 407037 155873 407071 155907
rect 296545 155533 296579 155567
rect 296637 155533 296671 155567
rect 296637 155193 296671 155227
rect 289369 154785 289403 154819
rect 293785 154989 293819 155023
rect 293785 154785 293819 154819
rect 425529 155805 425563 155839
rect 301513 155669 301547 155703
rect 301053 155329 301087 155363
rect 301513 155329 301547 155363
rect 301605 155669 301639 155703
rect 300593 155057 300627 155091
rect 296729 154717 296763 154751
rect 297649 154717 297683 154751
rect 282009 154173 282043 154207
rect 307309 155669 307343 155703
rect 407037 155669 407071 155703
rect 417341 155737 417375 155771
rect 301513 155125 301547 155159
rect 307309 154785 307343 154819
rect 307401 155329 307435 155363
rect 417433 155669 417467 155703
rect 425529 155601 425563 155635
rect 426541 155805 426575 155839
rect 428197 155805 428231 155839
rect 428565 155805 428599 155839
rect 426541 155601 426575 155635
rect 417433 154921 417467 154955
rect 417341 154853 417375 154887
rect 307401 154785 307435 154819
rect 417065 154785 417099 154819
rect 417525 154717 417559 154751
rect 301053 154649 301087 154683
rect 300869 154581 300903 154615
rect 578433 154581 578467 154615
rect 297649 153765 297683 153799
rect 272349 153629 272383 153663
rect 248705 153561 248739 153595
rect 130485 153221 130519 153255
rect 138213 153221 138247 153255
rect 166365 152949 166399 152983
rect 149069 152881 149103 152915
rect 166089 152881 166123 152915
rect 149345 152609 149379 152643
rect 578433 152473 578467 152507
rect 191113 152065 191147 152099
rect 43821 151929 43855 151963
rect 16313 151521 16347 151555
rect 57529 151929 57563 151963
rect 60841 151929 60875 151963
rect 64429 151929 64463 151963
rect 64429 151181 64463 151215
rect 67373 151929 67407 151963
rect 60841 151045 60875 151079
rect 57529 150977 57563 151011
rect 74549 151929 74583 151963
rect 78137 151929 78171 151963
rect 85037 151929 85071 151963
rect 91017 151929 91051 151963
rect 91017 151249 91051 151283
rect 95157 151929 95191 151963
rect 105645 151929 105679 151963
rect 190929 151929 190963 151963
rect 192033 151929 192067 151963
rect 192217 151861 192251 151895
rect 177221 151385 177255 151419
rect 177221 151249 177255 151283
rect 105645 150909 105679 150943
rect 95157 150841 95191 150875
rect 85037 150773 85071 150807
rect 78137 150705 78171 150739
rect 74549 150637 74583 150671
rect 67373 150569 67407 150603
rect 43821 150501 43855 150535
rect 16313 150433 16347 150467
rect 108405 5389 108439 5423
rect 86877 4981 86911 5015
rect 65993 4845 66027 4879
rect 65993 4233 66027 4267
rect 108221 5321 108255 5355
rect 108221 5049 108255 5083
rect 108313 5049 108347 5083
rect 108313 4777 108347 4811
rect 108405 4777 108439 4811
rect 168849 5117 168883 5151
rect 168849 4641 168883 4675
rect 474473 5117 474507 5151
rect 474473 4641 474507 4675
rect 518633 5049 518667 5083
rect 518633 4641 518667 4675
rect 108221 4505 108255 4539
rect 107945 4437 107979 4471
rect 125517 4029 125551 4063
rect 86877 3961 86911 3995
rect 107945 3961 107979 3995
rect 107945 3485 107979 3519
rect 114201 3961 114235 3995
rect 121653 3961 121687 3995
rect 114201 3485 114235 3519
rect 114753 3485 114787 3519
rect 114477 2873 114511 2907
rect 127633 4029 127667 4063
rect 125517 3485 125551 3519
rect 125609 3485 125643 3519
rect 125609 3009 125643 3043
rect 126989 3077 127023 3111
rect 121653 2873 121687 2907
rect 126989 2805 127023 2839
rect 127265 3009 127299 3043
rect 127449 3009 127483 3043
rect 127449 2873 127483 2907
rect 165077 3825 165111 3859
rect 165261 3825 165295 3859
rect 156705 3621 156739 3655
rect 141801 3485 141835 3519
rect 400873 3621 400907 3655
rect 431969 3349 432003 3383
rect 400873 3281 400907 3315
rect 417433 3281 417467 3315
rect 156705 3213 156739 3247
rect 141801 3145 141835 3179
rect 127633 2873 127667 2907
rect 127265 2805 127299 2839
rect 431969 3145 432003 3179
rect 417433 2805 417467 2839
<< metal1 >>
rect 26786 158856 26792 158908
rect 26844 158896 26850 158908
rect 137462 158896 137468 158908
rect 26844 158868 137468 158896
rect 26844 158856 26850 158868
rect 137462 158856 137468 158868
rect 137520 158856 137526 158908
rect 15194 158788 15200 158840
rect 15252 158828 15258 158840
rect 129734 158828 129740 158840
rect 15252 158800 129740 158828
rect 15252 158788 15258 158800
rect 129734 158788 129740 158800
rect 129792 158788 129798 158840
rect 22830 158720 22836 158772
rect 22888 158760 22894 158772
rect 134886 158760 134892 158772
rect 22888 158732 134892 158760
rect 22888 158720 22894 158732
rect 134886 158720 134892 158732
rect 134944 158720 134950 158772
rect 11146 158652 11152 158704
rect 11204 158692 11210 158704
rect 127066 158692 127072 158704
rect 11204 158664 127072 158692
rect 11204 158652 11210 158664
rect 127066 158652 127072 158664
rect 127124 158652 127130 158704
rect 82814 158584 82820 158636
rect 82872 158624 82878 158636
rect 164234 158624 164240 158636
rect 82872 158596 164240 158624
rect 82872 158584 82878 158596
rect 164234 158584 164240 158596
rect 164292 158584 164298 158636
rect 70394 158516 70400 158568
rect 70452 158556 70458 158568
rect 156322 158556 156328 158568
rect 70452 158528 156328 158556
rect 70452 158516 70458 158528
rect 156322 158516 156328 158528
rect 156380 158516 156386 158568
rect 74994 158448 75000 158500
rect 75052 158488 75058 158500
rect 161658 158488 161664 158500
rect 75052 158460 161664 158488
rect 75052 158448 75058 158460
rect 161658 158448 161664 158460
rect 161716 158448 161722 158500
rect 67358 158380 67364 158432
rect 67416 158420 67422 158432
rect 153746 158420 153752 158432
rect 67416 158392 153752 158420
rect 67416 158380 67422 158392
rect 153746 158380 153752 158392
rect 153804 158380 153810 158432
rect 51074 158312 51080 158364
rect 51132 158352 51138 158364
rect 148686 158352 148692 158364
rect 51132 158324 148692 158352
rect 51132 158312 51138 158324
rect 148686 158312 148692 158324
rect 148744 158312 148750 158364
rect 34514 158244 34520 158296
rect 34572 158284 34578 158296
rect 142798 158284 142804 158296
rect 34572 158256 142804 158284
rect 34572 158244 34578 158256
rect 142798 158244 142804 158256
rect 142856 158244 142862 158296
rect 12434 158176 12440 158228
rect 12492 158216 12498 158228
rect 122834 158216 122840 158228
rect 12492 158188 122840 158216
rect 12492 158176 12498 158188
rect 122834 158176 122840 158188
rect 122892 158176 122898 158228
rect 18966 158108 18972 158160
rect 19024 158148 19030 158160
rect 132586 158148 132592 158160
rect 19024 158120 132592 158148
rect 19024 158108 19030 158120
rect 132586 158108 132592 158120
rect 132644 158108 132650 158160
rect 112530 158040 112536 158092
rect 112588 158080 112594 158092
rect 194778 158080 194784 158092
rect 112588 158052 194784 158080
rect 112588 158040 112594 158052
rect 194778 158040 194784 158052
rect 194836 158040 194842 158092
rect 94038 157972 94044 158024
rect 94096 158012 94102 158024
rect 182358 158012 182364 158024
rect 94096 157984 182364 158012
rect 94096 157972 94102 157984
rect 182358 157972 182364 157984
rect 182416 157972 182422 158024
rect 82262 157904 82268 157956
rect 82320 157944 82326 157956
rect 174538 157944 174544 157956
rect 82320 157916 174544 157944
rect 82320 157904 82326 157916
rect 174538 157904 174544 157916
rect 174596 157904 174602 157956
rect 58894 157836 58900 157888
rect 58952 157876 58958 157888
rect 158990 157876 158996 157888
rect 58952 157848 158996 157876
rect 58952 157836 58958 157848
rect 158990 157836 158996 157848
rect 159048 157836 159054 157888
rect 47210 157768 47216 157820
rect 47268 157808 47274 157820
rect 151170 157808 151176 157820
rect 47268 157780 151176 157808
rect 47268 157768 47274 157780
rect 151170 157768 151176 157780
rect 151228 157768 151234 157820
rect 38470 157700 38476 157752
rect 38528 157740 38534 157752
rect 145282 157740 145288 157752
rect 38528 157712 145288 157740
rect 38528 157700 38534 157712
rect 145282 157700 145288 157712
rect 145340 157700 145346 157752
rect 148594 157700 148600 157752
rect 148652 157740 148658 157752
rect 218882 157740 218888 157752
rect 148652 157712 218888 157740
rect 148652 157700 148658 157712
rect 218882 157700 218888 157712
rect 218940 157700 218946 157752
rect 30650 157632 30656 157684
rect 30708 157672 30714 157684
rect 140130 157672 140136 157684
rect 30708 157644 140136 157672
rect 30708 157632 30714 157644
rect 140130 157632 140136 157644
rect 140188 157632 140194 157684
rect 140774 157632 140780 157684
rect 140832 157672 140838 157684
rect 214098 157672 214104 157684
rect 140832 157644 214104 157672
rect 140832 157632 140838 157644
rect 214098 157632 214104 157644
rect 214156 157632 214162 157684
rect 129090 157564 129096 157616
rect 129148 157604 129154 157616
rect 205818 157604 205824 157616
rect 129148 157576 205824 157604
rect 129148 157564 129154 157576
rect 205818 157564 205824 157576
rect 205876 157564 205882 157616
rect 113542 157496 113548 157548
rect 113600 157536 113606 157548
rect 195422 157536 195428 157548
rect 113600 157508 195428 157536
rect 113600 157496 113606 157508
rect 195422 157496 195428 157508
rect 195480 157496 195486 157548
rect 104710 157428 104716 157480
rect 104768 157468 104774 157480
rect 189626 157468 189632 157480
rect 104768 157440 189632 157468
rect 104768 157428 104774 157440
rect 189626 157428 189632 157440
rect 189684 157428 189690 157480
rect 119430 157360 119436 157412
rect 119488 157400 119494 157412
rect 511534 157400 511540 157412
rect 119488 157372 511540 157400
rect 119488 157360 119494 157372
rect 511534 157360 511540 157372
rect 511592 157360 511598 157412
rect 73522 157292 73528 157344
rect 73580 157332 73586 157344
rect 168742 157332 168748 157344
rect 73580 157304 168748 157332
rect 73580 157292 73586 157304
rect 168742 157292 168748 157304
rect 168800 157292 168806 157344
rect 175829 157335 175887 157341
rect 175829 157301 175841 157335
rect 175875 157332 175887 157335
rect 181070 157332 181076 157344
rect 175875 157304 181076 157332
rect 175875 157301 175887 157304
rect 175829 157295 175887 157301
rect 181070 157292 181076 157304
rect 181128 157292 181134 157344
rect 189534 157292 189540 157344
rect 189592 157332 189598 157344
rect 246114 157332 246120 157344
rect 189592 157304 246120 157332
rect 189592 157292 189598 157304
rect 246114 157292 246120 157304
rect 246172 157292 246178 157344
rect 426250 157292 426256 157344
rect 426308 157332 426314 157344
rect 458542 157332 458548 157344
rect 426308 157304 458548 157332
rect 426308 157292 426314 157304
rect 458542 157292 458548 157304
rect 458600 157292 458606 157344
rect 475010 157292 475016 157344
rect 475068 157332 475074 157344
rect 485133 157335 485191 157341
rect 475068 157304 485084 157332
rect 475068 157292 475074 157304
rect 68646 157224 68652 157276
rect 68704 157264 68710 157276
rect 165614 157264 165620 157276
rect 68704 157236 165620 157264
rect 68704 157224 68710 157236
rect 165614 157224 165620 157236
rect 165672 157224 165678 157276
rect 165985 157267 166043 157273
rect 165985 157233 165997 157267
rect 166031 157264 166043 157267
rect 170674 157264 170680 157276
rect 166031 157236 170680 157264
rect 166031 157233 166043 157236
rect 165985 157227 166043 157233
rect 170674 157224 170680 157236
rect 170732 157224 170738 157276
rect 172701 157267 172759 157273
rect 172701 157233 172713 157267
rect 172747 157264 172759 157267
rect 172747 157236 175872 157264
rect 172747 157233 172759 157236
rect 172701 157227 172759 157233
rect 65702 157156 65708 157208
rect 65760 157196 65766 157208
rect 163498 157196 163504 157208
rect 65760 157168 163504 157196
rect 65760 157156 65766 157168
rect 163498 157156 163504 157168
rect 163556 157156 163562 157208
rect 167086 157156 167092 157208
rect 167144 157196 167150 157208
rect 173437 157199 173495 157205
rect 173437 157196 173449 157199
rect 167144 157168 173449 157196
rect 167144 157156 167150 157168
rect 173437 157165 173449 157168
rect 173483 157165 173495 157199
rect 175844 157196 175872 157236
rect 175918 157224 175924 157276
rect 175976 157264 175982 157276
rect 237006 157264 237012 157276
rect 175976 157236 237012 157264
rect 175976 157224 175982 157236
rect 237006 157224 237012 157236
rect 237064 157224 237070 157276
rect 428918 157224 428924 157276
rect 428976 157264 428982 157276
rect 462498 157264 462504 157276
rect 428976 157236 462504 157264
rect 428976 157224 428982 157236
rect 462498 157224 462504 157236
rect 462556 157224 462562 157276
rect 473722 157224 473728 157276
rect 473780 157264 473786 157276
rect 473780 157236 476252 157264
rect 473780 157224 473786 157236
rect 176010 157196 176016 157208
rect 175844 157168 176016 157196
rect 173437 157159 173495 157165
rect 176010 157156 176016 157168
rect 176068 157156 176074 157208
rect 177850 157156 177856 157208
rect 177908 157196 177914 157208
rect 238386 157196 238392 157208
rect 177908 157168 238392 157196
rect 177908 157156 177914 157168
rect 238386 157156 238392 157168
rect 238444 157156 238450 157208
rect 436646 157156 436652 157208
rect 436704 157196 436710 157208
rect 474182 157196 474188 157208
rect 436704 157168 474188 157196
rect 436704 157156 436710 157168
rect 474182 157156 474188 157168
rect 474240 157156 474246 157208
rect 57974 157088 57980 157140
rect 58032 157128 58038 157140
rect 158438 157128 158444 157140
rect 58032 157100 158444 157128
rect 58032 157088 58038 157100
rect 158438 157088 158444 157100
rect 158496 157088 158502 157140
rect 163038 157088 163044 157140
rect 163096 157128 163102 157140
rect 173805 157131 173863 157137
rect 173805 157128 173817 157131
rect 163096 157100 173817 157128
rect 163096 157088 163102 157100
rect 173805 157097 173817 157100
rect 173851 157097 173863 157131
rect 173805 157091 173863 157097
rect 173894 157088 173900 157140
rect 173952 157128 173958 157140
rect 235994 157128 236000 157140
rect 173952 157100 236000 157128
rect 173952 157088 173958 157100
rect 235994 157088 236000 157100
rect 236052 157088 236058 157140
rect 251910 157088 251916 157140
rect 251968 157128 251974 157140
rect 287790 157128 287796 157140
rect 251968 157100 287796 157128
rect 251968 157088 251974 157100
rect 287790 157088 287796 157100
rect 287848 157088 287854 157140
rect 438026 157088 438032 157140
rect 438084 157128 438090 157140
rect 476114 157128 476120 157140
rect 438084 157100 476120 157128
rect 438084 157088 438090 157100
rect 476114 157088 476120 157100
rect 476172 157088 476178 157140
rect 56962 157020 56968 157072
rect 57020 157060 57026 157072
rect 157702 157060 157708 157072
rect 57020 157032 157708 157060
rect 57020 157020 57026 157032
rect 157702 157020 157708 157032
rect 157760 157020 157766 157072
rect 160094 157020 160100 157072
rect 160152 157060 160158 157072
rect 166077 157063 166135 157069
rect 166077 157060 166089 157063
rect 160152 157032 166089 157060
rect 160152 157020 160158 157032
rect 166077 157029 166089 157032
rect 166123 157029 166135 157063
rect 166077 157023 166135 157029
rect 166166 157020 166172 157072
rect 166224 157060 166230 157072
rect 230566 157060 230572 157072
rect 166224 157032 230572 157060
rect 166224 157020 166230 157032
rect 230566 157020 230572 157032
rect 230624 157020 230630 157072
rect 244090 157020 244096 157072
rect 244148 157060 244154 157072
rect 282546 157060 282552 157072
rect 244148 157032 282552 157060
rect 244148 157020 244154 157032
rect 282546 157020 282552 157032
rect 282604 157020 282610 157072
rect 437382 157020 437388 157072
rect 437440 157060 437446 157072
rect 475102 157060 475108 157072
rect 437440 157032 475108 157060
rect 437440 157020 437446 157032
rect 475102 157020 475108 157032
rect 475160 157020 475166 157072
rect 476224 157060 476252 157236
rect 477310 157224 477316 157276
rect 477368 157264 477374 157276
rect 485056 157264 485084 157304
rect 485133 157301 485145 157335
rect 485179 157332 485191 157335
rect 529750 157332 529756 157344
rect 485179 157304 529756 157332
rect 485179 157301 485191 157304
rect 485133 157295 485191 157301
rect 529750 157292 529756 157304
rect 529808 157292 529814 157344
rect 531682 157264 531688 157276
rect 477368 157236 484992 157264
rect 485056 157236 531688 157264
rect 477368 157224 477374 157236
rect 484964 157196 484992 157236
rect 531682 157224 531688 157236
rect 531740 157224 531746 157276
rect 535546 157196 535552 157208
rect 484964 157168 535552 157196
rect 535546 157156 535552 157168
rect 535604 157156 535610 157208
rect 478782 157088 478788 157140
rect 478840 157128 478846 157140
rect 537478 157128 537484 157140
rect 478840 157100 537484 157128
rect 478840 157088 478846 157100
rect 537478 157088 537484 157100
rect 537536 157088 537542 157140
rect 485133 157063 485191 157069
rect 485133 157060 485145 157063
rect 476224 157032 485145 157060
rect 485133 157029 485145 157032
rect 485179 157029 485191 157063
rect 485133 157023 485191 157029
rect 485225 157063 485283 157069
rect 485225 157029 485237 157063
rect 485271 157060 485283 157063
rect 541434 157060 541440 157072
rect 485271 157032 541440 157060
rect 485271 157029 485283 157032
rect 485225 157023 485283 157029
rect 541434 157020 541440 157032
rect 541492 157020 541498 157072
rect 53098 156952 53104 157004
rect 53156 156992 53162 157004
rect 155034 156992 155040 157004
rect 53156 156964 155040 156992
rect 53156 156952 53162 156964
rect 155034 156952 155040 156964
rect 155092 156952 155098 157004
rect 158346 156952 158352 157004
rect 158404 156992 158410 157004
rect 225322 156992 225328 157004
rect 158404 156964 225328 156992
rect 158404 156952 158410 156964
rect 225322 156952 225328 156964
rect 225380 156952 225386 157004
rect 236270 156952 236276 157004
rect 236328 156992 236334 157004
rect 277486 156992 277492 157004
rect 236328 156964 277492 156992
rect 236328 156952 236334 156964
rect 277486 156952 277492 156964
rect 277544 156952 277550 157004
rect 442534 156952 442540 157004
rect 442592 156992 442598 157004
rect 482922 156992 482928 157004
rect 442592 156964 482928 156992
rect 442592 156952 442598 156964
rect 482922 156952 482928 156964
rect 482980 156952 482986 157004
rect 483014 156952 483020 157004
rect 483072 156992 483078 157004
rect 543366 156992 543372 157004
rect 483072 156964 543372 156992
rect 483072 156952 483078 156964
rect 543366 156952 543372 156964
rect 543424 156952 543430 157004
rect 42334 156884 42340 156936
rect 42392 156924 42398 156936
rect 147950 156924 147956 156936
rect 42392 156896 147956 156924
rect 42392 156884 42398 156896
rect 147950 156884 147956 156896
rect 148008 156884 148014 156936
rect 150526 156884 150532 156936
rect 150584 156924 150590 156936
rect 220078 156924 220084 156936
rect 150584 156896 220084 156924
rect 150584 156884 150590 156896
rect 220078 156884 220084 156896
rect 220136 156884 220142 156936
rect 228542 156884 228548 156936
rect 228600 156924 228606 156936
rect 272150 156924 272156 156936
rect 228600 156896 272156 156924
rect 228600 156884 228606 156896
rect 272150 156884 272156 156896
rect 272208 156884 272214 156936
rect 442810 156884 442816 156936
rect 442868 156924 442874 156936
rect 483934 156924 483940 156936
rect 442868 156896 483940 156924
rect 442868 156884 442874 156896
rect 483934 156884 483940 156896
rect 483992 156884 483998 156936
rect 485498 156884 485504 156936
rect 485556 156924 485562 156936
rect 547230 156924 547236 156936
rect 485556 156896 547236 156924
rect 485556 156884 485562 156896
rect 547230 156884 547236 156896
rect 547288 156884 547294 156936
rect 25774 156816 25780 156868
rect 25832 156856 25838 156868
rect 136818 156856 136824 156868
rect 25832 156828 136824 156856
rect 25832 156816 25838 156828
rect 136818 156816 136824 156828
rect 136876 156816 136882 156868
rect 139854 156816 139860 156868
rect 139912 156856 139918 156868
rect 212994 156856 213000 156868
rect 139912 156828 213000 156856
rect 139912 156816 139918 156828
rect 212994 156816 213000 156828
rect 213052 156816 213058 156868
rect 218790 156816 218796 156868
rect 218848 156856 218854 156868
rect 265618 156856 265624 156868
rect 218848 156828 265624 156856
rect 218848 156816 218854 156828
rect 265618 156816 265624 156828
rect 265676 156816 265682 156868
rect 445110 156816 445116 156868
rect 445168 156856 445174 156868
rect 486786 156856 486792 156868
rect 445168 156828 486792 156856
rect 445168 156816 445174 156828
rect 486786 156816 486792 156828
rect 486844 156816 486850 156868
rect 486878 156816 486884 156868
rect 486936 156856 486942 156868
rect 549162 156856 549168 156868
rect 486936 156828 549168 156856
rect 486936 156816 486942 156828
rect 549162 156816 549168 156828
rect 549220 156816 549226 156868
rect 17954 156748 17960 156800
rect 18012 156788 18018 156800
rect 131666 156788 131672 156800
rect 18012 156760 131672 156788
rect 18012 156748 18018 156760
rect 131666 156748 131672 156760
rect 131724 156748 131730 156800
rect 134978 156748 134984 156800
rect 135036 156788 135042 156800
rect 209866 156788 209872 156800
rect 135036 156760 209872 156788
rect 135036 156748 135042 156760
rect 209866 156748 209872 156760
rect 209924 156748 209930 156800
rect 212353 156791 212411 156797
rect 212353 156757 212365 156791
rect 212399 156788 212411 156791
rect 218146 156788 218152 156800
rect 212399 156760 218152 156788
rect 212399 156757 212411 156760
rect 212353 156751 212411 156757
rect 218146 156748 218152 156760
rect 218204 156748 218210 156800
rect 221734 156748 221740 156800
rect 221792 156788 221798 156800
rect 267826 156788 267832 156800
rect 221792 156760 267832 156788
rect 221792 156748 221798 156760
rect 267826 156748 267832 156760
rect 267884 156748 267890 156800
rect 445662 156748 445668 156800
rect 445720 156788 445726 156800
rect 487798 156788 487804 156800
rect 445720 156760 487804 156788
rect 445720 156748 445726 156760
rect 487798 156748 487804 156760
rect 487856 156748 487862 156800
rect 490650 156748 490656 156800
rect 490708 156788 490714 156800
rect 555050 156788 555056 156800
rect 490708 156760 555056 156788
rect 490708 156748 490714 156760
rect 555050 156748 555056 156760
rect 555108 156748 555114 156800
rect 10134 156680 10140 156732
rect 10192 156720 10198 156732
rect 126422 156720 126428 156732
rect 10192 156692 126428 156720
rect 10192 156680 10198 156692
rect 126422 156680 126428 156692
rect 126480 156680 126486 156732
rect 132034 156680 132040 156732
rect 132092 156720 132098 156732
rect 207750 156720 207756 156732
rect 132092 156692 207756 156720
rect 132092 156680 132098 156692
rect 207750 156680 207756 156692
rect 207808 156680 207814 156732
rect 212902 156680 212908 156732
rect 212960 156720 212966 156732
rect 261754 156720 261760 156732
rect 212960 156692 261760 156720
rect 212960 156680 212966 156692
rect 261754 156680 261760 156692
rect 261812 156680 261818 156732
rect 449066 156680 449072 156732
rect 449124 156720 449130 156732
rect 492674 156720 492680 156732
rect 449124 156692 492680 156720
rect 449124 156680 449130 156692
rect 492674 156680 492680 156692
rect 492732 156680 492738 156732
rect 493318 156680 493324 156732
rect 493376 156720 493382 156732
rect 558914 156720 558920 156732
rect 493376 156692 558920 156720
rect 493376 156680 493382 156692
rect 558914 156680 558920 156692
rect 558972 156680 558978 156732
rect 6270 156612 6276 156664
rect 6328 156652 6334 156664
rect 123846 156652 123852 156664
rect 6328 156624 123852 156652
rect 6328 156612 6334 156624
rect 123846 156612 123852 156624
rect 123904 156612 123910 156664
rect 124214 156612 124220 156664
rect 124272 156652 124278 156664
rect 202506 156652 202512 156664
rect 124272 156624 202512 156652
rect 124272 156612 124278 156624
rect 202506 156612 202512 156624
rect 202564 156612 202570 156664
rect 209038 156612 209044 156664
rect 209096 156652 209102 156664
rect 259086 156652 259092 156664
rect 209096 156624 259092 156652
rect 209096 156612 209102 156624
rect 259086 156612 259092 156624
rect 259144 156612 259150 156664
rect 420730 156612 420736 156664
rect 420788 156652 420794 156664
rect 450722 156652 450728 156664
rect 420788 156624 450728 156652
rect 420788 156612 420794 156624
rect 450722 156612 450728 156624
rect 450780 156612 450786 156664
rect 456702 156612 456708 156664
rect 456760 156652 456766 156664
rect 504358 156652 504364 156664
rect 456760 156624 504364 156652
rect 456760 156612 456766 156624
rect 504358 156612 504364 156624
rect 504416 156612 504422 156664
rect 508774 156612 508780 156664
rect 508832 156652 508838 156664
rect 577498 156652 577504 156664
rect 508832 156624 577504 156652
rect 508832 156612 508838 156624
rect 577498 156612 577504 156624
rect 577556 156612 577562 156664
rect 76466 156544 76472 156596
rect 76524 156584 76530 156596
rect 165985 156587 166043 156593
rect 165985 156584 165997 156587
rect 76524 156556 165997 156584
rect 76524 156544 76530 156556
rect 165985 156553 165997 156556
rect 166031 156553 166043 156587
rect 165985 156547 166043 156553
rect 166077 156587 166135 156593
rect 166077 156553 166089 156587
rect 166123 156584 166135 156587
rect 223574 156584 223580 156596
rect 166123 156556 223580 156584
rect 166123 156553 166135 156556
rect 166077 156547 166135 156553
rect 223574 156544 223580 156556
rect 223632 156544 223638 156596
rect 469858 156544 469864 156596
rect 469916 156584 469922 156596
rect 523862 156584 523868 156596
rect 469916 156556 523868 156584
rect 469916 156544 469922 156556
rect 523862 156544 523868 156556
rect 523920 156544 523926 156596
rect 81342 156476 81348 156528
rect 81400 156516 81406 156528
rect 173437 156519 173495 156525
rect 81400 156488 172836 156516
rect 81400 156476 81406 156488
rect 84286 156408 84292 156460
rect 84344 156448 84350 156460
rect 172701 156451 172759 156457
rect 172701 156448 172713 156451
rect 84344 156420 172713 156448
rect 84344 156408 84350 156420
rect 172701 156417 172713 156420
rect 172747 156417 172759 156451
rect 172808 156448 172836 156488
rect 173437 156485 173449 156519
rect 173483 156516 173495 156519
rect 231118 156516 231124 156528
rect 173483 156488 231124 156516
rect 173483 156485 173495 156488
rect 173437 156479 173495 156485
rect 231118 156476 231124 156488
rect 231176 156476 231182 156528
rect 465994 156476 466000 156528
rect 466052 156516 466058 156528
rect 517974 156516 517980 156528
rect 466052 156488 517980 156516
rect 466052 156476 466058 156488
rect 517974 156476 517980 156488
rect 518032 156476 518038 156528
rect 173710 156448 173716 156460
rect 172808 156420 173716 156448
rect 172701 156411 172759 156417
rect 173710 156408 173716 156420
rect 173768 156408 173774 156460
rect 173805 156451 173863 156457
rect 173805 156417 173817 156451
rect 173851 156448 173863 156451
rect 225966 156448 225972 156460
rect 173851 156420 225972 156448
rect 173851 156417 173863 156420
rect 173805 156411 173863 156417
rect 225966 156408 225972 156420
rect 226024 156408 226030 156460
rect 440602 156408 440608 156460
rect 440660 156448 440666 156460
rect 479978 156448 479984 156460
rect 440660 156420 479984 156448
rect 440660 156408 440666 156420
rect 479978 156408 479984 156420
rect 480036 156408 480042 156460
rect 480070 156408 480076 156460
rect 480128 156448 480134 156460
rect 530670 156448 530676 156460
rect 480128 156420 530676 156448
rect 480128 156408 480134 156420
rect 530670 156408 530676 156420
rect 530728 156408 530734 156460
rect 92014 156340 92020 156392
rect 92072 156380 92078 156392
rect 175829 156383 175887 156389
rect 175829 156380 175841 156383
rect 92072 156352 175841 156380
rect 92072 156340 92078 156352
rect 175829 156349 175841 156352
rect 175875 156349 175887 156383
rect 175829 156343 175887 156349
rect 178770 156340 178776 156392
rect 178828 156380 178834 156392
rect 180797 156383 180855 156389
rect 180797 156380 180809 156383
rect 178828 156352 180809 156380
rect 178828 156340 178834 156352
rect 180797 156349 180809 156352
rect 180843 156349 180855 156383
rect 180797 156343 180855 156349
rect 180886 156340 180892 156392
rect 180944 156380 180950 156392
rect 191558 156380 191564 156392
rect 180944 156352 191564 156380
rect 180944 156340 180950 156352
rect 191558 156340 191564 156352
rect 191616 156340 191622 156392
rect 193398 156340 193404 156392
rect 193456 156380 193462 156392
rect 248690 156380 248696 156392
rect 193456 156352 248696 156380
rect 193456 156340 193462 156352
rect 248690 156340 248696 156352
rect 248748 156340 248754 156392
rect 481542 156340 481548 156392
rect 481600 156380 481606 156392
rect 485225 156383 485283 156389
rect 485225 156380 485237 156383
rect 481600 156352 485237 156380
rect 481600 156340 481606 156352
rect 485225 156349 485237 156352
rect 485271 156349 485283 156383
rect 485225 156343 485283 156349
rect 487154 156340 487160 156392
rect 487212 156380 487218 156392
rect 538490 156380 538496 156392
rect 487212 156352 538496 156380
rect 487212 156340 487218 156352
rect 538490 156340 538496 156352
rect 538548 156340 538554 156392
rect 99834 156272 99840 156324
rect 99892 156312 99898 156324
rect 186498 156312 186504 156324
rect 99892 156284 186504 156312
rect 99892 156272 99898 156284
rect 186498 156272 186504 156284
rect 186556 156272 186562 156324
rect 191469 156315 191527 156321
rect 191469 156281 191481 156315
rect 191515 156312 191527 156315
rect 197173 156315 197231 156321
rect 197173 156312 197185 156315
rect 191515 156284 197185 156312
rect 191515 156281 191527 156284
rect 191469 156275 191527 156281
rect 197173 156281 197185 156284
rect 197219 156281 197231 156315
rect 197173 156275 197231 156281
rect 197354 156272 197360 156324
rect 197412 156312 197418 156324
rect 251358 156312 251364 156324
rect 197412 156284 251364 156312
rect 197412 156272 197418 156284
rect 251358 156272 251364 156284
rect 251416 156272 251422 156324
rect 460658 156272 460664 156324
rect 460716 156312 460722 156324
rect 510246 156312 510252 156324
rect 460716 156284 510252 156312
rect 460716 156272 460722 156284
rect 510246 156272 510252 156284
rect 510304 156272 510310 156324
rect 107654 156204 107660 156256
rect 107712 156244 107718 156256
rect 180886 156244 180892 156256
rect 107712 156216 180892 156244
rect 107712 156204 107718 156216
rect 180886 156204 180892 156216
rect 180944 156204 180950 156256
rect 180981 156247 181039 156253
rect 180981 156213 180993 156247
rect 181027 156244 181039 156247
rect 183373 156247 183431 156253
rect 183373 156244 183385 156247
rect 181027 156216 183385 156244
rect 181027 156213 181039 156216
rect 180981 156207 181039 156213
rect 183373 156213 183385 156216
rect 183419 156213 183431 156247
rect 183373 156207 183431 156213
rect 183462 156204 183468 156256
rect 183520 156244 183526 156256
rect 236362 156244 236368 156256
rect 183520 156216 236368 156244
rect 183520 156204 183526 156216
rect 236362 156204 236368 156216
rect 236420 156204 236426 156256
rect 453574 156204 453580 156256
rect 453632 156244 453638 156256
rect 499482 156244 499488 156256
rect 453632 156216 499488 156244
rect 453632 156204 453638 156216
rect 499482 156204 499488 156216
rect 499540 156204 499546 156256
rect 111518 156136 111524 156188
rect 111576 156176 111582 156188
rect 111576 156148 191696 156176
rect 111576 156136 111582 156148
rect 116394 156068 116400 156120
rect 116452 156108 116458 156120
rect 191668 156108 191696 156148
rect 191742 156136 191748 156188
rect 191800 156176 191806 156188
rect 241606 156176 241612 156188
rect 191800 156148 241612 156176
rect 191800 156136 191806 156148
rect 241606 156136 241612 156148
rect 241664 156136 241670 156188
rect 452286 156136 452292 156188
rect 452344 156176 452350 156188
rect 497550 156176 497556 156188
rect 452344 156148 497556 156176
rect 452344 156136 452350 156148
rect 497550 156136 497556 156148
rect 497608 156136 497614 156188
rect 194042 156108 194048 156120
rect 116452 156080 191604 156108
rect 191668 156080 194048 156108
rect 116452 156068 116458 156080
rect 119338 156000 119344 156052
rect 119396 156040 119402 156052
rect 191469 156043 191527 156049
rect 191469 156040 191481 156043
rect 119396 156012 191481 156040
rect 119396 156000 119402 156012
rect 191469 156009 191481 156012
rect 191515 156009 191527 156043
rect 191576 156040 191604 156080
rect 194042 156068 194048 156080
rect 194100 156068 194106 156120
rect 197173 156111 197231 156117
rect 197173 156077 197185 156111
rect 197219 156108 197231 156111
rect 199378 156108 199384 156120
rect 197219 156080 199384 156108
rect 197219 156077 197231 156080
rect 197173 156071 197231 156077
rect 199378 156068 199384 156080
rect 199436 156068 199442 156120
rect 200025 156111 200083 156117
rect 200025 156077 200037 156111
rect 200071 156108 200083 156111
rect 244366 156108 244372 156120
rect 200071 156080 244372 156108
rect 200071 156077 200083 156080
rect 200025 156071 200083 156077
rect 244366 156068 244372 156080
rect 244424 156068 244430 156120
rect 450354 156068 450360 156120
rect 450412 156108 450418 156120
rect 494606 156108 494612 156120
rect 450412 156080 494612 156108
rect 450412 156068 450418 156080
rect 494606 156068 494612 156080
rect 494664 156068 494670 156120
rect 197446 156040 197452 156052
rect 191576 156012 197452 156040
rect 191469 156003 191527 156009
rect 197446 156000 197452 156012
rect 197504 156000 197510 156052
rect 205634 156000 205640 156052
rect 205692 156040 205698 156052
rect 214285 156043 214343 156049
rect 205692 156012 214236 156040
rect 205692 156000 205698 156012
rect 155862 155932 155868 155984
rect 155920 155972 155926 155984
rect 212353 155975 212411 155981
rect 212353 155972 212365 155975
rect 155920 155944 212365 155972
rect 155920 155932 155926 155944
rect 212353 155941 212365 155944
rect 212399 155941 212411 155975
rect 214009 155975 214067 155981
rect 214009 155972 214021 155975
rect 212353 155935 212411 155941
rect 212460 155944 214021 155972
rect 12158 155864 12164 155916
rect 12216 155904 12222 155916
rect 12216 155876 16574 155904
rect 12216 155864 12222 155876
rect 4338 155796 4344 155848
rect 4396 155836 4402 155848
rect 12434 155836 12440 155848
rect 4396 155808 12440 155836
rect 4396 155796 4402 155808
rect 12434 155796 12440 155808
rect 12492 155796 12498 155848
rect 16546 155836 16574 155876
rect 33594 155864 33600 155916
rect 33652 155904 33658 155916
rect 34698 155904 34704 155916
rect 33652 155876 34704 155904
rect 33652 155864 33658 155876
rect 34698 155864 34704 155876
rect 34756 155864 34762 155916
rect 66714 155864 66720 155916
rect 66772 155904 66778 155916
rect 82814 155904 82820 155916
rect 66772 155876 82820 155904
rect 66772 155864 66778 155876
rect 82814 155864 82820 155876
rect 82872 155864 82878 155916
rect 108301 155907 108359 155913
rect 108301 155873 108313 155907
rect 108347 155904 108359 155907
rect 175921 155907 175979 155913
rect 175921 155904 175933 155907
rect 108347 155876 175933 155904
rect 108347 155873 108359 155876
rect 108301 155867 108359 155873
rect 175921 155873 175933 155876
rect 175967 155873 175979 155907
rect 175921 155867 175979 155873
rect 176838 155864 176844 155916
rect 176896 155904 176902 155916
rect 179138 155904 179144 155916
rect 176896 155876 179144 155904
rect 176896 155864 176902 155876
rect 179138 155864 179144 155876
rect 179196 155864 179202 155916
rect 180794 155864 180800 155916
rect 180852 155904 180858 155916
rect 183370 155904 183376 155916
rect 180852 155876 183376 155904
rect 180852 155864 180858 155876
rect 183370 155864 183376 155876
rect 183428 155864 183434 155916
rect 183465 155907 183523 155913
rect 183465 155873 183477 155907
rect 183511 155904 183523 155907
rect 185305 155907 185363 155913
rect 185305 155904 185317 155907
rect 183511 155876 185317 155904
rect 183511 155873 183523 155876
rect 183465 155867 183523 155873
rect 185305 155873 185317 155876
rect 185351 155873 185363 155907
rect 186406 155904 186412 155916
rect 185305 155867 185363 155873
rect 185412 155876 186412 155904
rect 17862 155836 17868 155848
rect 16546 155808 17868 155836
rect 17862 155796 17868 155808
rect 17920 155796 17926 155848
rect 43346 155796 43352 155848
rect 43404 155836 43410 155848
rect 51074 155836 51080 155848
rect 43404 155808 51080 155836
rect 43404 155796 43410 155808
rect 51074 155796 51080 155808
rect 51132 155796 51138 155848
rect 63770 155796 63776 155848
rect 63828 155836 63834 155848
rect 137281 155839 137339 155845
rect 137281 155836 137293 155839
rect 63828 155808 137293 155836
rect 63828 155796 63834 155808
rect 137281 155805 137293 155808
rect 137327 155805 137339 155839
rect 185412 155836 185440 155876
rect 186406 155864 186412 155876
rect 186464 155864 186470 155916
rect 186590 155864 186596 155916
rect 186648 155904 186654 155916
rect 200025 155907 200083 155913
rect 200025 155904 200037 155907
rect 186648 155876 200037 155904
rect 186648 155864 186654 155876
rect 200025 155873 200037 155876
rect 200071 155873 200083 155907
rect 200025 155867 200083 155873
rect 200206 155864 200212 155916
rect 200264 155904 200270 155916
rect 202782 155904 202788 155916
rect 200264 155876 202788 155904
rect 200264 155864 200270 155876
rect 202782 155864 202788 155876
rect 202840 155864 202846 155916
rect 206094 155864 206100 155916
rect 206152 155904 206158 155916
rect 212460 155904 212488 155944
rect 214009 155941 214021 155944
rect 214055 155941 214067 155975
rect 214208 155972 214236 156012
rect 214285 156009 214297 156043
rect 214331 156040 214343 156043
rect 257154 156040 257160 156052
rect 214331 156012 257160 156040
rect 214331 156009 214343 156012
rect 214285 156003 214343 156009
rect 257154 156000 257160 156012
rect 257212 156000 257218 156052
rect 446490 156000 446496 156052
rect 446548 156040 446554 156052
rect 488810 156040 488816 156052
rect 446548 156012 488816 156040
rect 446548 156000 446554 156012
rect 488810 156000 488816 156012
rect 488868 156000 488874 156052
rect 249334 155972 249340 155984
rect 214208 155944 249340 155972
rect 214009 155935 214067 155941
rect 249334 155932 249340 155944
rect 249392 155932 249398 155984
rect 262861 155975 262919 155981
rect 262861 155972 262873 155975
rect 258644 155944 262873 155972
rect 206152 155876 212488 155904
rect 206152 155864 206158 155876
rect 215846 155864 215852 155916
rect 215904 155904 215910 155916
rect 216582 155904 216588 155916
rect 215904 155876 216588 155904
rect 215904 155864 215910 155876
rect 216582 155864 216588 155876
rect 216640 155864 216646 155916
rect 219621 155907 219679 155913
rect 219621 155873 219633 155907
rect 219667 155904 219679 155907
rect 219667 155876 222516 155904
rect 219667 155873 219679 155876
rect 219621 155867 219679 155873
rect 137281 155799 137339 155805
rect 142126 155808 185440 155836
rect 185489 155839 185547 155845
rect 55950 155728 55956 155780
rect 56008 155768 56014 155780
rect 136821 155771 136879 155777
rect 136821 155768 136833 155771
rect 56008 155740 136833 155768
rect 56008 155728 56014 155740
rect 136821 155737 136833 155740
rect 136867 155737 136879 155771
rect 136821 155731 136879 155737
rect 136910 155728 136916 155780
rect 136968 155768 136974 155780
rect 142126 155768 142154 155808
rect 185489 155805 185501 155839
rect 185535 155836 185547 155839
rect 222381 155839 222439 155845
rect 222381 155836 222393 155839
rect 185535 155808 222393 155836
rect 185535 155805 185547 155808
rect 185489 155799 185547 155805
rect 222381 155805 222393 155808
rect 222427 155805 222439 155839
rect 222381 155799 222439 155805
rect 136968 155740 142154 155768
rect 136968 155728 136974 155740
rect 143718 155728 143724 155780
rect 143776 155768 143782 155780
rect 144638 155768 144644 155780
rect 143776 155740 144644 155768
rect 143776 155728 143782 155740
rect 144638 155728 144644 155740
rect 144696 155728 144702 155780
rect 144730 155728 144736 155780
rect 144788 155768 144794 155780
rect 148229 155771 148287 155777
rect 148229 155768 148241 155771
rect 144788 155740 148241 155768
rect 144788 155728 144794 155740
rect 148229 155737 148241 155740
rect 148275 155737 148287 155771
rect 148229 155731 148287 155737
rect 149606 155728 149612 155780
rect 149664 155768 149670 155780
rect 153102 155768 153108 155780
rect 149664 155740 153108 155768
rect 149664 155728 149670 155740
rect 153102 155728 153108 155740
rect 153160 155728 153166 155780
rect 153470 155728 153476 155780
rect 153528 155768 153534 155780
rect 155313 155771 155371 155777
rect 155313 155768 155325 155771
rect 153528 155740 155325 155768
rect 153528 155728 153534 155740
rect 155313 155737 155325 155740
rect 155359 155737 155371 155771
rect 155313 155731 155371 155737
rect 155402 155728 155408 155780
rect 155460 155768 155466 155780
rect 160094 155768 160100 155780
rect 155460 155740 160100 155768
rect 155460 155728 155466 155740
rect 160094 155728 160100 155740
rect 160152 155728 160158 155780
rect 160278 155728 160284 155780
rect 160336 155768 160342 155780
rect 166261 155771 166319 155777
rect 166261 155768 166273 155771
rect 160336 155740 166273 155768
rect 160336 155728 160342 155740
rect 166261 155737 166273 155740
rect 166307 155737 166319 155771
rect 172146 155768 172152 155780
rect 166261 155731 166319 155737
rect 171888 155740 172152 155768
rect 74534 155660 74540 155712
rect 74592 155700 74598 155712
rect 167730 155700 167736 155712
rect 74592 155672 167736 155700
rect 74592 155660 74598 155672
rect 167730 155660 167736 155672
rect 167788 155660 167794 155712
rect 171042 155660 171048 155712
rect 171100 155700 171106 155712
rect 171888 155700 171916 155740
rect 172146 155728 172152 155740
rect 172204 155728 172210 155780
rect 172241 155771 172299 155777
rect 172241 155737 172253 155771
rect 172287 155768 172299 155771
rect 219621 155771 219679 155777
rect 219621 155768 219633 155771
rect 172287 155740 219633 155768
rect 172287 155737 172299 155740
rect 172241 155731 172299 155737
rect 219621 155737 219633 155740
rect 219667 155737 219679 155771
rect 219621 155731 219679 155737
rect 219710 155728 219716 155780
rect 219768 155768 219774 155780
rect 222102 155768 222108 155780
rect 219768 155740 222108 155768
rect 219768 155728 219774 155740
rect 222102 155728 222108 155740
rect 222160 155728 222166 155780
rect 222488 155768 222516 155876
rect 222654 155864 222660 155916
rect 222712 155904 222718 155916
rect 258644 155904 258672 155944
rect 262861 155941 262873 155944
rect 262907 155941 262919 155975
rect 262861 155935 262919 155941
rect 287793 155975 287851 155981
rect 287793 155941 287805 155975
rect 287839 155972 287851 155975
rect 289357 155975 289415 155981
rect 289357 155972 289369 155975
rect 287839 155944 289369 155972
rect 287839 155941 287851 155944
rect 287793 155935 287851 155941
rect 289357 155941 289369 155944
rect 289403 155941 289415 155975
rect 296809 155975 296867 155981
rect 296809 155972 296821 155975
rect 289357 155935 289415 155941
rect 296548 155944 296821 155972
rect 222712 155876 258672 155904
rect 222712 155864 222718 155876
rect 258718 155864 258724 155916
rect 258776 155904 258782 155916
rect 262122 155904 262128 155916
rect 258776 155876 262128 155904
rect 258776 155864 258782 155876
rect 262122 155864 262128 155876
rect 262180 155864 262186 155916
rect 262677 155907 262735 155913
rect 262677 155873 262689 155907
rect 262723 155904 262735 155907
rect 277857 155907 277915 155913
rect 277857 155904 277869 155907
rect 262723 155876 277869 155904
rect 262723 155873 262735 155876
rect 262677 155867 262735 155873
rect 277857 155873 277869 155876
rect 277903 155873 277915 155907
rect 280246 155904 280252 155916
rect 277857 155867 277915 155873
rect 277964 155876 280252 155904
rect 222565 155839 222623 155845
rect 222565 155805 222577 155839
rect 222611 155836 222623 155839
rect 229373 155839 229431 155845
rect 229373 155836 229385 155839
rect 222611 155808 229385 155836
rect 222611 155805 222623 155808
rect 222565 155799 222623 155805
rect 229373 155805 229385 155808
rect 229419 155805 229431 155839
rect 229373 155799 229431 155805
rect 229462 155796 229468 155848
rect 229520 155836 229526 155848
rect 239125 155839 239183 155845
rect 229520 155808 238754 155836
rect 229520 155796 229526 155808
rect 225046 155768 225052 155780
rect 222488 155740 225052 155768
rect 225046 155728 225052 155740
rect 225104 155728 225110 155780
rect 225598 155728 225604 155780
rect 225656 155768 225662 155780
rect 233881 155771 233939 155777
rect 233881 155768 233893 155771
rect 225656 155740 233893 155768
rect 225656 155728 225662 155740
rect 233881 155737 233893 155740
rect 233927 155737 233939 155771
rect 238726 155768 238754 155808
rect 239125 155805 239137 155839
rect 239171 155836 239183 155839
rect 241057 155839 241115 155845
rect 241057 155836 241069 155839
rect 239171 155808 241069 155836
rect 239171 155805 239183 155808
rect 239125 155799 239183 155805
rect 241057 155805 241069 155808
rect 241103 155805 241115 155839
rect 241057 155799 241115 155805
rect 241146 155796 241152 155848
rect 241204 155836 241210 155848
rect 248969 155839 249027 155845
rect 248969 155836 248981 155839
rect 241204 155808 248981 155836
rect 241204 155796 241210 155808
rect 248969 155805 248981 155808
rect 249015 155805 249027 155839
rect 277964 155836 277992 155876
rect 280246 155864 280252 155876
rect 280304 155864 280310 155916
rect 280341 155907 280399 155913
rect 280341 155873 280353 155907
rect 280387 155904 280399 155907
rect 280387 155876 284064 155904
rect 280387 155873 280399 155876
rect 280341 155867 280399 155873
rect 248969 155799 249027 155805
rect 249076 155808 277992 155836
rect 278041 155839 278099 155845
rect 248877 155771 248935 155777
rect 248877 155768 248889 155771
rect 238726 155740 248889 155768
rect 233881 155731 233939 155737
rect 248877 155737 248889 155740
rect 248923 155737 248935 155771
rect 248877 155731 248935 155737
rect 171100 155672 171916 155700
rect 171100 155660 171106 155672
rect 171962 155660 171968 155712
rect 172020 155700 172026 155712
rect 233329 155703 233387 155709
rect 233329 155700 233341 155703
rect 172020 155672 233341 155700
rect 172020 155660 172026 155672
rect 233329 155669 233341 155672
rect 233375 155669 233387 155703
rect 233329 155663 233387 155669
rect 233418 155660 233424 155712
rect 233476 155700 233482 155712
rect 243081 155703 243139 155709
rect 243081 155700 243093 155703
rect 233476 155672 243093 155700
rect 233476 155660 233482 155672
rect 243081 155669 243093 155672
rect 243127 155669 243139 155703
rect 243081 155663 243139 155669
rect 243170 155660 243176 155712
rect 243228 155700 243234 155712
rect 249076 155700 249104 155808
rect 278041 155805 278053 155839
rect 278087 155836 278099 155839
rect 281442 155836 281448 155848
rect 278087 155808 281448 155836
rect 278087 155805 278099 155808
rect 278041 155799 278099 155805
rect 281442 155796 281448 155808
rect 281500 155796 281506 155848
rect 284036 155836 284064 155876
rect 284110 155864 284116 155916
rect 284168 155904 284174 155916
rect 291746 155904 291752 155916
rect 284168 155876 291752 155904
rect 284168 155864 284174 155876
rect 291746 155864 291752 155876
rect 291804 155864 291810 155916
rect 292850 155864 292856 155916
rect 292908 155904 292914 155916
rect 296548 155904 296576 155944
rect 296809 155941 296821 155944
rect 296855 155941 296867 155975
rect 296809 155935 296867 155941
rect 447778 155932 447784 155984
rect 447836 155972 447842 155984
rect 490742 155972 490748 155984
rect 447836 155944 490748 155972
rect 447836 155932 447842 155944
rect 490742 155932 490748 155944
rect 490800 155932 490806 155984
rect 292908 155876 296576 155904
rect 296625 155907 296683 155913
rect 292908 155864 292914 155876
rect 296625 155873 296637 155907
rect 296671 155904 296683 155907
rect 313734 155904 313740 155916
rect 296671 155876 313740 155904
rect 296671 155873 296683 155876
rect 296625 155867 296683 155873
rect 313734 155864 313740 155876
rect 313792 155864 313798 155916
rect 316218 155864 316224 155916
rect 316276 155904 316282 155916
rect 328454 155904 328460 155916
rect 316276 155876 328460 155904
rect 316276 155864 316282 155876
rect 328454 155864 328460 155876
rect 328512 155864 328518 155916
rect 328914 155864 328920 155916
rect 328972 155904 328978 155916
rect 334342 155904 334348 155916
rect 328972 155876 334348 155904
rect 328972 155864 328978 155876
rect 334342 155864 334348 155876
rect 334400 155864 334406 155916
rect 334802 155864 334808 155916
rect 334860 155904 334866 155916
rect 340230 155904 340236 155916
rect 334860 155876 340236 155904
rect 334860 155864 334866 155876
rect 340230 155864 340236 155876
rect 340288 155864 340294 155916
rect 353294 155864 353300 155916
rect 353352 155904 353358 155916
rect 355410 155904 355416 155916
rect 353352 155876 355416 155904
rect 353352 155864 353358 155876
rect 355410 155864 355416 155876
rect 355468 155864 355474 155916
rect 382366 155864 382372 155916
rect 382424 155904 382430 155916
rect 385494 155904 385500 155916
rect 382424 155876 385500 155904
rect 382424 155864 382430 155876
rect 385494 155864 385500 155876
rect 385552 155864 385558 155916
rect 388438 155864 388444 155916
rect 388496 155904 388502 155916
rect 393222 155904 393228 155916
rect 388496 155876 393228 155904
rect 388496 155864 388502 155876
rect 393222 155864 393228 155876
rect 393280 155864 393286 155916
rect 404170 155864 404176 155916
rect 404228 155904 404234 155916
rect 406930 155904 406936 155916
rect 404228 155876 406936 155904
rect 404228 155864 404234 155876
rect 406930 155864 406936 155876
rect 406988 155864 406994 155916
rect 407025 155907 407083 155913
rect 407025 155873 407037 155907
rect 407071 155904 407083 155907
rect 426342 155904 426348 155916
rect 407071 155876 426348 155904
rect 407071 155873 407083 155876
rect 407025 155867 407083 155873
rect 426342 155864 426348 155876
rect 426400 155864 426406 155916
rect 457622 155904 457628 155916
rect 426452 155876 457628 155904
rect 284386 155836 284392 155848
rect 284036 155808 284392 155836
rect 284386 155796 284392 155808
rect 284444 155796 284450 155848
rect 286962 155796 286968 155848
rect 287020 155836 287026 155848
rect 311250 155836 311256 155848
rect 287020 155808 311256 155836
rect 287020 155796 287026 155808
rect 311250 155796 311256 155808
rect 311308 155796 311314 155848
rect 315298 155796 315304 155848
rect 315356 155836 315362 155848
rect 329650 155836 329656 155848
rect 315356 155808 329656 155836
rect 315356 155796 315362 155808
rect 329650 155796 329656 155808
rect 329708 155796 329714 155848
rect 330846 155796 330852 155848
rect 330904 155836 330910 155848
rect 336550 155836 336556 155848
rect 330904 155808 336556 155836
rect 330904 155796 330910 155808
rect 336550 155796 336556 155808
rect 336608 155796 336614 155848
rect 354214 155796 354220 155848
rect 354272 155836 354278 155848
rect 355962 155836 355968 155848
rect 354272 155808 355968 155836
rect 354272 155796 354278 155808
rect 355962 155796 355968 155808
rect 356020 155796 356026 155848
rect 387334 155796 387340 155848
rect 387392 155836 387398 155848
rect 391290 155836 391296 155848
rect 387392 155808 391296 155836
rect 387392 155796 387398 155808
rect 391290 155796 391296 155808
rect 391348 155796 391354 155848
rect 402238 155796 402244 155848
rect 402296 155836 402302 155848
rect 422478 155836 422484 155848
rect 402296 155808 422484 155836
rect 402296 155796 402302 155808
rect 422478 155796 422484 155808
rect 422536 155796 422542 155848
rect 424962 155796 424968 155848
rect 425020 155836 425026 155848
rect 425517 155839 425575 155845
rect 425517 155836 425529 155839
rect 425020 155808 425529 155836
rect 425020 155796 425026 155808
rect 425517 155805 425529 155808
rect 425563 155805 425575 155839
rect 425517 155799 425575 155805
rect 425606 155796 425612 155848
rect 425664 155836 425670 155848
rect 426452 155836 426480 155876
rect 457622 155864 457628 155876
rect 457680 155864 457686 155916
rect 466270 155864 466276 155916
rect 466328 155904 466334 155916
rect 518986 155904 518992 155916
rect 466328 155876 518992 155904
rect 466328 155864 466334 155876
rect 518986 155864 518992 155876
rect 519044 155864 519050 155916
rect 546494 155864 546500 155916
rect 546552 155904 546558 155916
rect 548242 155904 548248 155916
rect 546552 155876 548248 155904
rect 546552 155864 546558 155876
rect 548242 155864 548248 155876
rect 548300 155864 548306 155916
rect 425664 155808 426480 155836
rect 426529 155839 426587 155845
rect 425664 155796 425670 155808
rect 426529 155805 426541 155839
rect 426575 155836 426587 155839
rect 428185 155839 428243 155845
rect 428185 155836 428197 155839
rect 426575 155808 428197 155836
rect 426575 155805 426587 155808
rect 426529 155799 426587 155805
rect 428185 155805 428197 155808
rect 428231 155805 428243 155839
rect 428185 155799 428243 155805
rect 428274 155796 428280 155848
rect 428332 155836 428338 155848
rect 428553 155839 428611 155845
rect 428332 155808 428504 155836
rect 428332 155796 428338 155808
rect 249153 155771 249211 155777
rect 249153 155737 249165 155771
rect 249199 155768 249211 155771
rect 262769 155771 262827 155777
rect 262769 155768 262781 155771
rect 249199 155740 262781 155768
rect 249199 155737 249211 155740
rect 249153 155731 249211 155737
rect 262769 155737 262781 155740
rect 262815 155737 262827 155771
rect 262769 155731 262827 155737
rect 262861 155771 262919 155777
rect 262861 155737 262873 155771
rect 262907 155768 262919 155771
rect 263778 155768 263784 155780
rect 262907 155740 263784 155768
rect 262907 155737 262919 155740
rect 262861 155731 262919 155737
rect 263778 155728 263784 155740
rect 263836 155728 263842 155780
rect 264606 155728 264612 155780
rect 264664 155768 264670 155780
rect 268381 155771 268439 155777
rect 268381 155768 268393 155771
rect 264664 155740 268393 155768
rect 264664 155728 264670 155740
rect 268381 155737 268393 155740
rect 268427 155737 268439 155771
rect 268381 155731 268439 155737
rect 268470 155728 268476 155780
rect 268528 155768 268534 155780
rect 268528 155740 278176 155768
rect 268528 155728 268534 155740
rect 278041 155703 278099 155709
rect 278041 155700 278053 155703
rect 243228 155672 249104 155700
rect 249168 155672 278053 155700
rect 243228 155660 243234 155672
rect 39390 155592 39396 155644
rect 39448 155632 39454 155644
rect 133325 155635 133383 155641
rect 133325 155632 133337 155635
rect 39448 155604 133337 155632
rect 39448 155592 39454 155604
rect 133325 155601 133337 155604
rect 133371 155601 133383 155635
rect 133325 155595 133383 155601
rect 133417 155635 133475 155641
rect 133417 155601 133429 155635
rect 133463 155632 133475 155635
rect 182637 155635 182695 155641
rect 182637 155632 182649 155635
rect 133463 155604 182649 155632
rect 133463 155601 133475 155604
rect 133417 155595 133475 155601
rect 182637 155601 182649 155604
rect 182683 155601 182695 155635
rect 182637 155595 182695 155601
rect 182726 155592 182732 155644
rect 182784 155632 182790 155644
rect 187145 155635 187203 155641
rect 187145 155632 187157 155635
rect 182784 155604 187157 155632
rect 182784 155592 182790 155604
rect 187145 155601 187157 155604
rect 187191 155601 187203 155635
rect 187145 155595 187203 155601
rect 191466 155592 191472 155644
rect 191524 155632 191530 155644
rect 239125 155635 239183 155641
rect 239125 155632 239137 155635
rect 191524 155604 239137 155632
rect 191524 155592 191530 155604
rect 239125 155601 239137 155604
rect 239171 155601 239183 155635
rect 239125 155595 239183 155601
rect 239214 155592 239220 155644
rect 239272 155632 239278 155644
rect 241422 155632 241428 155644
rect 239272 155604 241428 155632
rect 239272 155592 239278 155604
rect 241422 155592 241428 155604
rect 241480 155592 241486 155644
rect 243633 155635 243691 155641
rect 243633 155632 243645 155635
rect 242084 155604 243645 155632
rect 16022 155524 16028 155576
rect 16080 155564 16086 155576
rect 117958 155564 117964 155576
rect 16080 155536 117964 155564
rect 16080 155524 16086 155536
rect 117958 155524 117964 155536
rect 118016 155524 118022 155576
rect 118326 155524 118332 155576
rect 118384 155564 118390 155576
rect 127713 155567 127771 155573
rect 127713 155564 127725 155567
rect 118384 155536 127725 155564
rect 118384 155524 118390 155536
rect 127713 155533 127725 155536
rect 127759 155533 127771 155567
rect 127713 155527 127771 155533
rect 127897 155567 127955 155573
rect 127897 155533 127909 155567
rect 127943 155564 127955 155567
rect 185581 155567 185639 155573
rect 185581 155564 185593 155567
rect 127943 155536 185593 155564
rect 127943 155533 127955 155536
rect 127897 155527 127955 155533
rect 185581 155533 185593 155536
rect 185627 155533 185639 155567
rect 185581 155527 185639 155533
rect 185673 155567 185731 155573
rect 185673 155533 185685 155567
rect 185719 155564 185731 155567
rect 187786 155564 187792 155576
rect 185719 155536 187792 155564
rect 185719 155533 185731 155536
rect 185673 155527 185731 155533
rect 187786 155524 187792 155536
rect 187844 155524 187850 155576
rect 190546 155524 190552 155576
rect 190604 155564 190610 155576
rect 195241 155567 195299 155573
rect 195241 155564 195253 155567
rect 190604 155536 195253 155564
rect 190604 155524 190610 155536
rect 195241 155533 195253 155536
rect 195287 155533 195299 155567
rect 195241 155527 195299 155533
rect 195330 155524 195336 155576
rect 195388 155564 195394 155576
rect 242084 155564 242112 155604
rect 243633 155601 243645 155604
rect 243679 155601 243691 155635
rect 243633 155595 243691 155601
rect 245102 155592 245108 155644
rect 245160 155632 245166 155644
rect 249061 155635 249119 155641
rect 249061 155632 249073 155635
rect 245160 155604 249073 155632
rect 245160 155592 245166 155604
rect 249061 155601 249073 155604
rect 249107 155601 249119 155635
rect 249061 155595 249119 155601
rect 195388 155536 242112 155564
rect 195388 155524 195394 155536
rect 242158 155524 242164 155576
rect 242216 155564 242222 155576
rect 249168 155564 249196 155672
rect 278041 155669 278053 155672
rect 278087 155669 278099 155703
rect 278148 155700 278176 155740
rect 278222 155728 278228 155780
rect 278280 155768 278286 155780
rect 296717 155771 296775 155777
rect 296717 155768 296729 155771
rect 278280 155740 296729 155768
rect 278280 155728 278286 155740
rect 296717 155737 296729 155740
rect 296763 155737 296775 155771
rect 296717 155731 296775 155737
rect 296809 155771 296867 155777
rect 296809 155737 296821 155771
rect 296855 155768 296867 155771
rect 304994 155768 305000 155780
rect 296855 155740 305000 155768
rect 296855 155737 296867 155740
rect 296809 155731 296867 155737
rect 304994 155728 305000 155740
rect 305052 155728 305058 155780
rect 305546 155728 305552 155780
rect 305604 155768 305610 155780
rect 323486 155768 323492 155780
rect 305604 155740 323492 155768
rect 305604 155728 305610 155740
rect 323486 155728 323492 155740
rect 323544 155728 323550 155780
rect 331858 155728 331864 155780
rect 331916 155768 331922 155780
rect 337930 155768 337936 155780
rect 331916 155740 337936 155768
rect 331916 155728 331922 155740
rect 337930 155728 337936 155740
rect 337988 155728 337994 155780
rect 385494 155728 385500 155780
rect 385552 155768 385558 155780
rect 390278 155768 390284 155780
rect 385552 155740 390284 155768
rect 385552 155728 385558 155740
rect 390278 155728 390284 155740
rect 390336 155728 390342 155780
rect 405826 155728 405832 155780
rect 405884 155768 405890 155780
rect 409782 155768 409788 155780
rect 405884 155740 409788 155768
rect 405884 155728 405890 155740
rect 409782 155728 409788 155740
rect 409840 155728 409846 155780
rect 411346 155728 411352 155780
rect 411404 155768 411410 155780
rect 412726 155768 412732 155780
rect 411404 155740 412732 155768
rect 411404 155728 411410 155740
rect 412726 155728 412732 155740
rect 412784 155728 412790 155780
rect 413278 155728 413284 155780
rect 413336 155768 413342 155780
rect 414658 155768 414664 155780
rect 413336 155740 414664 155768
rect 413336 155728 413342 155740
rect 414658 155728 414664 155740
rect 414716 155728 414722 155780
rect 417329 155771 417387 155777
rect 417329 155737 417341 155771
rect 417375 155768 417387 155771
rect 428366 155768 428372 155780
rect 417375 155740 428372 155768
rect 417375 155737 417387 155740
rect 417329 155731 417387 155737
rect 428366 155728 428372 155740
rect 428424 155728 428430 155780
rect 428476 155768 428504 155808
rect 428553 155805 428565 155839
rect 428599 155836 428611 155839
rect 456610 155836 456616 155848
rect 428599 155808 456616 155836
rect 428599 155805 428611 155808
rect 428553 155799 428611 155805
rect 456610 155796 456616 155808
rect 456668 155796 456674 155848
rect 469122 155796 469128 155848
rect 469180 155836 469186 155848
rect 522850 155836 522856 155848
rect 469180 155808 522856 155836
rect 469180 155796 469186 155808
rect 522850 155796 522856 155808
rect 522908 155796 522914 155848
rect 461486 155768 461492 155780
rect 428476 155740 461492 155768
rect 461486 155728 461492 155740
rect 461544 155728 461550 155780
rect 471146 155728 471152 155780
rect 471204 155768 471210 155780
rect 525794 155768 525800 155780
rect 471204 155740 525800 155768
rect 471204 155728 471210 155740
rect 525794 155728 525800 155740
rect 525852 155728 525858 155780
rect 282914 155700 282920 155712
rect 278148 155672 282920 155700
rect 278041 155663 278099 155669
rect 282914 155660 282920 155672
rect 282972 155660 282978 155712
rect 283098 155660 283104 155712
rect 283156 155700 283162 155712
rect 301501 155703 301559 155709
rect 301501 155700 301513 155703
rect 283156 155672 301513 155700
rect 283156 155660 283162 155672
rect 301501 155669 301513 155672
rect 301547 155669 301559 155703
rect 301501 155663 301559 155669
rect 301593 155703 301651 155709
rect 301593 155669 301605 155703
rect 301639 155700 301651 155703
rect 305914 155700 305920 155712
rect 301639 155672 305920 155700
rect 301639 155669 301651 155672
rect 301593 155663 301651 155669
rect 305914 155660 305920 155672
rect 305972 155660 305978 155712
rect 307297 155703 307355 155709
rect 307297 155669 307309 155703
rect 307343 155700 307355 155703
rect 313366 155700 313372 155712
rect 307343 155672 313372 155700
rect 307343 155669 307355 155672
rect 307297 155663 307355 155669
rect 313366 155660 313372 155672
rect 313424 155660 313430 155712
rect 314286 155660 314292 155712
rect 314344 155700 314350 155712
rect 329374 155700 329380 155712
rect 314344 155672 329380 155700
rect 314344 155660 314350 155672
rect 329374 155660 329380 155672
rect 329432 155660 329438 155712
rect 404814 155660 404820 155712
rect 404872 155700 404878 155712
rect 407025 155703 407083 155709
rect 407025 155700 407037 155703
rect 404872 155672 407037 155700
rect 404872 155660 404878 155672
rect 407025 155669 407037 155672
rect 407071 155669 407083 155703
rect 407025 155663 407083 155669
rect 411254 155660 411260 155712
rect 411312 155700 411318 155712
rect 413738 155700 413744 155712
rect 411312 155672 413744 155700
rect 411312 155660 411318 155672
rect 413738 155660 413744 155672
rect 413796 155660 413802 155712
rect 414106 155660 414112 155712
rect 414164 155700 414170 155712
rect 416682 155700 416688 155712
rect 414164 155672 416688 155700
rect 414164 155660 414170 155672
rect 416682 155660 416688 155672
rect 416740 155660 416746 155712
rect 417421 155703 417479 155709
rect 417421 155669 417433 155703
rect 417467 155700 417479 155703
rect 430298 155700 430304 155712
rect 417467 155672 430304 155700
rect 417467 155669 417479 155672
rect 417421 155663 417479 155669
rect 430298 155660 430304 155672
rect 430356 155660 430362 155712
rect 430390 155660 430396 155712
rect 430448 155700 430454 155712
rect 464430 155700 464436 155712
rect 430448 155672 464436 155700
rect 430448 155660 430454 155672
rect 464430 155660 464436 155672
rect 464488 155660 464494 155712
rect 475746 155660 475752 155712
rect 475804 155700 475810 155712
rect 532602 155700 532608 155712
rect 475804 155672 532608 155700
rect 475804 155660 475810 155672
rect 532602 155660 532608 155672
rect 532660 155660 532666 155712
rect 250898 155592 250904 155644
rect 250956 155632 250962 155644
rect 262677 155635 262735 155641
rect 262677 155632 262689 155635
rect 250956 155604 262689 155632
rect 250956 155592 250962 155604
rect 262677 155601 262689 155604
rect 262723 155601 262735 155635
rect 262677 155595 262735 155601
rect 262766 155592 262772 155644
rect 262824 155632 262830 155644
rect 287793 155635 287851 155641
rect 287793 155632 287805 155635
rect 262824 155604 287805 155632
rect 262824 155592 262830 155604
rect 287793 155601 287805 155604
rect 287839 155601 287851 155635
rect 287793 155595 287851 155601
rect 287885 155635 287943 155641
rect 287885 155601 287897 155635
rect 287931 155632 287943 155635
rect 295518 155632 295524 155644
rect 287931 155604 295524 155632
rect 287931 155601 287943 155604
rect 287885 155595 287943 155601
rect 295518 155592 295524 155604
rect 295576 155592 295582 155644
rect 295794 155592 295800 155644
rect 295852 155632 295858 155644
rect 317046 155632 317052 155644
rect 295852 155604 317052 155632
rect 295852 155592 295858 155604
rect 317046 155592 317052 155604
rect 317104 155592 317110 155644
rect 317230 155592 317236 155644
rect 317288 155632 317294 155644
rect 331306 155632 331312 155644
rect 317288 155604 331312 155632
rect 317288 155592 317294 155604
rect 331306 155592 331312 155604
rect 331364 155592 331370 155644
rect 333790 155592 333796 155644
rect 333848 155632 333854 155644
rect 338942 155632 338948 155644
rect 333848 155604 338948 155632
rect 333848 155592 333854 155604
rect 338942 155592 338948 155604
rect 339000 155592 339006 155644
rect 342530 155592 342536 155644
rect 342588 155632 342594 155644
rect 348234 155632 348240 155644
rect 342588 155604 348240 155632
rect 342588 155592 342594 155604
rect 348234 155592 348240 155604
rect 348292 155592 348298 155644
rect 379698 155592 379704 155644
rect 379756 155632 379762 155644
rect 382550 155632 382556 155644
rect 379756 155604 382556 155632
rect 379756 155592 379762 155604
rect 382550 155592 382556 155604
rect 382608 155592 382614 155644
rect 404078 155592 404084 155644
rect 404136 155632 404142 155644
rect 425422 155632 425428 155644
rect 404136 155604 425428 155632
rect 404136 155592 404142 155604
rect 425422 155592 425428 155604
rect 425480 155592 425486 155644
rect 425517 155635 425575 155641
rect 425517 155601 425529 155635
rect 425563 155632 425575 155635
rect 426529 155635 426587 155641
rect 426529 155632 426541 155635
rect 425563 155604 426541 155632
rect 425563 155601 425575 155604
rect 425517 155595 425575 155601
rect 426529 155601 426541 155604
rect 426575 155601 426587 155635
rect 426529 155595 426587 155601
rect 427630 155592 427636 155644
rect 427688 155632 427694 155644
rect 460474 155632 460480 155644
rect 427688 155604 429424 155632
rect 427688 155592 427694 155604
rect 242216 155536 249196 155564
rect 242216 155524 242222 155536
rect 249978 155524 249984 155576
rect 250036 155564 250042 155576
rect 280065 155567 280123 155573
rect 280065 155564 280077 155567
rect 250036 155536 280077 155564
rect 250036 155524 250042 155536
rect 280065 155533 280077 155536
rect 280111 155533 280123 155567
rect 280065 155527 280123 155533
rect 280154 155524 280160 155576
rect 280212 155564 280218 155576
rect 290826 155564 290832 155576
rect 280212 155536 290832 155564
rect 280212 155524 280218 155536
rect 290826 155524 290832 155536
rect 290884 155524 290890 155576
rect 290918 155524 290924 155576
rect 290976 155564 290982 155576
rect 296533 155567 296591 155573
rect 296533 155564 296545 155567
rect 290976 155536 296545 155564
rect 290976 155524 290982 155536
rect 296533 155533 296545 155536
rect 296579 155533 296591 155567
rect 296533 155527 296591 155533
rect 296625 155567 296683 155573
rect 296625 155533 296637 155567
rect 296671 155564 296683 155567
rect 311894 155564 311900 155576
rect 296671 155536 311900 155564
rect 296671 155533 296683 155536
rect 296625 155527 296683 155533
rect 311894 155524 311900 155536
rect 311952 155524 311958 155576
rect 313274 155524 313280 155576
rect 313332 155564 313338 155576
rect 328730 155564 328736 155576
rect 313332 155536 328736 155564
rect 313332 155524 313338 155536
rect 328730 155524 328736 155536
rect 328788 155524 328794 155576
rect 329926 155524 329932 155576
rect 329984 155564 329990 155576
rect 335630 155564 335636 155576
rect 329984 155536 335636 155564
rect 329984 155524 329990 155536
rect 335630 155524 335636 155536
rect 335688 155524 335694 155576
rect 335722 155524 335728 155576
rect 335780 155564 335786 155576
rect 340966 155564 340972 155576
rect 335780 155536 340972 155564
rect 335780 155524 335786 155536
rect 340966 155524 340972 155536
rect 341024 155524 341030 155576
rect 345474 155524 345480 155576
rect 345532 155564 345538 155576
rect 347590 155564 347596 155576
rect 345532 155536 347596 155564
rect 345532 155524 345538 155536
rect 347590 155524 347596 155536
rect 347648 155524 347654 155576
rect 356238 155524 356244 155576
rect 356296 155564 356302 155576
rect 357434 155564 357440 155576
rect 356296 155536 357440 155564
rect 356296 155524 356302 155536
rect 357434 155524 357440 155536
rect 357492 155524 357498 155576
rect 358170 155524 358176 155576
rect 358228 155564 358234 155576
rect 358814 155564 358820 155576
rect 358228 155536 358820 155564
rect 358228 155524 358234 155536
rect 358814 155524 358820 155536
rect 358872 155524 358878 155576
rect 378134 155524 378140 155576
rect 378192 155564 378198 155576
rect 380618 155564 380624 155576
rect 378192 155536 380624 155564
rect 378192 155524 378198 155536
rect 380618 155524 380624 155536
rect 380676 155524 380682 155576
rect 386322 155524 386328 155576
rect 386380 155564 386386 155576
rect 389358 155564 389364 155576
rect 386380 155536 389364 155564
rect 386380 155524 386386 155536
rect 389358 155524 389364 155536
rect 389416 155524 389422 155576
rect 406746 155524 406752 155576
rect 406804 155564 406810 155576
rect 429286 155564 429292 155576
rect 406804 155536 429292 155564
rect 406804 155524 406810 155536
rect 429286 155524 429292 155536
rect 429344 155524 429350 155576
rect 429396 155564 429424 155604
rect 430408 155604 460480 155632
rect 430408 155564 430436 155604
rect 460474 155592 460480 155604
rect 460532 155592 460538 155644
rect 478322 155592 478328 155644
rect 478380 155632 478386 155644
rect 536558 155632 536564 155644
rect 478380 155604 536564 155632
rect 478380 155592 478386 155604
rect 536558 155592 536564 155604
rect 536616 155592 536622 155644
rect 571978 155592 571984 155644
rect 572036 155632 572042 155644
rect 576486 155632 576492 155644
rect 572036 155604 576492 155632
rect 572036 155592 572042 155604
rect 576486 155592 576492 155604
rect 576544 155592 576550 155644
rect 429396 155536 430436 155564
rect 430482 155524 430488 155576
rect 430540 155564 430546 155576
rect 465350 155564 465356 155576
rect 430540 155536 465356 155564
rect 430540 155524 430546 155536
rect 465350 155524 465356 155536
rect 465408 155524 465414 155576
rect 480898 155524 480904 155576
rect 480956 155564 480962 155576
rect 540422 155564 540428 155576
rect 480956 155536 540428 155564
rect 480956 155524 480962 155536
rect 540422 155524 540428 155536
rect 540480 155524 540486 155576
rect 573358 155524 573364 155576
rect 573416 155564 573422 155576
rect 574554 155564 574560 155576
rect 573416 155536 574560 155564
rect 573416 155524 573422 155536
rect 574554 155524 574560 155536
rect 574612 155524 574618 155576
rect 27706 155456 27712 155508
rect 27764 155496 27770 155508
rect 27764 155468 127940 155496
rect 27764 155456 27770 155468
rect 23842 155388 23848 155440
rect 23900 155428 23906 155440
rect 125137 155431 125195 155437
rect 125137 155428 125149 155431
rect 23900 155400 125149 155428
rect 23900 155388 23906 155400
rect 125137 155397 125149 155400
rect 125183 155397 125195 155431
rect 125137 155391 125195 155397
rect 125226 155388 125232 155440
rect 125284 155428 125290 155440
rect 127621 155431 127679 155437
rect 127621 155428 127633 155431
rect 125284 155400 127633 155428
rect 125284 155388 125290 155400
rect 127621 155397 127633 155400
rect 127667 155397 127679 155431
rect 127621 155391 127679 155397
rect 19886 155320 19892 155372
rect 19944 155360 19950 155372
rect 126054 155360 126060 155372
rect 19944 155332 126060 155360
rect 19944 155320 19950 155332
rect 126054 155320 126060 155332
rect 126112 155320 126118 155372
rect 126146 155320 126152 155372
rect 126204 155360 126210 155372
rect 127805 155363 127863 155369
rect 127805 155360 127817 155363
rect 126204 155332 127817 155360
rect 126204 155320 126210 155332
rect 127805 155329 127817 155332
rect 127851 155329 127863 155363
rect 127912 155360 127940 155468
rect 132954 155456 132960 155508
rect 133012 155496 133018 155508
rect 137741 155499 137799 155505
rect 137741 155496 137753 155499
rect 133012 155468 137753 155496
rect 133012 155456 133018 155468
rect 137741 155465 137753 155468
rect 137787 155465 137799 155499
rect 137741 155459 137799 155465
rect 137830 155456 137836 155508
rect 137888 155496 137894 155508
rect 146849 155499 146907 155505
rect 146849 155496 146861 155499
rect 137888 155468 146861 155496
rect 137888 155456 137894 155468
rect 146849 155465 146861 155468
rect 146895 155465 146907 155499
rect 146849 155459 146907 155465
rect 147582 155456 147588 155508
rect 147640 155496 147646 155508
rect 155862 155496 155868 155508
rect 147640 155468 155868 155496
rect 147640 155456 147646 155468
rect 155862 155456 155868 155468
rect 155920 155456 155926 155508
rect 155957 155499 156015 155505
rect 155957 155465 155969 155499
rect 156003 155496 156015 155499
rect 156417 155499 156475 155505
rect 156417 155496 156429 155499
rect 156003 155468 156429 155496
rect 156003 155465 156015 155468
rect 155957 155459 156015 155465
rect 156417 155465 156429 155468
rect 156463 155465 156475 155499
rect 158714 155496 158720 155508
rect 156417 155459 156475 155465
rect 156524 155468 158720 155496
rect 127989 155431 128047 155437
rect 127989 155397 128001 155431
rect 128035 155428 128047 155431
rect 133417 155431 133475 155437
rect 133417 155428 133429 155431
rect 128035 155400 133429 155428
rect 128035 155397 128047 155400
rect 127989 155391 128047 155397
rect 133417 155397 133429 155400
rect 133463 155397 133475 155431
rect 133417 155391 133475 155397
rect 133509 155431 133567 155437
rect 133509 155397 133521 155431
rect 133555 155428 133567 155431
rect 135162 155428 135168 155440
rect 133555 155400 135168 155428
rect 133555 155397 133567 155400
rect 133509 155391 133567 155397
rect 135162 155388 135168 155400
rect 135220 155388 135226 155440
rect 137281 155431 137339 155437
rect 137281 155397 137293 155431
rect 137327 155428 137339 155431
rect 144730 155428 144736 155440
rect 137327 155400 144736 155428
rect 137327 155397 137339 155400
rect 137281 155391 137339 155397
rect 144730 155388 144736 155400
rect 144788 155388 144794 155440
rect 144822 155388 144828 155440
rect 144880 155428 144886 155440
rect 146754 155428 146760 155440
rect 144880 155400 146760 155428
rect 144880 155388 144886 155400
rect 146754 155388 146760 155400
rect 146812 155388 146818 155440
rect 146941 155431 146999 155437
rect 146941 155397 146953 155431
rect 146987 155428 146999 155431
rect 156524 155428 156552 155468
rect 158714 155456 158720 155468
rect 158772 155456 158778 155508
rect 159266 155456 159272 155508
rect 159324 155496 159330 155508
rect 163038 155496 163044 155508
rect 159324 155468 163044 155496
rect 159324 155456 159330 155468
rect 163038 155456 163044 155468
rect 163096 155456 163102 155508
rect 164142 155456 164148 155508
rect 164200 155496 164206 155508
rect 229278 155496 229284 155508
rect 164200 155468 229284 155496
rect 164200 155456 164206 155468
rect 229278 155456 229284 155468
rect 229336 155456 229342 155508
rect 230474 155456 230480 155508
rect 230532 155496 230538 155508
rect 233142 155496 233148 155508
rect 230532 155468 233148 155496
rect 230532 155456 230538 155468
rect 233142 155456 233148 155468
rect 233200 155456 233206 155508
rect 233881 155499 233939 155505
rect 233881 155465 233893 155499
rect 233927 155496 233939 155499
rect 265066 155496 265072 155508
rect 233927 155468 265072 155496
rect 233927 155465 233939 155468
rect 233881 155459 233939 155465
rect 265066 155456 265072 155468
rect 265124 155456 265130 155508
rect 265526 155456 265532 155508
rect 265584 155496 265590 155508
rect 266446 155496 266452 155508
rect 265584 155468 266452 155496
rect 265584 155456 265590 155468
rect 266446 155456 266452 155468
rect 266504 155456 266510 155508
rect 266538 155456 266544 155508
rect 266596 155496 266602 155508
rect 272521 155499 272579 155505
rect 272521 155496 272533 155499
rect 266596 155468 272533 155496
rect 266596 155456 266602 155468
rect 272521 155465 272533 155468
rect 272567 155465 272579 155499
rect 272521 155459 272579 155465
rect 274358 155456 274364 155508
rect 274416 155496 274422 155508
rect 274416 155468 296852 155496
rect 274416 155456 274422 155468
rect 146987 155400 156552 155428
rect 156601 155431 156659 155437
rect 146987 155397 146999 155400
rect 146941 155391 146999 155397
rect 156601 155397 156613 155431
rect 156647 155428 156659 155431
rect 162118 155428 162124 155440
rect 156647 155400 162124 155428
rect 156647 155397 156659 155400
rect 156601 155391 156659 155397
rect 162118 155388 162124 155400
rect 162176 155388 162182 155440
rect 163222 155388 163228 155440
rect 163280 155428 163286 155440
rect 165522 155428 165528 155440
rect 163280 155400 165528 155428
rect 163280 155388 163286 155400
rect 165522 155388 165528 155400
rect 165580 155388 165586 155440
rect 166261 155431 166319 155437
rect 166261 155397 166273 155431
rect 166307 155428 166319 155431
rect 226518 155428 226524 155440
rect 166307 155400 226524 155428
rect 166307 155397 166319 155400
rect 166261 155391 166319 155397
rect 226518 155388 226524 155400
rect 226576 155388 226582 155440
rect 226610 155388 226616 155440
rect 226668 155428 226674 155440
rect 233234 155428 233240 155440
rect 226668 155400 233240 155428
rect 226668 155388 226674 155400
rect 233234 155388 233240 155400
rect 233292 155388 233298 155440
rect 233329 155431 233387 155437
rect 233329 155397 233341 155431
rect 233375 155428 233387 155431
rect 234614 155428 234620 155440
rect 233375 155400 234620 155428
rect 233375 155397 233387 155400
rect 233329 155391 233387 155397
rect 234614 155388 234620 155400
rect 234672 155388 234678 155440
rect 238294 155388 238300 155440
rect 238352 155428 238358 155440
rect 272613 155431 272671 155437
rect 238352 155400 272564 155428
rect 238352 155388 238358 155400
rect 133782 155360 133788 155372
rect 127912 155332 133788 155360
rect 127805 155323 127863 155329
rect 133782 155320 133788 155332
rect 133840 155320 133846 155372
rect 133966 155320 133972 155372
rect 134024 155360 134030 155372
rect 209038 155360 209044 155372
rect 134024 155332 209044 155360
rect 134024 155320 134030 155332
rect 209038 155320 209044 155332
rect 209096 155320 209102 155372
rect 210970 155320 210976 155372
rect 211028 155360 211034 155372
rect 249061 155363 249119 155369
rect 249061 155360 249073 155363
rect 211028 155332 249073 155360
rect 211028 155320 211034 155332
rect 249061 155329 249073 155332
rect 249107 155329 249119 155363
rect 249061 155323 249119 155329
rect 249153 155363 249211 155369
rect 249153 155329 249165 155363
rect 249199 155360 249211 155363
rect 252649 155363 252707 155369
rect 252649 155360 252661 155363
rect 249199 155332 252661 155360
rect 249199 155329 249211 155332
rect 249153 155323 249211 155329
rect 252649 155329 252661 155332
rect 252695 155329 252707 155363
rect 252649 155323 252707 155329
rect 253198 155320 253204 155372
rect 253256 155360 253262 155372
rect 262861 155363 262919 155369
rect 262861 155360 262873 155363
rect 253256 155332 262873 155360
rect 253256 155320 253262 155332
rect 262861 155329 262873 155332
rect 262907 155329 262919 155363
rect 262861 155323 262919 155329
rect 262953 155363 263011 155369
rect 262953 155329 262965 155363
rect 262999 155360 263011 155363
rect 272429 155363 272487 155369
rect 272429 155360 272441 155363
rect 262999 155332 272441 155360
rect 262999 155329 263011 155332
rect 262953 155323 263011 155329
rect 272429 155329 272441 155332
rect 272475 155329 272487 155363
rect 272536 155360 272564 155400
rect 272613 155397 272625 155431
rect 272659 155428 272671 155431
rect 279142 155428 279148 155440
rect 272659 155400 279148 155428
rect 272659 155397 272671 155400
rect 272613 155391 272671 155397
rect 279142 155388 279148 155400
rect 279200 155388 279206 155440
rect 279234 155388 279240 155440
rect 279292 155428 279298 155440
rect 296714 155428 296720 155440
rect 279292 155400 296720 155428
rect 279292 155388 279298 155400
rect 296714 155388 296720 155400
rect 296772 155388 296778 155440
rect 296824 155428 296852 155468
rect 296898 155456 296904 155508
rect 296956 155496 296962 155508
rect 308398 155496 308404 155508
rect 296956 155468 308404 155496
rect 296956 155456 296962 155468
rect 308398 155456 308404 155468
rect 308456 155456 308462 155508
rect 308490 155456 308496 155508
rect 308548 155496 308554 155508
rect 324406 155496 324412 155508
rect 308548 155468 324412 155496
rect 308548 155456 308554 155468
rect 324406 155456 324412 155468
rect 324464 155456 324470 155508
rect 325970 155456 325976 155508
rect 326028 155496 326034 155508
rect 337194 155496 337200 155508
rect 326028 155468 337200 155496
rect 326028 155456 326034 155468
rect 337194 155456 337200 155468
rect 337252 155456 337258 155508
rect 337654 155456 337660 155508
rect 337712 155496 337718 155508
rect 342530 155496 342536 155508
rect 337712 155468 342536 155496
rect 337712 155456 337718 155468
rect 342530 155456 342536 155468
rect 342588 155456 342594 155508
rect 344554 155456 344560 155508
rect 344612 155496 344618 155508
rect 349522 155496 349528 155508
rect 344612 155468 349528 155496
rect 344612 155456 344618 155468
rect 349522 155456 349528 155468
rect 349580 155456 349586 155508
rect 380894 155456 380900 155508
rect 380952 155496 380958 155508
rect 384482 155496 384488 155508
rect 380952 155468 384488 155496
rect 380952 155456 380958 155468
rect 384482 155456 384488 155468
rect 384540 155456 384546 155508
rect 384758 155456 384764 155508
rect 384816 155496 384822 155508
rect 388346 155496 388352 155508
rect 384816 155468 388352 155496
rect 384816 155456 384822 155468
rect 388346 155456 388352 155468
rect 388404 155456 388410 155508
rect 404630 155456 404636 155508
rect 404688 155496 404694 155508
rect 407850 155496 407856 155508
rect 404688 155468 407856 155496
rect 404688 155456 404694 155468
rect 407850 155456 407856 155468
rect 407908 155456 407914 155508
rect 408310 155456 408316 155508
rect 408368 155496 408374 155508
rect 432230 155496 432236 155508
rect 408368 155468 432236 155496
rect 408368 155456 408374 155468
rect 432230 155456 432236 155468
rect 432288 155456 432294 155508
rect 433058 155456 433064 155508
rect 433116 155496 433122 155508
rect 469306 155496 469312 155508
rect 433116 155468 469312 155496
rect 433116 155456 433122 155468
rect 469306 155456 469312 155468
rect 469364 155456 469370 155508
rect 484854 155456 484860 155508
rect 484912 155496 484918 155508
rect 546310 155496 546316 155508
rect 484912 155468 546316 155496
rect 484912 155456 484918 155468
rect 546310 155456 546316 155468
rect 546368 155456 546374 155508
rect 296824 155400 301176 155428
rect 277302 155360 277308 155372
rect 272536 155332 277308 155360
rect 272429 155323 272487 155329
rect 277302 155320 277308 155332
rect 277360 155320 277366 155372
rect 277581 155363 277639 155369
rect 277581 155329 277593 155363
rect 277627 155360 277639 155363
rect 301041 155363 301099 155369
rect 301041 155360 301053 155363
rect 277627 155332 301053 155360
rect 277627 155329 277639 155332
rect 277581 155323 277639 155329
rect 301041 155329 301053 155332
rect 301087 155329 301099 155363
rect 301041 155323 301099 155329
rect 14090 155252 14096 155304
rect 14148 155292 14154 155304
rect 24854 155292 24860 155304
rect 14148 155264 24860 155292
rect 14148 155252 14154 155264
rect 24854 155252 24860 155264
rect 24912 155252 24918 155304
rect 31662 155252 31668 155304
rect 31720 155292 31726 155304
rect 133325 155295 133383 155301
rect 31720 155264 133276 155292
rect 31720 155252 31726 155264
rect 474 155184 480 155236
rect 532 155224 538 155236
rect 1302 155224 1308 155236
rect 532 155196 1308 155224
rect 532 155184 538 155196
rect 1302 155184 1308 155196
rect 1360 155184 1366 155236
rect 8202 155184 8208 155236
rect 8260 155224 8266 155236
rect 125042 155224 125048 155236
rect 8260 155196 125048 155224
rect 8260 155184 8266 155196
rect 125042 155184 125048 155196
rect 125100 155184 125106 155236
rect 125137 155227 125195 155233
rect 125137 155193 125149 155227
rect 125183 155224 125195 155227
rect 127529 155227 127587 155233
rect 127529 155224 127541 155227
rect 125183 155196 127541 155224
rect 125183 155193 125195 155196
rect 125137 155187 125195 155193
rect 127529 155193 127541 155196
rect 127575 155193 127587 155227
rect 127529 155187 127587 155193
rect 127621 155227 127679 155233
rect 127621 155193 127633 155227
rect 127667 155224 127679 155227
rect 133141 155227 133199 155233
rect 133141 155224 133153 155227
rect 127667 155196 133153 155224
rect 127667 155193 127679 155196
rect 127621 155187 127679 155193
rect 133141 155193 133153 155196
rect 133187 155193 133199 155227
rect 133248 155224 133276 155264
rect 133325 155261 133337 155295
rect 133371 155292 133383 155295
rect 138014 155292 138020 155304
rect 133371 155264 138020 155292
rect 133371 155261 133383 155264
rect 133325 155255 133383 155261
rect 138014 155252 138020 155264
rect 138072 155252 138078 155304
rect 138109 155295 138167 155301
rect 138109 155261 138121 155295
rect 138155 155292 138167 155295
rect 138155 155264 140912 155292
rect 138155 155261 138167 155264
rect 138109 155255 138167 155261
rect 136726 155224 136732 155236
rect 133248 155196 136732 155224
rect 133141 155187 133199 155193
rect 136726 155184 136732 155196
rect 136784 155184 136790 155236
rect 136821 155227 136879 155233
rect 136821 155193 136833 155227
rect 136867 155224 136879 155227
rect 140774 155224 140780 155236
rect 136867 155196 140780 155224
rect 136867 155193 136879 155196
rect 136821 155187 136879 155193
rect 140774 155184 140780 155196
rect 140832 155184 140838 155236
rect 140884 155224 140912 155264
rect 141786 155252 141792 155304
rect 141844 155292 141850 155304
rect 213825 155295 213883 155301
rect 213825 155292 213837 155295
rect 141844 155264 213837 155292
rect 141844 155252 141850 155264
rect 213825 155261 213837 155264
rect 213871 155261 213883 155295
rect 213825 155255 213883 155261
rect 213914 155252 213920 155304
rect 213972 155292 213978 155304
rect 262398 155292 262404 155304
rect 213972 155264 262404 155292
rect 213972 155252 213978 155264
rect 262398 155252 262404 155264
rect 262456 155252 262462 155304
rect 262769 155295 262827 155301
rect 262769 155261 262781 155295
rect 262815 155292 262827 155295
rect 270310 155292 270316 155304
rect 262815 155264 270316 155292
rect 262815 155261 262827 155264
rect 262769 155255 262827 155261
rect 270310 155252 270316 155264
rect 270368 155252 270374 155304
rect 270402 155252 270408 155304
rect 270460 155292 270466 155304
rect 300118 155292 300124 155304
rect 270460 155264 300124 155292
rect 270460 155252 270466 155264
rect 300118 155252 300124 155264
rect 300176 155252 300182 155304
rect 301148 155292 301176 155400
rect 306466 155388 306472 155440
rect 306524 155428 306530 155440
rect 324222 155428 324228 155440
rect 306524 155400 324228 155428
rect 306524 155388 306530 155400
rect 324222 155388 324228 155400
rect 324280 155388 324286 155440
rect 327902 155388 327908 155440
rect 327960 155428 327966 155440
rect 338482 155428 338488 155440
rect 327960 155400 338488 155428
rect 327960 155388 327966 155400
rect 338482 155388 338488 155400
rect 338540 155388 338546 155440
rect 409690 155388 409696 155440
rect 409748 155428 409754 155440
rect 434162 155428 434168 155440
rect 409748 155400 434168 155428
rect 409748 155388 409754 155400
rect 434162 155388 434168 155400
rect 434220 155388 434226 155440
rect 436002 155388 436008 155440
rect 436060 155428 436066 155440
rect 473170 155428 473176 155440
rect 436060 155400 473176 155428
rect 436060 155388 436066 155400
rect 473170 155388 473176 155400
rect 473228 155388 473234 155440
rect 483566 155388 483572 155440
rect 483624 155428 483630 155440
rect 544286 155428 544292 155440
rect 483624 155400 544292 155428
rect 483624 155388 483630 155400
rect 544286 155388 544292 155400
rect 544344 155388 544350 155440
rect 549162 155388 549168 155440
rect 549220 155428 549226 155440
rect 572622 155428 572628 155440
rect 549220 155400 572628 155428
rect 549220 155388 549226 155400
rect 572622 155388 572628 155400
rect 572680 155388 572686 155440
rect 301501 155363 301559 155369
rect 301501 155329 301513 155363
rect 301547 155360 301559 155363
rect 307389 155363 307447 155369
rect 307389 155360 307401 155363
rect 301547 155332 307401 155360
rect 301547 155329 301559 155332
rect 301501 155323 301559 155329
rect 307389 155329 307401 155332
rect 307435 155329 307447 155363
rect 307389 155323 307447 155329
rect 307478 155320 307484 155372
rect 307536 155360 307542 155372
rect 324130 155360 324136 155372
rect 307536 155332 324136 155360
rect 307536 155320 307542 155332
rect 324130 155320 324136 155332
rect 324188 155320 324194 155372
rect 325050 155320 325056 155372
rect 325108 155360 325114 155372
rect 336642 155360 336648 155372
rect 325108 155332 336648 155360
rect 325108 155320 325114 155332
rect 336642 155320 336648 155332
rect 336700 155320 336706 155372
rect 401594 155320 401600 155372
rect 401652 155360 401658 155372
rect 404906 155360 404912 155372
rect 401652 155332 404912 155360
rect 401652 155320 401658 155332
rect 404906 155320 404912 155332
rect 404964 155320 404970 155372
rect 411162 155320 411168 155372
rect 411220 155360 411226 155372
rect 436094 155360 436100 155372
rect 411220 155332 436100 155360
rect 411220 155320 411226 155332
rect 436094 155320 436100 155332
rect 436152 155320 436158 155372
rect 438670 155320 438676 155372
rect 438728 155360 438734 155372
rect 477034 155360 477040 155372
rect 438728 155332 477040 155360
rect 438728 155320 438734 155332
rect 477034 155320 477040 155332
rect 477092 155320 477098 155372
rect 491202 155320 491208 155372
rect 491260 155360 491266 155372
rect 556062 155360 556068 155372
rect 491260 155332 556068 155360
rect 491260 155320 491266 155332
rect 556062 155320 556068 155332
rect 556120 155320 556126 155372
rect 302510 155292 302516 155304
rect 301148 155264 302516 155292
rect 302510 155252 302516 155264
rect 302568 155252 302574 155304
rect 302602 155252 302608 155304
rect 302660 155292 302666 155304
rect 321646 155292 321652 155304
rect 302660 155264 321652 155292
rect 302660 155252 302666 155264
rect 321646 155252 321652 155264
rect 321704 155252 321710 155304
rect 326982 155252 326988 155304
rect 327040 155292 327046 155304
rect 338022 155292 338028 155304
rect 327040 155264 338028 155292
rect 327040 155252 327046 155264
rect 338022 155252 338028 155264
rect 338080 155252 338086 155304
rect 414566 155252 414572 155304
rect 414624 155292 414630 155304
rect 440970 155292 440976 155304
rect 414624 155264 440976 155292
rect 414624 155252 414630 155264
rect 440970 155252 440976 155264
rect 441028 155252 441034 155304
rect 441246 155252 441252 155304
rect 441304 155292 441310 155304
rect 480990 155292 480996 155304
rect 441304 155264 480996 155292
rect 441304 155252 441310 155264
rect 480990 155252 480996 155264
rect 481048 155252 481054 155304
rect 488350 155252 488356 155304
rect 488408 155292 488414 155304
rect 552106 155292 552112 155304
rect 488408 155264 552112 155292
rect 488408 155252 488414 155264
rect 552106 155252 552112 155264
rect 552164 155252 552170 155304
rect 554774 155252 554780 155304
rect 554832 155292 554838 155304
rect 569678 155292 569684 155304
rect 554832 155264 569684 155292
rect 554832 155252 554838 155264
rect 569678 155252 569684 155264
rect 569736 155252 569742 155304
rect 208394 155224 208400 155236
rect 140884 155196 208400 155224
rect 208394 155184 208400 155196
rect 208452 155184 208458 155236
rect 209958 155184 209964 155236
rect 210016 155224 210022 155236
rect 259822 155224 259828 155236
rect 210016 155196 259828 155224
rect 210016 155184 210022 155196
rect 259822 155184 259828 155196
rect 259880 155184 259886 155236
rect 260650 155184 260656 155236
rect 260708 155224 260714 155236
rect 263505 155227 263563 155233
rect 263505 155224 263517 155227
rect 260708 155196 263517 155224
rect 260708 155184 260714 155196
rect 263505 155193 263517 155196
rect 263551 155193 263563 155227
rect 263505 155187 263563 155193
rect 263594 155184 263600 155236
rect 263652 155224 263658 155236
rect 287885 155227 287943 155233
rect 287885 155224 287897 155227
rect 263652 155196 287897 155224
rect 263652 155184 263658 155196
rect 287885 155193 287897 155196
rect 287931 155193 287943 155227
rect 287885 155187 287943 155193
rect 287974 155184 287980 155236
rect 288032 155224 288038 155236
rect 296625 155227 296683 155233
rect 296625 155224 296637 155227
rect 288032 155196 296637 155224
rect 288032 155184 288038 155196
rect 296625 155193 296637 155196
rect 296671 155193 296683 155227
rect 296625 155187 296683 155193
rect 296714 155184 296720 155236
rect 296772 155224 296778 155236
rect 296772 155196 298692 155224
rect 296772 155184 296778 155196
rect 29638 155116 29644 155168
rect 29696 155156 29702 155168
rect 31662 155156 31668 155168
rect 29696 155128 31668 155156
rect 29696 155116 29702 155128
rect 31662 155116 31668 155128
rect 31720 155116 31726 155168
rect 55030 155116 55036 155168
rect 55088 155156 55094 155168
rect 70394 155156 70400 155168
rect 55088 155128 70400 155156
rect 55088 155116 55094 155128
rect 70394 155116 70400 155128
rect 70452 155116 70458 155168
rect 90082 155116 90088 155168
rect 90140 155156 90146 155168
rect 168374 155156 168380 155168
rect 90140 155128 168380 155156
rect 90140 155116 90146 155128
rect 168374 155116 168380 155128
rect 168432 155116 168438 155168
rect 169018 155116 169024 155168
rect 169076 155156 169082 155168
rect 172422 155156 172428 155168
rect 169076 155128 172428 155156
rect 169076 155116 169082 155128
rect 172422 155116 172428 155128
rect 172480 155116 172486 155168
rect 172974 155116 172980 155168
rect 173032 155156 173038 155168
rect 229186 155156 229192 155168
rect 173032 155128 229192 155156
rect 173032 155116 173038 155128
rect 229186 155116 229192 155128
rect 229244 155116 229250 155168
rect 229373 155159 229431 155165
rect 229373 155125 229385 155159
rect 229419 155156 229431 155159
rect 239582 155156 239588 155168
rect 229419 155128 239588 155156
rect 229419 155125 229431 155128
rect 229373 155119 229431 155125
rect 239582 155116 239588 155128
rect 239640 155116 239646 155168
rect 241057 155159 241115 155165
rect 241057 155125 241069 155159
rect 241103 155156 241115 155159
rect 243449 155159 243507 155165
rect 243449 155156 243461 155159
rect 241103 155128 243461 155156
rect 241103 155125 241115 155128
rect 241057 155119 241115 155125
rect 243449 155125 243461 155128
rect 243495 155125 243507 155159
rect 243449 155119 243507 155125
rect 243541 155159 243599 155165
rect 243541 155125 243553 155159
rect 243587 155156 243599 155159
rect 269301 155159 269359 155165
rect 269301 155156 269313 155159
rect 243587 155128 269313 155156
rect 243587 155125 243599 155128
rect 243541 155119 243599 155125
rect 269301 155125 269313 155128
rect 269347 155125 269359 155159
rect 269301 155119 269359 155125
rect 269390 155116 269396 155168
rect 269448 155156 269454 155168
rect 274634 155156 274640 155168
rect 269448 155128 274640 155156
rect 269448 155116 269454 155128
rect 274634 155116 274640 155128
rect 274692 155116 274698 155168
rect 275278 155116 275284 155168
rect 275336 155156 275342 155168
rect 277581 155159 277639 155165
rect 277581 155156 277593 155159
rect 275336 155128 277593 155156
rect 275336 155116 275342 155128
rect 277581 155125 277593 155128
rect 277627 155125 277639 155159
rect 298002 155156 298008 155168
rect 277581 155119 277639 155125
rect 277688 155128 298008 155156
rect 51166 155048 51172 155100
rect 51224 155088 51230 155100
rect 67358 155088 67364 155100
rect 51224 155060 67364 155088
rect 51224 155048 51230 155060
rect 67358 155048 67364 155060
rect 67416 155048 67422 155100
rect 83274 155048 83280 155100
rect 83332 155088 83338 155100
rect 146941 155091 146999 155097
rect 146941 155088 146953 155091
rect 83332 155060 146953 155088
rect 83332 155048 83338 155060
rect 146941 155057 146953 155060
rect 146987 155057 146999 155091
rect 146941 155051 146999 155057
rect 148229 155091 148287 155097
rect 148229 155057 148241 155091
rect 148275 155088 148287 155091
rect 187694 155088 187700 155100
rect 148275 155060 187700 155088
rect 148275 155057 148287 155060
rect 148229 155051 148287 155057
rect 187694 155048 187700 155060
rect 187752 155048 187758 155100
rect 188522 155048 188528 155100
rect 188580 155088 188586 155100
rect 242986 155088 242992 155100
rect 188580 155060 242992 155088
rect 188580 155048 188586 155060
rect 242986 155048 242992 155060
rect 243044 155048 243050 155100
rect 243081 155091 243139 155097
rect 243081 155057 243093 155091
rect 243127 155088 243139 155091
rect 248969 155091 249027 155097
rect 243127 155060 243676 155088
rect 243127 155057 243139 155060
rect 243081 155051 243139 155057
rect 62850 154980 62856 155032
rect 62908 155020 62914 155032
rect 74994 155020 75000 155032
rect 62908 154992 75000 155020
rect 62908 154980 62914 154992
rect 74994 154980 75000 154992
rect 75052 154980 75058 155032
rect 101766 154980 101772 155032
rect 101824 155020 101830 155032
rect 108301 155023 108359 155029
rect 108301 155020 108313 155023
rect 101824 154992 108313 155020
rect 101824 154980 101830 154992
rect 108301 154989 108313 154992
rect 108347 154989 108359 155023
rect 108301 154983 108359 154989
rect 109865 155023 109923 155029
rect 109865 154989 109877 155023
rect 109911 155020 109923 155023
rect 182082 155020 182088 155032
rect 109911 154992 182088 155020
rect 109911 154989 109923 154992
rect 109865 154983 109923 154989
rect 182082 154980 182088 154992
rect 182140 154980 182146 155032
rect 182637 155023 182695 155029
rect 182637 154989 182649 155023
rect 182683 155020 182695 155023
rect 185486 155020 185492 155032
rect 182683 154992 185492 155020
rect 182683 154989 182695 154992
rect 182637 154983 182695 154989
rect 185486 154980 185492 154992
rect 185544 154980 185550 155032
rect 185581 155023 185639 155029
rect 185581 154989 185593 155023
rect 185627 155020 185639 155023
rect 193122 155020 193128 155032
rect 185627 154992 193128 155020
rect 185627 154989 185639 154992
rect 185581 154983 185639 154989
rect 193122 154980 193128 154992
rect 193180 154980 193186 155032
rect 195149 155023 195207 155029
rect 195149 154989 195161 155023
rect 195195 155020 195207 155023
rect 237190 155020 237196 155032
rect 195195 154992 237196 155020
rect 195195 154989 195207 154992
rect 195149 154983 195207 154989
rect 237190 154980 237196 154992
rect 237248 154980 237254 155032
rect 237282 154980 237288 155032
rect 237340 155020 237346 155032
rect 243541 155023 243599 155029
rect 243541 155020 243553 155023
rect 237340 154992 243553 155020
rect 237340 154980 237346 154992
rect 243541 154989 243553 154992
rect 243587 154989 243599 155023
rect 243648 155020 243676 155060
rect 248969 155057 248981 155091
rect 249015 155088 249027 155091
rect 272337 155091 272395 155097
rect 272337 155088 272349 155091
rect 249015 155060 272349 155088
rect 249015 155057 249027 155060
rect 248969 155051 249027 155057
rect 272337 155057 272349 155060
rect 272383 155057 272395 155091
rect 272337 155051 272395 155057
rect 272429 155091 272487 155097
rect 272429 155057 272441 155091
rect 272475 155088 272487 155091
rect 272705 155091 272763 155097
rect 272705 155088 272717 155091
rect 272475 155060 272717 155088
rect 272475 155057 272487 155060
rect 272429 155051 272487 155057
rect 272705 155057 272717 155060
rect 272751 155057 272763 155091
rect 272705 155051 272763 155057
rect 273346 155048 273352 155100
rect 273404 155088 273410 155100
rect 277688 155088 277716 155128
rect 298002 155116 298008 155128
rect 298060 155116 298066 155168
rect 298664 155156 298692 155196
rect 298738 155184 298744 155236
rect 298796 155224 298802 155236
rect 318978 155224 318984 155236
rect 298796 155196 318984 155224
rect 298796 155184 298802 155196
rect 318978 155184 318984 155196
rect 319036 155184 319042 155236
rect 323026 155184 323032 155236
rect 323084 155224 323090 155236
rect 334066 155224 334072 155236
rect 323084 155196 334072 155224
rect 323084 155184 323090 155196
rect 334066 155184 334072 155196
rect 334124 155184 334130 155236
rect 338666 155184 338672 155236
rect 338724 155224 338730 155236
rect 343634 155224 343640 155236
rect 338724 155196 343640 155224
rect 338724 155184 338730 155196
rect 343634 155184 343640 155196
rect 343692 155184 343698 155236
rect 382274 155184 382280 155236
rect 382332 155224 382338 155236
rect 386414 155224 386420 155236
rect 382332 155196 386420 155224
rect 382332 155184 382338 155196
rect 386414 155184 386420 155196
rect 386472 155184 386478 155236
rect 401502 155184 401508 155236
rect 401560 155224 401566 155236
rect 421558 155224 421564 155236
rect 401560 155196 421564 155224
rect 401560 155184 401566 155196
rect 421558 155184 421564 155196
rect 421616 155184 421622 155236
rect 422202 155184 422208 155236
rect 422260 155224 422266 155236
rect 452746 155224 452752 155236
rect 422260 155196 452752 155224
rect 422260 155184 422266 155196
rect 452746 155184 452752 155196
rect 452804 155184 452810 155236
rect 454862 155184 454868 155236
rect 454920 155224 454926 155236
rect 501414 155224 501420 155236
rect 454920 155196 501420 155224
rect 454920 155184 454926 155196
rect 501414 155184 501420 155196
rect 501472 155184 501478 155236
rect 503070 155184 503076 155236
rect 503128 155224 503134 155236
rect 573542 155224 573548 155236
rect 503128 155196 573548 155224
rect 503128 155184 503134 155196
rect 573542 155184 573548 155196
rect 573600 155184 573606 155236
rect 301501 155159 301559 155165
rect 301501 155156 301513 155159
rect 298664 155128 301513 155156
rect 301501 155125 301513 155128
rect 301547 155125 301559 155159
rect 301501 155119 301559 155125
rect 301590 155116 301596 155168
rect 301648 155156 301654 155168
rect 317322 155156 317328 155168
rect 301648 155128 317328 155156
rect 301648 155116 301654 155128
rect 317322 155116 317328 155128
rect 317380 155116 317386 155168
rect 318150 155116 318156 155168
rect 318208 155156 318214 155168
rect 329742 155156 329748 155168
rect 318208 155128 329748 155156
rect 318208 155116 318214 155128
rect 329742 155116 329748 155128
rect 329800 155116 329806 155168
rect 332778 155116 332784 155168
rect 332836 155156 332842 155168
rect 338574 155156 338580 155168
rect 332836 155128 338580 155156
rect 332836 155116 332842 155128
rect 338574 155116 338580 155128
rect 338632 155116 338638 155168
rect 343542 155116 343548 155168
rect 343600 155156 343606 155168
rect 349062 155156 349068 155168
rect 343600 155128 349068 155156
rect 343600 155116 343606 155128
rect 349062 155116 349068 155128
rect 349120 155116 349126 155168
rect 398558 155116 398564 155168
rect 398616 155156 398622 155168
rect 417602 155156 417608 155168
rect 398616 155128 417608 155156
rect 398616 155116 398622 155128
rect 417602 155116 417608 155128
rect 417660 155116 417666 155168
rect 419442 155116 419448 155168
rect 419500 155156 419506 155168
rect 448790 155156 448796 155168
rect 419500 155128 448796 155156
rect 419500 155116 419506 155128
rect 448790 155116 448796 155128
rect 448848 155116 448854 155168
rect 467190 155116 467196 155168
rect 467248 155156 467254 155168
rect 519998 155156 520004 155168
rect 467248 155128 520004 155156
rect 467248 155116 467254 155128
rect 519998 155116 520004 155128
rect 520056 155116 520062 155168
rect 273404 155060 277716 155088
rect 277857 155091 277915 155097
rect 273404 155048 273410 155060
rect 277857 155057 277869 155091
rect 277903 155088 277915 155091
rect 281997 155091 282055 155097
rect 281997 155088 282009 155091
rect 277903 155060 282009 155088
rect 277903 155057 277915 155060
rect 277857 155051 277915 155057
rect 281997 155057 282009 155060
rect 282043 155057 282055 155091
rect 281997 155051 282055 155057
rect 282086 155048 282092 155100
rect 282144 155088 282150 155100
rect 300581 155091 300639 155097
rect 300581 155088 300593 155091
rect 282144 155060 300593 155088
rect 282144 155048 282150 155060
rect 300581 155057 300593 155060
rect 300627 155057 300639 155091
rect 300581 155051 300639 155057
rect 300670 155048 300676 155100
rect 300728 155088 300734 155100
rect 309318 155088 309324 155100
rect 300728 155060 309324 155088
rect 300728 155048 300734 155060
rect 309318 155048 309324 155060
rect 309376 155048 309382 155100
rect 309410 155048 309416 155100
rect 309468 155088 309474 155100
rect 323210 155088 323216 155100
rect 309468 155060 323216 155088
rect 309468 155048 309474 155060
rect 323210 155048 323216 155060
rect 323268 155048 323274 155100
rect 398926 155048 398932 155100
rect 398984 155088 398990 155100
rect 401042 155088 401048 155100
rect 398984 155060 401048 155088
rect 398984 155048 398990 155060
rect 401042 155048 401048 155060
rect 401100 155048 401106 155100
rect 420546 155088 420552 155100
rect 401336 155060 420552 155088
rect 266354 155020 266360 155032
rect 243648 154992 266360 155020
rect 243541 154983 243599 154989
rect 266354 154980 266360 154992
rect 266412 154980 266418 155032
rect 268381 155023 268439 155029
rect 268381 154989 268393 155023
rect 268427 155020 268439 155023
rect 269301 155023 269359 155029
rect 269301 155020 269313 155023
rect 268427 154992 269313 155020
rect 268427 154989 268439 154992
rect 268381 154983 268439 154989
rect 269301 154989 269313 154992
rect 269347 154989 269359 155023
rect 269301 154983 269359 154989
rect 269482 154980 269488 155032
rect 269540 155020 269546 155032
rect 292574 155020 292580 155032
rect 269540 154992 292580 155020
rect 269540 154980 269546 154992
rect 292574 154980 292580 154992
rect 292632 154980 292638 155032
rect 293773 155023 293831 155029
rect 293773 154989 293785 155023
rect 293819 155020 293831 155023
rect 294690 155020 294696 155032
rect 293819 154992 294696 155020
rect 293819 154989 293831 154992
rect 293773 154983 293831 154989
rect 294690 154980 294696 154992
rect 294748 154980 294754 155032
rect 294782 154980 294788 155032
rect 294840 155020 294846 155032
rect 316402 155020 316408 155032
rect 294840 154992 316408 155020
rect 294840 154980 294846 154992
rect 316402 154980 316408 154992
rect 316460 154980 316466 155032
rect 321094 154980 321100 155032
rect 321152 155020 321158 155032
rect 332318 155020 332324 155032
rect 321152 154992 332324 155020
rect 321152 154980 321158 154992
rect 332318 154980 332324 154992
rect 332376 154980 332382 155032
rect 355226 154980 355232 155032
rect 355284 155020 355290 155032
rect 356698 155020 356704 155032
rect 355284 154992 356704 155020
rect 355284 154980 355290 154992
rect 356698 154980 356704 154992
rect 356756 154980 356762 155032
rect 400950 154980 400956 155032
rect 401008 155020 401014 155032
rect 401336 155020 401364 155060
rect 420546 155048 420552 155060
rect 420604 155048 420610 155100
rect 423030 155048 423036 155100
rect 423088 155088 423094 155100
rect 453666 155088 453672 155100
rect 423088 155060 453672 155088
rect 423088 155048 423094 155060
rect 453666 155048 453672 155060
rect 453724 155048 453730 155100
rect 463602 155048 463608 155100
rect 463660 155088 463666 155100
rect 515122 155088 515128 155100
rect 463660 155060 515128 155088
rect 463660 155048 463666 155060
rect 515122 155048 515128 155060
rect 515180 155048 515186 155100
rect 401008 154992 401364 155020
rect 401008 154980 401014 154992
rect 401686 154980 401692 155032
rect 401744 155020 401750 155032
rect 403986 155020 403992 155032
rect 401744 154992 403992 155020
rect 401744 154980 401750 154992
rect 403986 154980 403992 154992
rect 404044 154980 404050 155032
rect 418614 155020 418620 155032
rect 407776 154992 418620 155020
rect 87138 154912 87144 154964
rect 87196 154952 87202 154964
rect 156601 154955 156659 154961
rect 156601 154952 156613 154955
rect 87196 154924 156613 154952
rect 87196 154912 87202 154924
rect 156601 154921 156613 154924
rect 156647 154921 156659 154955
rect 156601 154915 156659 154921
rect 156693 154955 156751 154961
rect 156693 154921 156705 154955
rect 156739 154952 156751 154955
rect 197354 154952 197360 154964
rect 156739 154924 197360 154952
rect 156739 154921 156751 154924
rect 156693 154915 156751 154921
rect 197354 154912 197360 154924
rect 197412 154912 197418 154964
rect 207106 154912 207112 154964
rect 207164 154952 207170 154964
rect 256694 154952 256700 154964
rect 207164 154924 256700 154952
rect 207164 154912 207170 154924
rect 256694 154912 256700 154924
rect 256752 154912 256758 154964
rect 257798 154912 257804 154964
rect 257856 154952 257862 154964
rect 261389 154955 261447 154961
rect 261389 154952 261401 154955
rect 257856 154924 261401 154952
rect 257856 154912 257862 154924
rect 261389 154921 261401 154924
rect 261435 154921 261447 154955
rect 261389 154915 261447 154921
rect 262861 154955 262919 154961
rect 262861 154921 262873 154955
rect 262907 154952 262919 154955
rect 269390 154952 269396 154964
rect 262907 154924 269396 154952
rect 262907 154921 262919 154924
rect 262861 154915 262919 154921
rect 269390 154912 269396 154924
rect 269448 154912 269454 154964
rect 269577 154955 269635 154961
rect 269577 154921 269589 154955
rect 269623 154952 269635 154955
rect 271690 154952 271696 154964
rect 269623 154924 271696 154952
rect 269623 154921 269635 154924
rect 269577 154915 269635 154921
rect 271690 154912 271696 154924
rect 271748 154912 271754 154964
rect 272334 154912 272340 154964
rect 272392 154952 272398 154964
rect 275281 154955 275339 154961
rect 272392 154924 275232 154952
rect 272392 154912 272398 154924
rect 71590 154844 71596 154896
rect 71648 154884 71654 154896
rect 144822 154884 144828 154896
rect 71648 154856 144828 154884
rect 71648 154844 71654 154856
rect 144822 154844 144828 154856
rect 144880 154844 144886 154896
rect 146849 154887 146907 154893
rect 146849 154853 146861 154887
rect 146895 154884 146907 154887
rect 195974 154884 195980 154896
rect 146895 154856 195980 154884
rect 146895 154853 146907 154856
rect 146849 154847 146907 154853
rect 195974 154844 195980 154856
rect 196032 154844 196038 154896
rect 202230 154844 202236 154896
rect 202288 154884 202294 154896
rect 243541 154887 243599 154893
rect 243541 154884 243553 154887
rect 202288 154856 243553 154884
rect 202288 154844 202294 154856
rect 243541 154853 243553 154856
rect 243587 154853 243599 154887
rect 243541 154847 243599 154853
rect 243633 154887 243691 154893
rect 243633 154853 243645 154887
rect 243679 154884 243691 154887
rect 248785 154887 248843 154893
rect 248785 154884 248797 154887
rect 243679 154856 248797 154884
rect 243679 154853 243691 154856
rect 243633 154847 243691 154853
rect 248785 154853 248797 154856
rect 248831 154853 248843 154887
rect 248785 154847 248843 154853
rect 249061 154887 249119 154893
rect 249061 154853 249073 154887
rect 249107 154884 249119 154887
rect 259362 154884 259368 154896
rect 249107 154856 259368 154884
rect 249107 154853 249119 154856
rect 249061 154847 249119 154853
rect 259362 154844 259368 154856
rect 259420 154844 259426 154896
rect 262953 154887 263011 154893
rect 262953 154884 262965 154887
rect 261220 154856 262965 154884
rect 106642 154776 106648 154828
rect 106700 154816 106706 154828
rect 109865 154819 109923 154825
rect 109865 154816 109877 154819
rect 106700 154788 109877 154816
rect 106700 154776 106706 154788
rect 109865 154785 109877 154788
rect 109911 154785 109923 154819
rect 109865 154779 109923 154785
rect 117406 154776 117412 154828
rect 117464 154816 117470 154828
rect 185578 154816 185584 154828
rect 117464 154788 185584 154816
rect 117464 154776 117470 154788
rect 185578 154776 185584 154788
rect 185636 154776 185642 154828
rect 187053 154819 187111 154825
rect 187053 154785 187065 154819
rect 187099 154816 187111 154819
rect 195241 154819 195299 154825
rect 195241 154816 195253 154819
rect 187099 154788 195253 154816
rect 187099 154785 187111 154788
rect 187053 154779 187111 154785
rect 195241 154785 195253 154788
rect 195287 154785 195299 154819
rect 195241 154779 195299 154785
rect 196342 154776 196348 154828
rect 196400 154816 196406 154828
rect 245562 154816 245568 154828
rect 196400 154788 245568 154816
rect 196400 154776 196406 154788
rect 245562 154776 245568 154788
rect 245620 154776 245626 154828
rect 245933 154819 245991 154825
rect 245933 154785 245945 154819
rect 245979 154816 245991 154819
rect 248877 154819 248935 154825
rect 248877 154816 248889 154819
rect 245979 154788 248889 154816
rect 245979 154785 245991 154788
rect 245933 154779 245991 154785
rect 248877 154785 248889 154788
rect 248923 154785 248935 154819
rect 248877 154779 248935 154785
rect 248966 154776 248972 154828
rect 249024 154816 249030 154828
rect 261113 154819 261171 154825
rect 261113 154816 261125 154819
rect 249024 154788 261125 154816
rect 249024 154776 249030 154788
rect 261113 154785 261125 154788
rect 261159 154785 261171 154819
rect 261113 154779 261171 154785
rect 98914 154708 98920 154760
rect 98972 154748 98978 154760
rect 164878 154748 164884 154760
rect 98972 154720 164884 154748
rect 98972 154708 98978 154720
rect 164878 154708 164884 154720
rect 164936 154708 164942 154760
rect 165154 154708 165160 154760
rect 165212 154748 165218 154760
rect 172241 154751 172299 154757
rect 172241 154748 172253 154751
rect 165212 154720 172253 154748
rect 165212 154708 165218 154720
rect 172241 154717 172253 154720
rect 172287 154717 172299 154751
rect 172241 154711 172299 154717
rect 175921 154751 175979 154757
rect 175921 154717 175933 154751
rect 175967 154748 175979 154751
rect 179506 154748 179512 154760
rect 175967 154720 179512 154748
rect 175967 154717 175979 154720
rect 175921 154711 175979 154717
rect 179506 154708 179512 154720
rect 179564 154708 179570 154760
rect 179782 154708 179788 154760
rect 179840 154748 179846 154760
rect 185489 154751 185547 154757
rect 185489 154748 185501 154751
rect 179840 154720 185501 154748
rect 179840 154708 179846 154720
rect 185489 154717 185501 154720
rect 185535 154717 185547 154751
rect 185489 154711 185547 154717
rect 185670 154708 185676 154760
rect 185728 154748 185734 154760
rect 189074 154748 189080 154760
rect 185728 154720 189080 154748
rect 185728 154708 185734 154720
rect 189074 154708 189080 154720
rect 189132 154708 189138 154760
rect 194410 154708 194416 154760
rect 194468 154748 194474 154760
rect 194468 154720 197308 154748
rect 194468 154708 194474 154720
rect 86218 154640 86224 154692
rect 86276 154680 86282 154692
rect 91002 154680 91008 154692
rect 86276 154652 91008 154680
rect 86276 154640 86282 154652
rect 91002 154640 91008 154652
rect 91060 154640 91066 154692
rect 96890 154640 96896 154692
rect 96948 154680 96954 154692
rect 127621 154683 127679 154689
rect 127621 154680 127633 154683
rect 96948 154652 127633 154680
rect 96948 154640 96954 154652
rect 127621 154649 127633 154652
rect 127667 154649 127679 154683
rect 127621 154643 127679 154649
rect 127713 154683 127771 154689
rect 127713 154649 127725 154683
rect 127759 154680 127771 154683
rect 184290 154680 184296 154692
rect 127759 154652 184296 154680
rect 127759 154649 127771 154652
rect 127713 154643 127771 154649
rect 184290 154640 184296 154652
rect 184348 154640 184354 154692
rect 184658 154640 184664 154692
rect 184716 154680 184722 154692
rect 195149 154683 195207 154689
rect 195149 154680 195161 154683
rect 184716 154652 195161 154680
rect 184716 154640 184722 154652
rect 195149 154649 195161 154652
rect 195195 154649 195207 154683
rect 195149 154643 195207 154649
rect 195333 154683 195391 154689
rect 195333 154649 195345 154683
rect 195379 154680 195391 154683
rect 196526 154680 196532 154692
rect 195379 154652 196532 154680
rect 195379 154649 195391 154652
rect 195333 154643 195391 154649
rect 196526 154640 196532 154652
rect 196584 154640 196590 154692
rect 197280 154680 197308 154720
rect 198274 154708 198280 154760
rect 198332 154748 198338 154760
rect 211062 154748 211068 154760
rect 198332 154720 211068 154748
rect 198332 154708 198338 154720
rect 211062 154708 211068 154720
rect 211120 154708 211126 154760
rect 211982 154708 211988 154760
rect 212040 154748 212046 154760
rect 255314 154748 255320 154760
rect 212040 154720 255320 154748
rect 212040 154708 212046 154720
rect 255314 154708 255320 154720
rect 255372 154708 255378 154760
rect 256786 154708 256792 154760
rect 256844 154748 256850 154760
rect 261220 154748 261248 154856
rect 262953 154853 262965 154856
rect 262999 154853 263011 154887
rect 262953 154847 263011 154853
rect 263505 154887 263563 154893
rect 263505 154853 263517 154887
rect 263551 154884 263563 154887
rect 272613 154887 272671 154893
rect 272613 154884 272625 154887
rect 263551 154856 272625 154884
rect 263551 154853 263563 154856
rect 263505 154847 263563 154853
rect 272613 154853 272625 154856
rect 272659 154853 272671 154887
rect 272613 154847 272671 154853
rect 272705 154887 272763 154893
rect 272705 154853 272717 154887
rect 272751 154884 272763 154887
rect 275097 154887 275155 154893
rect 275097 154884 275109 154887
rect 272751 154856 275109 154884
rect 272751 154853 272763 154856
rect 272705 154847 272763 154853
rect 275097 154853 275109 154856
rect 275143 154853 275155 154887
rect 275204 154884 275232 154924
rect 275281 154921 275293 154955
rect 275327 154952 275339 154955
rect 276750 154952 276756 154964
rect 275327 154924 276756 154952
rect 275327 154921 275339 154924
rect 275281 154915 275339 154921
rect 276750 154912 276756 154924
rect 276808 154912 276814 154964
rect 277210 154912 277216 154964
rect 277268 154952 277274 154964
rect 297910 154952 297916 154964
rect 277268 154924 297916 154952
rect 277268 154912 277274 154924
rect 297910 154912 297916 154924
rect 297968 154912 297974 154964
rect 299658 154912 299664 154964
rect 299716 154952 299722 154964
rect 319622 154952 319628 154964
rect 299716 154924 319628 154952
rect 299716 154912 299722 154924
rect 319622 154912 319628 154924
rect 319680 154912 319686 154964
rect 322106 154912 322112 154964
rect 322164 154952 322170 154964
rect 333882 154952 333888 154964
rect 322164 154924 333888 154952
rect 322164 154912 322170 154924
rect 333882 154912 333888 154924
rect 333940 154912 333946 154964
rect 357158 154912 357164 154964
rect 357216 154952 357222 154964
rect 357986 154952 357992 154964
rect 357216 154924 357992 154952
rect 357216 154912 357222 154924
rect 357986 154912 357992 154924
rect 358044 154912 358050 154964
rect 365254 154912 365260 154964
rect 365312 154952 365318 154964
rect 365990 154952 365996 154964
rect 365312 154924 365996 154952
rect 365312 154912 365318 154924
rect 365990 154912 365996 154924
rect 366048 154912 366054 154964
rect 400306 154912 400312 154964
rect 400364 154952 400370 154964
rect 402974 154952 402980 154964
rect 400364 154924 402980 154952
rect 400364 154912 400370 154924
rect 402974 154912 402980 154924
rect 403032 154912 403038 154964
rect 285674 154884 285680 154896
rect 275204 154856 285680 154884
rect 275097 154847 275155 154853
rect 285674 154844 285680 154856
rect 285732 154844 285738 154896
rect 286042 154844 286048 154896
rect 286100 154884 286106 154896
rect 307662 154884 307668 154896
rect 286100 154856 307668 154884
rect 286100 154844 286106 154856
rect 307662 154844 307668 154856
rect 307720 154844 307726 154896
rect 311342 154844 311348 154896
rect 311400 154884 311406 154896
rect 321554 154884 321560 154896
rect 311400 154856 321560 154884
rect 311400 154844 311406 154856
rect 321554 154844 321560 154856
rect 321612 154844 321618 154896
rect 261297 154819 261355 154825
rect 261297 154785 261309 154819
rect 261343 154816 261355 154819
rect 276014 154816 276020 154828
rect 261343 154788 276020 154816
rect 261343 154785 261355 154788
rect 261297 154779 261355 154785
rect 276014 154776 276020 154788
rect 276072 154776 276078 154828
rect 276290 154776 276296 154828
rect 276348 154816 276354 154828
rect 289262 154816 289268 154828
rect 276348 154788 289268 154816
rect 276348 154776 276354 154788
rect 289262 154776 289268 154788
rect 289320 154776 289326 154828
rect 289357 154819 289415 154825
rect 289357 154785 289369 154819
rect 289403 154816 289415 154819
rect 293773 154819 293831 154825
rect 293773 154816 293785 154819
rect 289403 154788 293785 154816
rect 289403 154785 289415 154788
rect 289357 154779 289415 154785
rect 293773 154785 293785 154788
rect 293819 154785 293831 154819
rect 293773 154779 293831 154785
rect 293862 154776 293868 154828
rect 293920 154816 293926 154828
rect 307297 154819 307355 154825
rect 307297 154816 307309 154819
rect 293920 154788 307309 154816
rect 293920 154776 293926 154788
rect 307297 154785 307309 154788
rect 307343 154785 307355 154819
rect 307297 154779 307355 154785
rect 307389 154819 307447 154825
rect 307389 154785 307401 154819
rect 307435 154816 307447 154819
rect 308582 154816 308588 154828
rect 307435 154788 308588 154816
rect 307435 154785 307447 154788
rect 307389 154779 307447 154785
rect 308582 154776 308588 154788
rect 308640 154776 308646 154828
rect 310422 154776 310428 154828
rect 310480 154816 310486 154828
rect 323026 154816 323032 154828
rect 310480 154788 323032 154816
rect 310480 154776 310486 154788
rect 323026 154776 323032 154788
rect 323084 154776 323090 154828
rect 324038 154776 324044 154828
rect 324096 154816 324102 154828
rect 333974 154816 333980 154828
rect 324096 154788 333980 154816
rect 324096 154776 324102 154788
rect 333974 154776 333980 154788
rect 334032 154776 334038 154828
rect 341610 154776 341616 154828
rect 341668 154816 341674 154828
rect 347498 154816 347504 154828
rect 341668 154788 347504 154816
rect 341668 154776 341674 154788
rect 347498 154776 347504 154788
rect 347556 154776 347562 154828
rect 384574 154776 384580 154828
rect 384632 154816 384638 154828
rect 387426 154816 387432 154828
rect 384632 154788 387432 154816
rect 384632 154776 384638 154788
rect 387426 154776 387432 154788
rect 387484 154776 387490 154828
rect 400214 154776 400220 154828
rect 400272 154816 400278 154828
rect 402054 154816 402060 154828
rect 400272 154788 402060 154816
rect 400272 154776 400278 154788
rect 402054 154776 402060 154788
rect 402112 154776 402118 154828
rect 407776 154816 407804 154992
rect 418614 154980 418620 154992
rect 418672 154980 418678 155032
rect 420454 154980 420460 155032
rect 420512 155020 420518 155032
rect 449802 155020 449808 155032
rect 420512 154992 449808 155020
rect 420512 154980 420518 154992
rect 449802 154980 449808 154992
rect 449860 154980 449866 155032
rect 462038 154980 462044 155032
rect 462096 155020 462102 155032
rect 512178 155020 512184 155032
rect 462096 154992 512184 155020
rect 462096 154980 462102 154992
rect 512178 154980 512184 154992
rect 512236 154980 512242 155032
rect 417421 154955 417479 154961
rect 417421 154952 417433 154955
rect 402946 154788 407804 154816
rect 407868 154924 417433 154952
rect 256844 154720 261248 154748
rect 261389 154751 261447 154757
rect 256844 154708 256850 154720
rect 261389 154717 261401 154751
rect 261435 154748 261447 154751
rect 281077 154751 281135 154757
rect 281077 154748 281089 154751
rect 261435 154720 281089 154748
rect 261435 154717 261447 154720
rect 261389 154711 261447 154717
rect 281077 154717 281089 154720
rect 281123 154717 281135 154751
rect 281077 154711 281135 154717
rect 281166 154708 281172 154760
rect 281224 154748 281230 154760
rect 295334 154748 295340 154760
rect 281224 154720 295340 154748
rect 281224 154708 281230 154720
rect 295334 154708 295340 154720
rect 295392 154708 295398 154760
rect 296717 154751 296775 154757
rect 296717 154717 296729 154751
rect 296763 154748 296775 154751
rect 297637 154751 297695 154757
rect 297637 154748 297649 154751
rect 296763 154720 297649 154748
rect 296763 154717 296775 154720
rect 296717 154711 296775 154717
rect 297637 154717 297649 154720
rect 297683 154717 297695 154751
rect 297637 154711 297695 154717
rect 297726 154708 297732 154760
rect 297784 154748 297790 154760
rect 314746 154748 314752 154760
rect 297784 154720 314752 154748
rect 297784 154708 297790 154720
rect 314746 154708 314752 154720
rect 314804 154708 314810 154760
rect 319162 154708 319168 154760
rect 319220 154748 319226 154760
rect 319220 154720 331076 154748
rect 319220 154708 319226 154720
rect 205634 154680 205640 154692
rect 197280 154652 205640 154680
rect 205634 154640 205640 154652
rect 205692 154640 205698 154692
rect 213825 154683 213883 154689
rect 213825 154649 213837 154683
rect 213871 154680 213883 154683
rect 214282 154680 214288 154692
rect 213871 154652 214288 154680
rect 213871 154649 213883 154652
rect 213825 154643 213883 154649
rect 214282 154640 214288 154652
rect 214340 154640 214346 154692
rect 223666 154640 223672 154692
rect 223724 154680 223730 154692
rect 269022 154680 269028 154692
rect 223724 154652 269028 154680
rect 223724 154640 223730 154652
rect 269022 154640 269028 154652
rect 269080 154640 269086 154692
rect 269301 154683 269359 154689
rect 269301 154649 269313 154683
rect 269347 154680 269359 154683
rect 283282 154680 283288 154692
rect 269347 154652 283288 154680
rect 269347 154649 269359 154652
rect 269301 154643 269359 154649
rect 283282 154640 283288 154652
rect 283340 154640 283346 154692
rect 285030 154640 285036 154692
rect 285088 154680 285094 154692
rect 301041 154683 301099 154689
rect 285088 154652 300808 154680
rect 285088 154640 285094 154652
rect 1302 154572 1308 154624
rect 1360 154612 1366 154624
rect 106182 154612 106188 154624
rect 1360 154584 106188 154612
rect 1360 154572 1366 154584
rect 106182 154572 106188 154584
rect 106240 154572 106246 154624
rect 110598 154572 110604 154624
rect 110656 154612 110662 154624
rect 110656 154584 175228 154612
rect 110656 154572 110662 154584
rect 67726 154504 67732 154556
rect 67784 154544 67790 154556
rect 164786 154544 164792 154556
rect 67784 154516 164792 154544
rect 67784 154504 67790 154516
rect 164786 154504 164792 154516
rect 164844 154504 164850 154556
rect 59906 154436 59912 154488
rect 59964 154476 59970 154488
rect 59964 154448 158576 154476
rect 59964 154436 59970 154448
rect 48222 154368 48228 154420
rect 48280 154408 48286 154420
rect 151998 154408 152004 154420
rect 48280 154380 152004 154408
rect 48280 154368 48286 154380
rect 151998 154368 152004 154380
rect 152056 154368 152062 154420
rect 158548 154408 158576 154448
rect 158714 154436 158720 154488
rect 158772 154476 158778 154488
rect 175200 154476 175228 154584
rect 175274 154572 175280 154624
rect 175332 154612 175338 154624
rect 183462 154612 183468 154624
rect 175332 154584 183468 154612
rect 175332 154572 175338 154584
rect 183462 154572 183468 154584
rect 183520 154572 183526 154624
rect 183646 154572 183652 154624
rect 183704 154612 183710 154624
rect 187053 154615 187111 154621
rect 187053 154612 187065 154615
rect 183704 154584 187065 154612
rect 183704 154572 183710 154584
rect 187053 154581 187065 154584
rect 187099 154581 187111 154615
rect 187053 154575 187111 154581
rect 187145 154615 187203 154621
rect 187145 154581 187157 154615
rect 187191 154612 187203 154615
rect 191742 154612 191748 154624
rect 187191 154584 191748 154612
rect 187191 154581 187203 154584
rect 187145 154575 187203 154581
rect 191742 154572 191748 154584
rect 191800 154572 191806 154624
rect 195241 154615 195299 154621
rect 195241 154581 195253 154615
rect 195287 154612 195299 154615
rect 242250 154612 242256 154624
rect 195287 154584 242256 154612
rect 195287 154581 195299 154584
rect 195241 154575 195299 154581
rect 242250 154572 242256 154584
rect 242308 154572 242314 154624
rect 243541 154615 243599 154621
rect 243541 154581 243553 154615
rect 243587 154612 243599 154615
rect 245933 154615 245991 154621
rect 245933 154612 245945 154615
rect 243587 154584 245945 154612
rect 243587 154581 243599 154584
rect 243541 154575 243599 154581
rect 245933 154581 245945 154584
rect 245979 154581 245991 154615
rect 245933 154575 245991 154581
rect 246022 154572 246028 154624
rect 246080 154612 246086 154624
rect 252649 154615 252707 154621
rect 246080 154584 252600 154612
rect 246080 154572 246086 154584
rect 179414 154504 179420 154556
rect 179472 154544 179478 154556
rect 184934 154544 184940 154556
rect 179472 154516 184940 154544
rect 179472 154504 179478 154516
rect 184934 154504 184940 154516
rect 184992 154504 184998 154556
rect 186314 154504 186320 154556
rect 186372 154544 186378 154556
rect 201494 154544 201500 154556
rect 186372 154516 201500 154544
rect 186372 154504 186378 154516
rect 201494 154504 201500 154516
rect 201552 154504 201558 154556
rect 202782 154504 202788 154556
rect 202840 154544 202846 154556
rect 248693 154547 248751 154553
rect 248693 154544 248705 154547
rect 202840 154516 248705 154544
rect 202840 154504 202846 154516
rect 248693 154513 248705 154516
rect 248739 154513 248751 154547
rect 248693 154507 248751 154513
rect 248877 154547 248935 154553
rect 248877 154513 248889 154547
rect 248923 154544 248935 154547
rect 249794 154544 249800 154556
rect 248923 154516 249800 154544
rect 248923 154513 248935 154516
rect 248877 154507 248935 154513
rect 249794 154504 249800 154516
rect 249852 154504 249858 154556
rect 252572 154544 252600 154584
rect 252649 154581 252661 154615
rect 252695 154612 252707 154615
rect 271782 154612 271788 154624
rect 252695 154584 271788 154612
rect 252695 154581 252707 154584
rect 252649 154575 252707 154581
rect 271782 154572 271788 154584
rect 271840 154572 271846 154624
rect 272521 154615 272579 154621
rect 272521 154581 272533 154615
rect 272567 154612 272579 154615
rect 288342 154612 288348 154624
rect 272567 154584 288348 154612
rect 272567 154581 272579 154584
rect 272521 154575 272579 154581
rect 288342 154572 288348 154584
rect 288400 154572 288406 154624
rect 288986 154572 288992 154624
rect 289044 154612 289050 154624
rect 289044 154584 300716 154612
rect 289044 154572 289050 154584
rect 281077 154547 281135 154553
rect 252572 154516 277394 154544
rect 158772 154448 175136 154476
rect 175200 154448 180794 154476
rect 158772 154436 158778 154448
rect 159634 154408 159640 154420
rect 158548 154380 159640 154408
rect 159634 154368 159640 154380
rect 159692 154368 159698 154420
rect 161661 154411 161719 154417
rect 161661 154377 161673 154411
rect 161707 154408 161719 154411
rect 171962 154408 171968 154420
rect 161707 154380 171968 154408
rect 161707 154377 161719 154380
rect 161661 154371 161719 154377
rect 171962 154368 171968 154380
rect 172020 154368 172026 154420
rect 175108 154408 175136 154448
rect 175274 154408 175280 154420
rect 175108 154380 175280 154408
rect 175274 154368 175280 154380
rect 175332 154368 175338 154420
rect 180766 154408 180794 154448
rect 184290 154436 184296 154488
rect 184348 154476 184354 154488
rect 198734 154476 198740 154488
rect 184348 154448 198740 154476
rect 184348 154436 184354 154448
rect 198734 154436 198740 154448
rect 198792 154436 198798 154488
rect 203150 154436 203156 154488
rect 203208 154476 203214 154488
rect 249061 154479 249119 154485
rect 249061 154476 249073 154479
rect 203208 154448 249073 154476
rect 203208 154436 203214 154448
rect 249061 154445 249073 154448
rect 249107 154445 249119 154479
rect 249061 154439 249119 154445
rect 255314 154436 255320 154488
rect 255372 154476 255378 154488
rect 261110 154476 261116 154488
rect 255372 154448 261116 154476
rect 255372 154436 255378 154448
rect 261110 154436 261116 154448
rect 261168 154436 261174 154488
rect 266354 154436 266360 154488
rect 266412 154476 266418 154488
rect 275370 154476 275376 154488
rect 266412 154448 275376 154476
rect 266412 154436 266418 154448
rect 275370 154436 275376 154448
rect 275428 154436 275434 154488
rect 277366 154476 277394 154516
rect 281077 154513 281089 154547
rect 281123 154544 281135 154547
rect 281534 154544 281540 154556
rect 281123 154516 281540 154544
rect 281123 154513 281135 154516
rect 281077 154507 281135 154513
rect 281534 154504 281540 154516
rect 281592 154504 281598 154556
rect 282914 154504 282920 154556
rect 282972 154544 282978 154556
rect 298830 154544 298836 154556
rect 282972 154516 298836 154544
rect 282972 154504 282978 154516
rect 298830 154504 298836 154516
rect 298888 154504 298894 154556
rect 284018 154476 284024 154488
rect 277366 154448 284024 154476
rect 284018 154436 284024 154448
rect 284076 154436 284082 154488
rect 285674 154436 285680 154488
rect 285732 154476 285738 154488
rect 300688 154476 300716 154584
rect 300780 154544 300808 154652
rect 301041 154649 301053 154683
rect 301087 154680 301099 154683
rect 303522 154680 303528 154692
rect 301087 154652 303528 154680
rect 301087 154649 301099 154652
rect 301041 154643 301099 154649
rect 303522 154640 303528 154652
rect 303580 154640 303586 154692
rect 303614 154640 303620 154692
rect 303672 154680 303678 154692
rect 318702 154680 318708 154692
rect 303672 154652 318708 154680
rect 303672 154640 303678 154652
rect 318702 154640 318708 154652
rect 318760 154640 318766 154692
rect 320174 154640 320180 154692
rect 320232 154680 320238 154692
rect 320232 154652 330984 154680
rect 320232 154640 320238 154652
rect 300857 154615 300915 154621
rect 300857 154581 300869 154615
rect 300903 154612 300915 154615
rect 303798 154612 303804 154624
rect 300903 154584 303804 154612
rect 300903 154581 300915 154584
rect 300857 154575 300915 154581
rect 303798 154572 303804 154584
rect 303856 154572 303862 154624
rect 304534 154572 304540 154624
rect 304592 154612 304598 154624
rect 311158 154612 311164 154624
rect 304592 154584 311164 154612
rect 304592 154572 304598 154584
rect 311158 154572 311164 154584
rect 311216 154572 311222 154624
rect 312354 154572 312360 154624
rect 312412 154612 312418 154624
rect 322934 154612 322940 154624
rect 312412 154584 322940 154612
rect 312412 154572 312418 154584
rect 322934 154572 322940 154584
rect 322992 154572 322998 154624
rect 300780 154516 306374 154544
rect 300854 154476 300860 154488
rect 285732 154448 296714 154476
rect 300688 154448 300860 154476
rect 285732 154436 285738 154448
rect 193398 154408 193404 154420
rect 180766 154380 193404 154408
rect 193398 154368 193404 154380
rect 193456 154368 193462 154420
rect 199286 154368 199292 154420
rect 199344 154408 199350 154420
rect 252646 154408 252652 154420
rect 199344 154380 252652 154408
rect 199344 154368 199350 154380
rect 252646 154368 252652 154380
rect 252704 154368 252710 154420
rect 253842 154368 253848 154420
rect 253900 154408 253906 154420
rect 289078 154408 289084 154420
rect 253900 154380 289084 154408
rect 253900 154368 253906 154380
rect 289078 154368 289084 154380
rect 289136 154368 289142 154420
rect 296686 154408 296714 154448
rect 300854 154436 300860 154448
rect 300912 154436 300918 154488
rect 301406 154408 301412 154420
rect 296686 154380 301412 154408
rect 301406 154368 301412 154380
rect 301464 154368 301470 154420
rect 44266 154300 44272 154352
rect 44324 154340 44330 154352
rect 149238 154340 149244 154352
rect 44324 154312 149244 154340
rect 44324 154300 44330 154312
rect 149238 154300 149244 154312
rect 149296 154300 149302 154352
rect 164789 154343 164847 154349
rect 164789 154340 164801 154343
rect 161446 154312 164801 154340
rect 40402 154232 40408 154284
rect 40460 154272 40466 154284
rect 146570 154272 146576 154284
rect 40460 154244 146576 154272
rect 40460 154232 40466 154244
rect 146570 154232 146576 154244
rect 146628 154232 146634 154284
rect 149054 154232 149060 154284
rect 149112 154272 149118 154284
rect 161446 154272 161474 154312
rect 164789 154309 164801 154312
rect 164835 154309 164847 154343
rect 164789 154303 164847 154309
rect 164878 154300 164884 154352
rect 164936 154340 164942 154352
rect 185670 154340 185676 154352
rect 164936 154312 185676 154340
rect 164936 154300 164942 154312
rect 185670 154300 185676 154312
rect 185728 154300 185734 154352
rect 186406 154300 186412 154352
rect 186464 154340 186470 154352
rect 187789 154343 187847 154349
rect 187789 154340 187801 154343
rect 186464 154312 187801 154340
rect 186464 154300 186470 154312
rect 187789 154309 187801 154312
rect 187835 154309 187847 154343
rect 187789 154303 187847 154309
rect 192478 154300 192484 154352
rect 192536 154340 192542 154352
rect 243357 154343 243415 154349
rect 243357 154340 243369 154343
rect 192536 154312 243369 154340
rect 192536 154300 192542 154312
rect 243357 154309 243369 154312
rect 243403 154309 243415 154343
rect 243357 154303 243415 154309
rect 243449 154343 243507 154349
rect 243449 154309 243461 154343
rect 243495 154340 243507 154343
rect 247402 154340 247408 154352
rect 243495 154312 247408 154340
rect 243495 154309 243507 154312
rect 243449 154303 243507 154309
rect 247402 154300 247408 154312
rect 247460 154300 247466 154352
rect 248785 154343 248843 154349
rect 248785 154309 248797 154343
rect 248831 154340 248843 154343
rect 249978 154340 249984 154352
rect 248831 154312 249984 154340
rect 248831 154309 248843 154312
rect 248785 154303 248843 154309
rect 249978 154300 249984 154312
rect 250036 154300 250042 154352
rect 254854 154300 254860 154352
rect 254912 154340 254918 154352
rect 289814 154340 289820 154352
rect 254912 154312 289820 154340
rect 254912 154300 254918 154312
rect 289814 154300 289820 154312
rect 289872 154300 289878 154352
rect 292574 154300 292580 154352
rect 292632 154340 292638 154352
rect 299474 154340 299480 154352
rect 292632 154312 299480 154340
rect 292632 154300 292638 154312
rect 299474 154300 299480 154312
rect 299532 154300 299538 154352
rect 306346 154340 306374 154516
rect 330956 154476 330984 154652
rect 331048 154544 331076 154720
rect 340598 154708 340604 154760
rect 340656 154748 340662 154760
rect 340656 154720 346440 154748
rect 340656 154708 340662 154720
rect 339678 154640 339684 154692
rect 339736 154680 339742 154692
rect 346302 154680 346308 154692
rect 339736 154652 346308 154680
rect 339736 154640 339742 154652
rect 346302 154640 346308 154652
rect 346360 154640 346366 154692
rect 336734 154572 336740 154624
rect 336792 154612 336798 154624
rect 336792 154584 343588 154612
rect 336792 154572 336798 154584
rect 332594 154544 332600 154556
rect 331048 154516 332600 154544
rect 332594 154504 332600 154516
rect 332652 154504 332658 154556
rect 343560 154544 343588 154584
rect 344370 154544 344376 154556
rect 343560 154516 344376 154544
rect 344370 154504 344376 154516
rect 344428 154504 344434 154556
rect 346412 154544 346440 154720
rect 399478 154708 399484 154760
rect 399536 154748 399542 154760
rect 402946 154748 402974 154788
rect 399536 154720 402974 154748
rect 399536 154708 399542 154720
rect 407022 154708 407028 154760
rect 407080 154748 407086 154760
rect 407868 154748 407896 154924
rect 417421 154921 417433 154924
rect 417467 154921 417479 154955
rect 417421 154915 417479 154921
rect 417786 154912 417792 154964
rect 417844 154952 417850 154964
rect 445846 154952 445852 154964
rect 417844 154924 445852 154952
rect 417844 154912 417850 154924
rect 445846 154912 445852 154924
rect 445904 154912 445910 154964
rect 464614 154912 464620 154964
rect 464672 154952 464678 154964
rect 516042 154952 516048 154964
rect 464672 154924 516048 154952
rect 464672 154912 464678 154924
rect 516042 154912 516048 154924
rect 516100 154912 516106 154964
rect 417329 154887 417387 154893
rect 417329 154884 417341 154887
rect 407080 154720 407896 154748
rect 407960 154856 417341 154884
rect 407080 154708 407086 154720
rect 352282 154640 352288 154692
rect 352340 154680 352346 154692
rect 353386 154680 353392 154692
rect 352340 154652 353392 154680
rect 352340 154640 352346 154652
rect 353386 154640 353392 154652
rect 353444 154640 353450 154692
rect 406102 154640 406108 154692
rect 406160 154680 406166 154692
rect 407960 154680 407988 154856
rect 417329 154853 417341 154856
rect 417375 154853 417387 154887
rect 441982 154884 441988 154896
rect 417329 154847 417387 154853
rect 417436 154856 441988 154884
rect 413830 154776 413836 154828
rect 413888 154816 413894 154828
rect 417053 154819 417111 154825
rect 417053 154816 417065 154819
rect 413888 154788 417065 154816
rect 413888 154776 413894 154788
rect 417053 154785 417065 154788
rect 417099 154785 417111 154819
rect 417053 154779 417111 154785
rect 415210 154708 415216 154760
rect 415268 154748 415274 154760
rect 417436 154748 417464 154856
rect 441982 154844 441988 154856
rect 442040 154844 442046 154896
rect 463326 154844 463332 154896
rect 463384 154884 463390 154896
rect 514110 154884 514116 154896
rect 463384 154856 514116 154884
rect 463384 154844 463390 154856
rect 514110 154844 514116 154856
rect 514168 154844 514174 154896
rect 417970 154776 417976 154828
rect 418028 154816 418034 154828
rect 444926 154816 444932 154828
rect 418028 154788 444932 154816
rect 418028 154776 418034 154788
rect 444926 154776 444932 154788
rect 444984 154776 444990 154828
rect 459462 154776 459468 154828
rect 459520 154816 459526 154828
rect 508222 154816 508228 154828
rect 459520 154788 508228 154816
rect 459520 154776 459526 154788
rect 508222 154776 508228 154788
rect 508280 154776 508286 154828
rect 415268 154720 417464 154748
rect 417513 154751 417571 154757
rect 415268 154708 415274 154720
rect 417513 154717 417525 154751
rect 417559 154748 417571 154751
rect 438118 154748 438124 154760
rect 417559 154720 438124 154748
rect 417559 154717 417571 154720
rect 417513 154711 417571 154717
rect 438118 154708 438124 154720
rect 438176 154708 438182 154760
rect 460106 154708 460112 154760
rect 460164 154748 460170 154760
rect 509234 154748 509240 154760
rect 460164 154720 509240 154748
rect 460164 154708 460170 154720
rect 509234 154708 509240 154720
rect 509292 154708 509298 154760
rect 406160 154652 407988 154680
rect 406160 154640 406166 154652
rect 411990 154640 411996 154692
rect 412048 154680 412054 154692
rect 437106 154680 437112 154692
rect 412048 154652 437112 154680
rect 412048 154640 412054 154652
rect 437106 154640 437112 154652
rect 437164 154640 437170 154692
rect 461394 154640 461400 154692
rect 461452 154680 461458 154692
rect 511166 154680 511172 154692
rect 461452 154652 511172 154680
rect 461452 154640 461458 154652
rect 511166 154640 511172 154652
rect 511224 154640 511230 154692
rect 346486 154572 346492 154624
rect 346544 154612 346550 154624
rect 346544 154584 348372 154612
rect 346544 154572 346550 154584
rect 347038 154544 347044 154556
rect 346412 154516 347044 154544
rect 347038 154504 347044 154516
rect 347096 154504 347102 154556
rect 333238 154476 333244 154488
rect 330956 154448 333244 154476
rect 333238 154436 333244 154448
rect 333296 154436 333302 154488
rect 340966 154436 340972 154488
rect 341024 154476 341030 154488
rect 343726 154476 343732 154488
rect 341024 154448 343732 154476
rect 341024 154436 341030 154448
rect 343726 154436 343732 154448
rect 343784 154436 343790 154488
rect 309870 154340 309876 154352
rect 306346 154312 309876 154340
rect 309870 154300 309876 154312
rect 309928 154300 309934 154352
rect 167454 154272 167460 154284
rect 149112 154244 161474 154272
rect 161952 154244 167460 154272
rect 149112 154232 149118 154244
rect 35526 154164 35532 154216
rect 35584 154204 35590 154216
rect 143534 154204 143540 154216
rect 35584 154176 143540 154204
rect 35584 154164 35590 154176
rect 143534 154164 143540 154176
rect 143592 154164 143598 154216
rect 144730 154164 144736 154216
rect 144788 154204 144794 154216
rect 161842 154204 161848 154216
rect 144788 154176 161848 154204
rect 144788 154164 144794 154176
rect 161842 154164 161848 154176
rect 161900 154164 161906 154216
rect 32582 154096 32588 154148
rect 32640 154136 32646 154148
rect 141418 154136 141424 154148
rect 32640 154108 141424 154136
rect 32640 154096 32646 154108
rect 141418 154096 141424 154108
rect 141476 154096 141482 154148
rect 144822 154096 144828 154148
rect 144880 154136 144886 154148
rect 161952 154136 161980 154244
rect 167454 154232 167460 154244
rect 167512 154232 167518 154284
rect 168374 154232 168380 154284
rect 168432 154272 168438 154284
rect 179782 154272 179788 154284
rect 168432 154244 179788 154272
rect 168432 154232 168438 154244
rect 179782 154232 179788 154244
rect 179840 154232 179846 154284
rect 183370 154232 183376 154284
rect 183428 154272 183434 154284
rect 240226 154272 240232 154284
rect 183428 154244 240232 154272
rect 183428 154232 183434 154244
rect 240226 154232 240232 154244
rect 240284 154232 240290 154284
rect 247034 154232 247040 154284
rect 247092 154272 247098 154284
rect 284478 154272 284484 154284
rect 247092 154244 284484 154272
rect 247092 154232 247098 154244
rect 284478 154232 284484 154244
rect 284536 154232 284542 154284
rect 289262 154232 289268 154284
rect 289320 154272 289326 154284
rect 303982 154272 303988 154284
rect 289320 154244 303988 154272
rect 289320 154232 289326 154244
rect 303982 154232 303988 154244
rect 304040 154232 304046 154284
rect 304994 154232 305000 154284
rect 305052 154272 305058 154284
rect 315022 154272 315028 154284
rect 305052 154244 315028 154272
rect 305052 154232 305058 154244
rect 315022 154232 315028 154244
rect 315080 154232 315086 154284
rect 348344 154272 348372 154584
rect 348418 154572 348424 154624
rect 348476 154612 348482 154624
rect 348476 154584 349292 154612
rect 348476 154572 348482 154584
rect 349264 154340 349292 154584
rect 349338 154572 349344 154624
rect 349396 154612 349402 154624
rect 349396 154584 350304 154612
rect 349396 154572 349402 154584
rect 350276 154544 350304 154584
rect 350350 154572 350356 154624
rect 350408 154612 350414 154624
rect 350408 154584 351316 154612
rect 350408 154572 350414 154584
rect 350276 154516 351224 154544
rect 351196 154408 351224 154516
rect 351288 154476 351316 154584
rect 351362 154572 351368 154624
rect 351420 154612 351426 154624
rect 367922 154612 367928 154624
rect 351420 154584 353248 154612
rect 351420 154572 351426 154584
rect 353220 154544 353248 154584
rect 365732 154584 367928 154612
rect 354122 154544 354128 154556
rect 353220 154516 354128 154544
rect 354122 154504 354128 154516
rect 354180 154504 354186 154556
rect 361482 154504 361488 154556
rect 361540 154544 361546 154556
rect 362034 154544 362040 154556
rect 361540 154516 362040 154544
rect 361540 154504 361546 154516
rect 362034 154504 362040 154516
rect 362092 154504 362098 154556
rect 362586 154504 362592 154556
rect 362644 154544 362650 154556
rect 363046 154544 363052 154556
rect 362644 154516 363052 154544
rect 362644 154504 362650 154516
rect 363046 154504 363052 154516
rect 363104 154504 363110 154556
rect 365622 154504 365628 154556
rect 365680 154544 365686 154556
rect 365732 154544 365760 154584
rect 367922 154572 367928 154584
rect 367980 154572 367986 154624
rect 368842 154612 368848 154624
rect 368032 154584 368848 154612
rect 365680 154516 365760 154544
rect 365680 154504 365686 154516
rect 366450 154504 366456 154556
rect 366508 154544 366514 154556
rect 368032 154544 368060 154584
rect 368842 154572 368848 154584
rect 368900 154572 368906 154624
rect 370866 154612 370872 154624
rect 369964 154584 370872 154612
rect 366508 154516 368060 154544
rect 366508 154504 366514 154516
rect 353478 154476 353484 154488
rect 351288 154448 353484 154476
rect 353478 154436 353484 154448
rect 353536 154436 353542 154488
rect 362862 154436 362868 154488
rect 362920 154476 362926 154488
rect 363966 154476 363972 154488
rect 362920 154448 363972 154476
rect 362920 154436 362926 154448
rect 363966 154436 363972 154448
rect 364024 154436 364030 154488
rect 367002 154436 367008 154488
rect 367060 154476 367066 154488
rect 369854 154476 369860 154488
rect 367060 154448 369860 154476
rect 367060 154436 367066 154448
rect 369854 154436 369860 154448
rect 369912 154436 369918 154488
rect 352834 154408 352840 154420
rect 351196 154380 352840 154408
rect 352834 154368 352840 154380
rect 352892 154368 352898 154420
rect 367738 154368 367744 154420
rect 367796 154408 367802 154420
rect 369964 154408 369992 154584
rect 370866 154572 370872 154584
rect 370924 154572 370930 154624
rect 381538 154612 381544 154624
rect 379532 154584 381544 154612
rect 374914 154504 374920 154556
rect 374972 154544 374978 154556
rect 379532 154544 379560 154584
rect 381538 154572 381544 154584
rect 381596 154572 381602 154624
rect 383470 154612 383476 154624
rect 381648 154584 383476 154612
rect 374972 154516 379560 154544
rect 374972 154504 374978 154516
rect 372982 154436 372988 154488
rect 373040 154476 373046 154488
rect 378594 154476 378600 154488
rect 373040 154448 378600 154476
rect 373040 154436 373046 154448
rect 378594 154436 378600 154448
rect 378652 154436 378658 154488
rect 367796 154380 369992 154408
rect 367796 154368 367802 154380
rect 375190 154368 375196 154420
rect 375248 154408 375254 154420
rect 379698 154408 379704 154420
rect 375248 154380 379704 154408
rect 375248 154368 375254 154380
rect 379698 154368 379704 154380
rect 379756 154368 379762 154420
rect 352098 154340 352104 154352
rect 349264 154312 352104 154340
rect 352098 154300 352104 154312
rect 352156 154300 352162 154352
rect 368382 154300 368388 154352
rect 368440 154340 368446 154352
rect 371786 154340 371792 154352
rect 368440 154312 371792 154340
rect 368440 154300 368446 154312
rect 371786 154300 371792 154312
rect 371844 154300 371850 154352
rect 376202 154300 376208 154352
rect 376260 154340 376266 154352
rect 381648 154340 381676 154584
rect 383470 154572 383476 154584
rect 383528 154572 383534 154624
rect 403986 154572 403992 154624
rect 404044 154612 404050 154624
rect 405918 154612 405924 154624
rect 404044 154584 405924 154612
rect 404044 154572 404050 154584
rect 405918 154572 405924 154584
rect 405976 154572 405982 154624
rect 409414 154572 409420 154624
rect 409472 154612 409478 154624
rect 433242 154612 433248 154624
rect 409472 154584 433248 154612
rect 409472 154572 409478 154584
rect 433242 154572 433248 154584
rect 433300 154572 433306 154624
rect 457530 154572 457536 154624
rect 457588 154612 457594 154624
rect 505370 154612 505376 154624
rect 457588 154584 505376 154612
rect 457588 154572 457594 154584
rect 505370 154572 505376 154584
rect 505428 154572 505434 154624
rect 578418 154612 578424 154624
rect 578379 154584 578424 154612
rect 578418 154572 578424 154584
rect 578476 154572 578482 154624
rect 382090 154504 382096 154556
rect 382148 154544 382154 154556
rect 392302 154544 392308 154556
rect 382148 154516 392308 154544
rect 382148 154504 382154 154516
rect 392302 154504 392308 154516
rect 392360 154504 392366 154556
rect 395982 154504 395988 154556
rect 396040 154544 396046 154556
rect 411254 154544 411260 154556
rect 396040 154516 411260 154544
rect 396040 154504 396046 154516
rect 411254 154504 411260 154516
rect 411312 154504 411318 154556
rect 415854 154504 415860 154556
rect 415912 154544 415918 154556
rect 442994 154544 443000 154556
rect 415912 154516 443000 154544
rect 415912 154504 415918 154516
rect 442994 154504 443000 154516
rect 443052 154504 443058 154556
rect 471790 154504 471796 154556
rect 471848 154544 471854 154556
rect 526806 154544 526812 154556
rect 471848 154516 526812 154544
rect 471848 154504 471854 154516
rect 526806 154504 526812 154516
rect 526864 154504 526870 154556
rect 384022 154436 384028 154488
rect 384080 154476 384086 154488
rect 395154 154476 395160 154488
rect 384080 154448 395160 154476
rect 384080 154436 384086 154448
rect 395154 154436 395160 154448
rect 395212 154436 395218 154488
rect 395706 154436 395712 154488
rect 395764 154476 395770 154488
rect 411346 154476 411352 154488
rect 395764 154448 411352 154476
rect 395764 154436 395770 154448
rect 411346 154436 411352 154448
rect 411404 154436 411410 154488
rect 416498 154436 416504 154488
rect 416556 154476 416562 154488
rect 443914 154476 443920 154488
rect 416556 154448 443920 154476
rect 416556 154436 416562 154448
rect 443914 154436 443920 154448
rect 443972 154436 443978 154488
rect 500402 154436 500408 154488
rect 500460 154476 500466 154488
rect 554774 154476 554780 154488
rect 500460 154448 554780 154476
rect 500460 154436 500466 154448
rect 554774 154436 554780 154448
rect 554832 154436 554838 154488
rect 384666 154368 384672 154420
rect 384724 154408 384730 154420
rect 396166 154408 396172 154420
rect 384724 154380 396172 154408
rect 384724 154368 384730 154380
rect 396166 154368 396172 154380
rect 396224 154368 396230 154420
rect 396994 154368 397000 154420
rect 397052 154408 397058 154420
rect 413278 154408 413284 154420
rect 397052 154380 413284 154408
rect 397052 154368 397058 154380
rect 413278 154368 413284 154380
rect 413336 154368 413342 154420
rect 419166 154368 419172 154420
rect 419224 154408 419230 154420
rect 447870 154408 447876 154420
rect 419224 154380 447876 154408
rect 419224 154368 419230 154380
rect 447870 154368 447876 154380
rect 447928 154368 447934 154420
rect 482186 154368 482192 154420
rect 482244 154408 482250 154420
rect 542262 154408 542268 154420
rect 482244 154380 542268 154408
rect 482244 154368 482250 154380
rect 542262 154368 542268 154380
rect 542320 154368 542326 154420
rect 376260 154312 381676 154340
rect 376260 154300 376266 154312
rect 385954 154300 385960 154352
rect 386012 154340 386018 154352
rect 398098 154340 398104 154352
rect 386012 154312 398104 154340
rect 386012 154300 386018 154312
rect 398098 154300 398104 154312
rect 398156 154300 398162 154352
rect 398282 154300 398288 154352
rect 398340 154340 398346 154352
rect 414106 154340 414112 154352
rect 398340 154312 414112 154340
rect 398340 154300 398346 154312
rect 414106 154300 414112 154312
rect 414164 154300 414170 154352
rect 421742 154300 421748 154352
rect 421800 154340 421806 154352
rect 451734 154340 451740 154352
rect 421800 154312 451740 154340
rect 421800 154300 421806 154312
rect 451734 154300 451740 154312
rect 451792 154300 451798 154352
rect 486142 154300 486148 154352
rect 486200 154340 486206 154352
rect 546494 154340 546500 154352
rect 486200 154312 546500 154340
rect 486200 154300 486206 154312
rect 546494 154300 546500 154312
rect 546552 154300 546558 154352
rect 548518 154300 548524 154352
rect 548576 154340 548582 154352
rect 575566 154340 575572 154352
rect 548576 154312 575572 154340
rect 548576 154300 548582 154312
rect 575566 154300 575572 154312
rect 575624 154300 575630 154352
rect 350810 154272 350816 154284
rect 348344 154244 350816 154272
rect 350810 154232 350816 154244
rect 350868 154232 350874 154284
rect 369670 154232 369676 154284
rect 369728 154272 369734 154284
rect 373718 154272 373724 154284
rect 369728 154244 373724 154272
rect 369728 154232 369734 154244
rect 373718 154232 373724 154244
rect 373776 154232 373782 154284
rect 384942 154232 384948 154284
rect 385000 154272 385006 154284
rect 397178 154272 397184 154284
rect 385000 154244 397184 154272
rect 385000 154232 385006 154244
rect 397178 154232 397184 154244
rect 397236 154232 397242 154284
rect 397270 154232 397276 154284
rect 397328 154272 397334 154284
rect 415670 154272 415676 154284
rect 397328 154244 415676 154272
rect 397328 154232 397334 154244
rect 415670 154232 415676 154244
rect 415728 154232 415734 154284
rect 424318 154232 424324 154284
rect 424376 154272 424382 154284
rect 455598 154272 455604 154284
rect 424376 154244 455604 154272
rect 424376 154232 424382 154244
rect 455598 154232 455604 154244
rect 455656 154232 455662 154284
rect 487062 154232 487068 154284
rect 487120 154272 487126 154284
rect 550174 154272 550180 154284
rect 487120 154244 550180 154272
rect 487120 154232 487126 154244
rect 550174 154232 550180 154244
rect 550232 154232 550238 154284
rect 162118 154164 162124 154216
rect 162176 154204 162182 154216
rect 178034 154204 178040 154216
rect 162176 154176 178040 154204
rect 162176 154164 162182 154176
rect 178034 154164 178040 154176
rect 178092 154164 178098 154216
rect 179138 154164 179144 154216
rect 179196 154204 179202 154216
rect 237650 154204 237656 154216
rect 179196 154176 237656 154204
rect 179196 154164 179202 154176
rect 237650 154164 237656 154176
rect 237708 154164 237714 154216
rect 241422 154164 241428 154216
rect 241480 154204 241486 154216
rect 279326 154204 279332 154216
rect 241480 154176 279332 154204
rect 241480 154164 241486 154176
rect 279326 154164 279332 154176
rect 279384 154164 279390 154216
rect 281997 154207 282055 154213
rect 281997 154173 282009 154207
rect 282043 154204 282055 154207
rect 285674 154204 285680 154216
rect 282043 154176 285680 154204
rect 282043 154173 282055 154176
rect 281997 154167 282055 154173
rect 285674 154164 285680 154176
rect 285732 154164 285738 154216
rect 290826 154164 290832 154216
rect 290884 154204 290890 154216
rect 306650 154204 306656 154216
rect 290884 154176 306656 154204
rect 290884 154164 290890 154176
rect 306650 154164 306656 154176
rect 306708 154164 306714 154216
rect 308398 154164 308404 154216
rect 308456 154204 308462 154216
rect 317690 154204 317696 154216
rect 308456 154176 317696 154204
rect 308456 154164 308462 154176
rect 317690 154164 317696 154176
rect 317748 154164 317754 154216
rect 347590 154164 347596 154216
rect 347648 154204 347654 154216
rect 350166 154204 350172 154216
rect 347648 154176 350172 154204
rect 347648 154164 347654 154176
rect 350166 154164 350172 154176
rect 350224 154164 350230 154216
rect 372338 154164 372344 154216
rect 372396 154204 372402 154216
rect 377674 154204 377680 154216
rect 372396 154176 377680 154204
rect 372396 154164 372402 154176
rect 377674 154164 377680 154176
rect 377732 154164 377738 154216
rect 386230 154164 386236 154216
rect 386288 154204 386294 154216
rect 398742 154204 398748 154216
rect 386288 154176 398748 154204
rect 386288 154164 386294 154176
rect 398742 154164 398748 154176
rect 398800 154164 398806 154216
rect 400122 154164 400128 154216
rect 400180 154204 400186 154216
rect 419534 154204 419540 154216
rect 400180 154176 419540 154204
rect 400180 154164 400186 154176
rect 419534 154164 419540 154176
rect 419592 154164 419598 154216
rect 426894 154164 426900 154216
rect 426952 154204 426958 154216
rect 459554 154204 459560 154216
rect 426952 154176 459560 154204
rect 426952 154164 426958 154176
rect 459554 154164 459560 154176
rect 459612 154164 459618 154216
rect 489638 154164 489644 154216
rect 489696 154204 489702 154216
rect 554038 154204 554044 154216
rect 489696 154176 554044 154204
rect 489696 154164 489702 154176
rect 554038 154164 554044 154176
rect 554096 154164 554102 154216
rect 144880 154108 161980 154136
rect 164789 154139 164847 154145
rect 144880 154096 144886 154108
rect 164789 154105 164801 154139
rect 164835 154136 164847 154139
rect 166994 154136 167000 154148
rect 164835 154108 167000 154136
rect 164835 154105 164847 154108
rect 164789 154099 164847 154105
rect 166994 154096 167000 154108
rect 167052 154096 167058 154148
rect 172422 154096 172428 154148
rect 172480 154136 172486 154148
rect 232498 154136 232504 154148
rect 172480 154108 232504 154136
rect 172480 154096 172486 154108
rect 232498 154096 232504 154108
rect 232556 154096 232562 154148
rect 235350 154096 235356 154148
rect 235408 154136 235414 154148
rect 235408 154108 275968 154136
rect 235408 154096 235414 154108
rect 28718 154028 28724 154080
rect 28776 154068 28782 154080
rect 138842 154068 138848 154080
rect 28776 154040 138848 154068
rect 28776 154028 28782 154040
rect 138842 154028 138848 154040
rect 138900 154028 138906 154080
rect 140774 154028 140780 154080
rect 140832 154068 140838 154080
rect 156966 154068 156972 154080
rect 140832 154040 156972 154068
rect 140832 154028 140838 154040
rect 156966 154028 156972 154040
rect 157024 154028 157030 154080
rect 157334 154028 157340 154080
rect 157392 154068 157398 154080
rect 224954 154068 224960 154080
rect 157392 154040 224960 154068
rect 157392 154028 157398 154040
rect 224954 154028 224960 154040
rect 225012 154028 225018 154080
rect 233142 154028 233148 154080
rect 233200 154068 233206 154080
rect 273438 154068 273444 154080
rect 233200 154040 273444 154068
rect 233200 154028 233206 154040
rect 273438 154028 273444 154040
rect 273496 154028 273502 154080
rect 275940 154068 275968 154108
rect 276014 154096 276020 154148
rect 276072 154136 276078 154148
rect 285766 154136 285772 154148
rect 276072 154108 285772 154136
rect 276072 154096 276078 154108
rect 285766 154096 285772 154108
rect 285824 154096 285830 154148
rect 291746 154096 291752 154148
rect 291804 154136 291810 154148
rect 309226 154136 309232 154148
rect 291804 154108 309232 154136
rect 291804 154096 291810 154108
rect 309226 154096 309232 154108
rect 309284 154096 309290 154148
rect 309318 154096 309324 154148
rect 309376 154136 309382 154148
rect 320266 154136 320272 154148
rect 309376 154108 320272 154136
rect 309376 154096 309382 154108
rect 320266 154096 320272 154108
rect 320324 154096 320330 154148
rect 381446 154096 381452 154148
rect 381504 154136 381510 154148
rect 387334 154136 387340 154148
rect 381504 154108 387340 154136
rect 381504 154096 381510 154108
rect 387334 154096 387340 154108
rect 387392 154096 387398 154148
rect 390462 154096 390468 154148
rect 390520 154136 390526 154148
rect 401594 154136 401600 154148
rect 390520 154108 401600 154136
rect 390520 154096 390526 154108
rect 401594 154096 401600 154108
rect 401652 154096 401658 154148
rect 403526 154096 403532 154148
rect 403584 154136 403590 154148
rect 424410 154136 424416 154148
rect 403584 154108 424416 154136
rect 403584 154096 403590 154108
rect 424410 154096 424416 154108
rect 424468 154096 424474 154148
rect 429562 154096 429568 154148
rect 429620 154136 429626 154148
rect 463418 154136 463424 154148
rect 429620 154108 463424 154136
rect 429620 154096 429626 154108
rect 463418 154096 463424 154108
rect 463476 154096 463482 154148
rect 474458 154096 474464 154148
rect 474516 154136 474522 154148
rect 480070 154136 480076 154148
rect 474516 154108 480076 154136
rect 474516 154096 474522 154108
rect 480070 154096 480076 154108
rect 480128 154096 480134 154148
rect 492582 154096 492588 154148
rect 492640 154136 492646 154148
rect 557994 154136 558000 154148
rect 492640 154108 558000 154136
rect 492640 154096 492646 154108
rect 557994 154096 558000 154108
rect 558052 154096 558058 154148
rect 276658 154068 276664 154080
rect 275940 154040 276664 154068
rect 276658 154028 276664 154040
rect 276716 154028 276722 154080
rect 276750 154028 276756 154080
rect 276808 154068 276814 154080
rect 291194 154068 291200 154080
rect 276808 154040 291200 154068
rect 276808 154028 276814 154040
rect 291194 154028 291200 154040
rect 291252 154028 291258 154080
rect 291838 154028 291844 154080
rect 291896 154068 291902 154080
rect 314654 154068 314660 154080
rect 291896 154040 314660 154068
rect 291896 154028 291902 154040
rect 314654 154028 314660 154040
rect 314712 154028 314718 154080
rect 387702 154028 387708 154080
rect 387760 154068 387766 154080
rect 398926 154068 398932 154080
rect 387760 154040 398932 154068
rect 387760 154028 387766 154040
rect 398926 154028 398932 154040
rect 398984 154028 398990 154080
rect 402698 154028 402704 154080
rect 402756 154068 402762 154080
rect 423490 154068 423496 154080
rect 402756 154040 423496 154068
rect 402756 154028 402762 154040
rect 423490 154028 423496 154040
rect 423548 154028 423554 154080
rect 431770 154028 431776 154080
rect 431828 154068 431834 154080
rect 467282 154068 467288 154080
rect 431828 154040 467288 154068
rect 431828 154028 431834 154040
rect 467282 154028 467288 154040
rect 467340 154028 467346 154080
rect 495250 154028 495256 154080
rect 495308 154068 495314 154080
rect 561582 154068 561588 154080
rect 495308 154040 561588 154068
rect 495308 154028 495314 154040
rect 561582 154028 561588 154040
rect 561640 154028 561646 154080
rect 20898 153960 20904 154012
rect 20956 154000 20962 154012
rect 133874 154000 133880 154012
rect 20956 153972 133880 154000
rect 20956 153960 20962 153972
rect 133874 153960 133880 153972
rect 133932 153960 133938 154012
rect 135162 153960 135168 154012
rect 135220 154000 135226 154012
rect 137925 154003 137983 154009
rect 137925 154000 137937 154003
rect 135220 153972 137937 154000
rect 135220 153960 135226 153972
rect 137925 153969 137937 153972
rect 137971 153969 137983 154003
rect 137925 153963 137983 153969
rect 138014 153960 138020 154012
rect 138072 154000 138078 154012
rect 145926 154000 145932 154012
rect 138072 153972 145932 154000
rect 138072 153960 138078 153972
rect 145926 153960 145932 153972
rect 145984 153960 145990 154012
rect 153102 153960 153108 154012
rect 153160 154000 153166 154012
rect 219618 154000 219624 154012
rect 153160 153972 219624 154000
rect 153160 153960 153166 153972
rect 219618 153960 219624 153972
rect 219676 153960 219682 154012
rect 227530 153960 227536 154012
rect 227588 154000 227594 154012
rect 271506 154000 271512 154012
rect 227588 153972 271512 154000
rect 227588 153960 227594 153972
rect 271506 153960 271512 153972
rect 271564 153960 271570 154012
rect 274634 153960 274640 154012
rect 274692 154000 274698 154012
rect 288434 154000 288440 154012
rect 274692 153972 288440 154000
rect 274692 153960 274698 153972
rect 288434 153960 288440 153972
rect 288492 153960 288498 154012
rect 289906 153960 289912 154012
rect 289964 154000 289970 154012
rect 313274 154000 313280 154012
rect 289964 153972 313280 154000
rect 289964 153960 289970 153972
rect 313274 153960 313280 153972
rect 313332 153960 313338 154012
rect 369026 153960 369032 154012
rect 369084 154000 369090 154012
rect 372798 154000 372804 154012
rect 369084 153972 372804 154000
rect 369084 153960 369090 153972
rect 372798 153960 372804 153972
rect 372856 153960 372862 154012
rect 373902 153960 373908 154012
rect 373960 154000 373966 154012
rect 378134 154000 378140 154012
rect 373960 153972 378140 154000
rect 373960 153960 373966 153972
rect 378134 153960 378140 153972
rect 378192 153960 378198 154012
rect 388530 153960 388536 154012
rect 388588 154000 388594 154012
rect 400214 154000 400220 154012
rect 388588 153972 400220 154000
rect 388588 153960 388594 153972
rect 400214 153960 400220 153972
rect 400272 153960 400278 154012
rect 405458 153960 405464 154012
rect 405516 154000 405522 154012
rect 427354 154000 427360 154012
rect 405516 153972 427360 154000
rect 405516 153960 405522 153972
rect 427354 153960 427360 153972
rect 427412 153960 427418 154012
rect 432782 153960 432788 154012
rect 432840 154000 432846 154012
rect 468294 154000 468300 154012
rect 432840 153972 468300 154000
rect 432840 153960 432846 153972
rect 468294 153960 468300 153972
rect 468352 153960 468358 154012
rect 497826 153960 497832 154012
rect 497884 154000 497890 154012
rect 565722 154000 565728 154012
rect 497884 153972 565728 154000
rect 497884 153960 497890 153972
rect 565722 153960 565728 153972
rect 565780 153960 565786 154012
rect 13078 153892 13084 153944
rect 13136 153932 13142 153944
rect 128354 153932 128360 153944
rect 13136 153904 128360 153932
rect 13136 153892 13142 153904
rect 128354 153892 128360 153904
rect 128412 153892 128418 153944
rect 135530 153932 135536 153944
rect 128464 153904 135536 153932
rect 9214 153824 9220 153876
rect 9272 153864 9278 153876
rect 125778 153864 125784 153876
rect 9272 153836 125784 153864
rect 9272 153824 9278 153836
rect 125778 153824 125784 153836
rect 125836 153824 125842 153876
rect 126054 153824 126060 153876
rect 126112 153864 126118 153876
rect 127437 153867 127495 153873
rect 127437 153864 127449 153867
rect 126112 153836 127449 153864
rect 126112 153824 126118 153836
rect 127437 153833 127449 153836
rect 127483 153833 127495 153867
rect 127437 153827 127495 153833
rect 127529 153867 127587 153873
rect 127529 153833 127541 153867
rect 127575 153864 127587 153867
rect 128464 153864 128492 153904
rect 135530 153892 135536 153904
rect 135588 153892 135594 153944
rect 136726 153892 136732 153944
rect 136784 153932 136790 153944
rect 140774 153932 140780 153944
rect 136784 153904 140780 153932
rect 136784 153892 136790 153904
rect 140774 153892 140780 153904
rect 140832 153892 140838 153944
rect 140866 153892 140872 153944
rect 140924 153932 140930 153944
rect 143994 153932 144000 153944
rect 140924 153904 144000 153932
rect 140924 153892 140930 153904
rect 143994 153892 144000 153904
rect 144052 153892 144058 153944
rect 145650 153892 145656 153944
rect 145708 153932 145714 153944
rect 216858 153932 216864 153944
rect 145708 153904 216864 153932
rect 145708 153892 145714 153904
rect 216858 153892 216864 153904
rect 216916 153892 216922 153944
rect 222102 153892 222108 153944
rect 222160 153932 222166 153944
rect 266354 153932 266360 153944
rect 222160 153904 266360 153932
rect 222160 153892 222166 153904
rect 266354 153892 266360 153904
rect 266412 153892 266418 153944
rect 266446 153892 266452 153944
rect 266504 153932 266510 153944
rect 296990 153932 296996 153944
rect 266504 153904 296996 153932
rect 266504 153892 266510 153904
rect 296990 153892 296996 153904
rect 297048 153892 297054 153944
rect 300854 153892 300860 153944
rect 300912 153932 300918 153944
rect 312446 153932 312452 153944
rect 300912 153904 312452 153932
rect 300912 153892 300918 153904
rect 312446 153892 312452 153904
rect 312504 153892 312510 153944
rect 328454 153892 328460 153944
rect 328512 153932 328518 153944
rect 330662 153932 330668 153944
rect 328512 153904 330668 153932
rect 328512 153892 328518 153904
rect 330662 153892 330668 153904
rect 330720 153892 330726 153944
rect 334342 153892 334348 153944
rect 334400 153932 334406 153944
rect 339126 153932 339132 153944
rect 334400 153904 339132 153932
rect 334400 153892 334406 153904
rect 339126 153892 339132 153904
rect 339184 153892 339190 153944
rect 340230 153892 340236 153944
rect 340288 153932 340294 153944
rect 342990 153932 342996 153944
rect 340288 153904 342996 153932
rect 340288 153892 340294 153904
rect 342990 153892 342996 153904
rect 343048 153892 343054 153944
rect 377490 153892 377496 153944
rect 377548 153932 377554 153944
rect 382366 153932 382372 153944
rect 377548 153904 382372 153932
rect 377548 153892 377554 153904
rect 382366 153892 382372 153904
rect 382424 153892 382430 153944
rect 383286 153892 383292 153944
rect 383344 153932 383350 153944
rect 394234 153932 394240 153944
rect 383344 153904 394240 153932
rect 383344 153892 383350 153904
rect 394234 153892 394240 153904
rect 394292 153892 394298 153944
rect 394418 153892 394424 153944
rect 394476 153932 394482 153944
rect 410794 153932 410800 153944
rect 394476 153904 410800 153932
rect 394476 153892 394482 153904
rect 410794 153892 410800 153904
rect 410852 153892 410858 153944
rect 435358 153892 435364 153944
rect 435416 153932 435422 153944
rect 472158 153932 472164 153944
rect 435416 153904 472164 153932
rect 435416 153892 435422 153904
rect 472158 153892 472164 153904
rect 472216 153892 472222 153944
rect 499114 153892 499120 153944
rect 499172 153932 499178 153944
rect 567746 153932 567752 153944
rect 499172 153904 567752 153932
rect 499172 153892 499178 153904
rect 567746 153892 567752 153904
rect 567804 153892 567810 153944
rect 127575 153836 128492 153864
rect 128541 153867 128599 153873
rect 127575 153833 127587 153836
rect 127529 153827 127587 153833
rect 128541 153833 128553 153867
rect 128587 153864 128599 153867
rect 130013 153867 130071 153873
rect 130013 153864 130025 153867
rect 128587 153836 130025 153864
rect 128587 153833 128599 153836
rect 128541 153827 128599 153833
rect 130013 153833 130025 153836
rect 130059 153833 130071 153867
rect 130013 153827 130071 153833
rect 130102 153824 130108 153876
rect 130160 153864 130166 153876
rect 206462 153864 206468 153876
rect 130160 153836 206468 153864
rect 130160 153824 130166 153836
rect 206462 153824 206468 153836
rect 206520 153824 206526 153876
rect 208026 153824 208032 153876
rect 208084 153864 208090 153876
rect 258442 153864 258448 153876
rect 208084 153836 258448 153864
rect 208084 153824 208090 153836
rect 258442 153824 258448 153836
rect 258500 153824 258506 153876
rect 262122 153824 262128 153876
rect 262180 153864 262186 153876
rect 292574 153864 292580 153876
rect 262180 153836 292580 153864
rect 262180 153824 262186 153836
rect 292574 153824 292580 153836
rect 292632 153824 292638 153876
rect 295334 153824 295340 153876
rect 295392 153864 295398 153876
rect 307294 153864 307300 153876
rect 295392 153836 307300 153864
rect 295392 153824 295398 153836
rect 307294 153824 307300 153836
rect 307352 153824 307358 153876
rect 311158 153824 311164 153876
rect 311216 153864 311222 153876
rect 323118 153864 323124 153876
rect 311216 153836 323124 153864
rect 311216 153824 311222 153836
rect 323118 153824 323124 153836
rect 323176 153824 323182 153876
rect 373626 153824 373632 153876
rect 373684 153864 373690 153876
rect 379422 153864 379428 153876
rect 373684 153836 379428 153864
rect 373684 153824 373690 153836
rect 379422 153824 379428 153836
rect 379480 153824 379486 153876
rect 391198 153824 391204 153876
rect 391256 153864 391262 153876
rect 403986 153864 403992 153876
rect 391256 153836 403992 153864
rect 391256 153824 391262 153836
rect 403986 153824 403992 153836
rect 404044 153824 404050 153876
rect 408034 153824 408040 153876
rect 408092 153864 408098 153876
rect 431218 153864 431224 153876
rect 408092 153836 431224 153864
rect 408092 153824 408098 153836
rect 431218 153824 431224 153836
rect 431276 153824 431282 153876
rect 434622 153824 434628 153876
rect 434680 153864 434686 153876
rect 471238 153864 471244 153876
rect 434680 153836 471244 153864
rect 434680 153824 434686 153836
rect 471238 153824 471244 153836
rect 471296 153824 471302 153876
rect 479610 153824 479616 153876
rect 479668 153864 479674 153876
rect 487154 153864 487160 153876
rect 479668 153836 487160 153864
rect 479668 153824 479674 153836
rect 487154 153824 487160 153836
rect 487212 153824 487218 153876
rect 501690 153824 501696 153876
rect 501748 153864 501754 153876
rect 571242 153864 571248 153876
rect 501748 153836 571248 153864
rect 501748 153824 501754 153836
rect 571242 153824 571248 153836
rect 571300 153824 571306 153876
rect 78398 153756 78404 153808
rect 78456 153796 78462 153808
rect 161661 153799 161719 153805
rect 161661 153796 161673 153799
rect 78456 153768 161673 153796
rect 78456 153756 78462 153768
rect 161661 153765 161673 153768
rect 161707 153765 161719 153799
rect 172606 153796 172612 153808
rect 161661 153759 161719 153765
rect 161768 153768 172612 153796
rect 79410 153688 79416 153740
rect 79468 153728 79474 153740
rect 161768 153728 161796 153768
rect 172606 153756 172612 153768
rect 172664 153756 172670 153808
rect 179506 153756 179512 153808
rect 179564 153796 179570 153808
rect 179564 153768 185532 153796
rect 179564 153756 179570 153768
rect 79468 153700 161796 153728
rect 79468 153688 79474 153700
rect 167730 153688 167736 153740
rect 167788 153728 167794 153740
rect 169386 153728 169392 153740
rect 167788 153700 169392 153728
rect 167788 153688 167794 153700
rect 169386 153688 169392 153700
rect 169444 153688 169450 153740
rect 183002 153728 183008 153740
rect 171106 153700 183008 153728
rect 94958 153620 94964 153672
rect 95016 153660 95022 153672
rect 171106 153660 171134 153700
rect 183002 153688 183008 153700
rect 183060 153688 183066 153740
rect 95016 153632 171134 153660
rect 185504 153660 185532 153768
rect 187694 153756 187700 153808
rect 187752 153796 187758 153808
rect 216214 153796 216220 153808
rect 187752 153768 216220 153796
rect 187752 153756 187758 153768
rect 216214 153756 216220 153768
rect 216272 153756 216278 153808
rect 216582 153756 216588 153808
rect 216640 153796 216646 153808
rect 263686 153796 263692 153808
rect 216640 153768 263692 153796
rect 216640 153756 216646 153768
rect 263686 153756 263692 153768
rect 263744 153756 263750 153808
rect 271782 153756 271788 153808
rect 271840 153796 271846 153808
rect 283190 153796 283196 153808
rect 271840 153768 283196 153796
rect 271840 153756 271846 153768
rect 283190 153756 283196 153768
rect 283248 153756 283254 153808
rect 283282 153756 283288 153808
rect 283340 153796 283346 153808
rect 296162 153796 296168 153808
rect 283340 153768 296168 153796
rect 283340 153756 283346 153768
rect 296162 153756 296168 153768
rect 296220 153756 296226 153808
rect 297637 153799 297695 153805
rect 297637 153765 297649 153799
rect 297683 153796 297695 153799
rect 305270 153796 305276 153808
rect 297683 153768 305276 153796
rect 297683 153765 297695 153768
rect 297637 153759 297695 153765
rect 305270 153756 305276 153768
rect 305328 153756 305334 153808
rect 337930 153756 337936 153808
rect 337988 153796 337994 153808
rect 341058 153796 341064 153808
rect 337988 153768 341064 153796
rect 337988 153756 337994 153768
rect 341058 153756 341064 153768
rect 341116 153756 341122 153808
rect 347774 153756 347780 153808
rect 347832 153796 347838 153808
rect 351454 153796 351460 153808
rect 347832 153768 351460 153796
rect 347832 153756 347838 153768
rect 351454 153756 351460 153768
rect 351512 153756 351518 153808
rect 382734 153756 382740 153808
rect 382792 153796 382798 153808
rect 388438 153796 388444 153808
rect 382792 153768 388444 153796
rect 382792 153756 382798 153768
rect 388438 153756 388444 153768
rect 388496 153756 388502 153808
rect 395062 153756 395068 153808
rect 395120 153796 395126 153808
rect 411806 153796 411812 153808
rect 395120 153768 411812 153796
rect 395120 153756 395126 153768
rect 411806 153756 411812 153768
rect 411864 153756 411870 153808
rect 418522 153756 418528 153808
rect 418580 153796 418586 153808
rect 446858 153796 446864 153808
rect 418580 153768 446864 153796
rect 418580 153756 418586 153768
rect 446858 153756 446864 153768
rect 446916 153756 446922 153808
rect 470318 153756 470324 153808
rect 470376 153796 470382 153808
rect 524874 153796 524880 153808
rect 470376 153768 524880 153796
rect 470376 153756 470382 153768
rect 524874 153756 524880 153768
rect 524932 153756 524938 153808
rect 185578 153688 185584 153740
rect 185636 153728 185642 153740
rect 197265 153731 197323 153737
rect 197265 153728 197277 153731
rect 185636 153700 197277 153728
rect 185636 153688 185642 153700
rect 197265 153697 197277 153700
rect 197311 153697 197323 153731
rect 197265 153691 197323 153697
rect 197354 153688 197360 153740
rect 197412 153728 197418 153740
rect 222194 153728 222200 153740
rect 197412 153700 222200 153728
rect 197412 153688 197418 153700
rect 222194 153688 222200 153700
rect 222252 153688 222258 153740
rect 233234 153688 233240 153740
rect 233292 153728 233298 153740
rect 270862 153728 270868 153740
rect 233292 153700 270868 153728
rect 233292 153688 233298 153700
rect 270862 153688 270868 153700
rect 270920 153688 270926 153740
rect 271966 153688 271972 153740
rect 272024 153728 272030 153740
rect 274082 153728 274088 153740
rect 272024 153700 274088 153728
rect 272024 153688 272030 153700
rect 274082 153688 274088 153700
rect 274140 153688 274146 153740
rect 279142 153688 279148 153740
rect 279200 153728 279206 153740
rect 293586 153728 293592 153740
rect 279200 153700 293592 153728
rect 279200 153688 279206 153700
rect 293586 153688 293592 153700
rect 293644 153688 293650 153740
rect 335630 153688 335636 153740
rect 335688 153728 335694 153740
rect 339770 153728 339776 153740
rect 335688 153700 339776 153728
rect 335688 153688 335694 153700
rect 339770 153688 339776 153700
rect 339828 153688 339834 153740
rect 393038 153688 393044 153740
rect 393096 153728 393102 153740
rect 408862 153728 408868 153740
rect 393096 153700 408868 153728
rect 393096 153688 393102 153700
rect 408862 153688 408868 153700
rect 408920 153688 408926 153740
rect 413278 153688 413284 153740
rect 413336 153728 413342 153740
rect 439038 153728 439044 153740
rect 413336 153700 439044 153728
rect 413336 153688 413342 153700
rect 439038 153688 439044 153700
rect 439096 153688 439102 153740
rect 467742 153688 467748 153740
rect 467800 153728 467806 153740
rect 520918 153728 520924 153740
rect 467800 153700 520924 153728
rect 467800 153688 467806 153700
rect 520918 153688 520924 153700
rect 520976 153688 520982 153740
rect 187694 153660 187700 153672
rect 185504 153632 187700 153660
rect 95016 153620 95022 153632
rect 187694 153620 187700 153632
rect 187752 153620 187758 153672
rect 187789 153663 187847 153669
rect 187789 153629 187801 153663
rect 187835 153660 187847 153663
rect 211154 153660 211160 153672
rect 187835 153632 211160 153660
rect 187835 153629 187847 153632
rect 187789 153623 187847 153629
rect 211154 153620 211160 153632
rect 211212 153620 211218 153672
rect 237374 153620 237380 153672
rect 237432 153660 237438 153672
rect 242894 153660 242900 153672
rect 237432 153632 242900 153660
rect 237432 153620 237438 153632
rect 242894 153620 242900 153632
rect 242952 153620 242958 153672
rect 243357 153663 243415 153669
rect 243357 153629 243369 153663
rect 243403 153660 243415 153663
rect 248046 153660 248052 153672
rect 243403 153632 248052 153660
rect 243403 153629 243415 153632
rect 243357 153623 243415 153629
rect 248046 153620 248052 153632
rect 248104 153620 248110 153672
rect 249061 153663 249119 153669
rect 249061 153629 249073 153663
rect 249107 153660 249119 153663
rect 255314 153660 255320 153672
rect 249107 153632 255320 153660
rect 249107 153629 249119 153632
rect 249061 153623 249119 153629
rect 255314 153620 255320 153632
rect 255372 153620 255378 153672
rect 262214 153620 262220 153672
rect 262272 153660 262278 153672
rect 264974 153660 264980 153672
rect 262272 153632 264980 153660
rect 262272 153620 262278 153632
rect 264974 153620 264980 153632
rect 265032 153620 265038 153672
rect 272337 153663 272395 153669
rect 272337 153629 272349 153663
rect 272383 153660 272395 153663
rect 280614 153660 280620 153672
rect 272383 153632 280620 153660
rect 272383 153629 272395 153632
rect 272337 153623 272395 153629
rect 280614 153620 280620 153632
rect 280672 153620 280678 153672
rect 281534 153620 281540 153672
rect 281592 153660 281598 153672
rect 291654 153660 291660 153672
rect 281592 153632 291660 153660
rect 281592 153620 281598 153632
rect 291654 153620 291660 153632
rect 291712 153620 291718 153672
rect 292758 153620 292764 153672
rect 292816 153660 292822 153672
rect 294230 153660 294236 153672
rect 292816 153632 294236 153660
rect 292816 153620 292822 153632
rect 294230 153620 294236 153632
rect 294288 153620 294294 153672
rect 324130 153620 324136 153672
rect 324188 153660 324194 153672
rect 324866 153660 324872 153672
rect 324188 153632 324872 153660
rect 324188 153620 324194 153632
rect 324866 153620 324872 153632
rect 324924 153620 324930 153672
rect 338942 153620 338948 153672
rect 339000 153660 339006 153672
rect 342346 153660 342352 153672
rect 339000 153632 342352 153660
rect 339000 153620 339006 153632
rect 342346 153620 342352 153632
rect 342404 153620 342410 153672
rect 376478 153620 376484 153672
rect 376536 153660 376542 153672
rect 380894 153660 380900 153672
rect 376536 153632 380900 153660
rect 376536 153620 376542 153632
rect 380894 153620 380900 153632
rect 380952 153620 380958 153672
rect 389082 153620 389088 153672
rect 389140 153660 389146 153672
rect 400306 153660 400312 153672
rect 389140 153632 400312 153660
rect 389140 153620 389146 153632
rect 400306 153620 400312 153632
rect 400364 153620 400370 153672
rect 413922 153620 413928 153672
rect 413980 153660 413986 153672
rect 440050 153660 440056 153672
rect 413980 153632 440056 153660
rect 413980 153620 413986 153632
rect 440050 153620 440056 153632
rect 440108 153620 440114 153672
rect 464982 153620 464988 153672
rect 465040 153660 465046 153672
rect 517054 153660 517060 153672
rect 465040 153632 517060 153660
rect 465040 153620 465046 153632
rect 517054 153620 517060 153632
rect 517112 153620 517118 153672
rect 93026 153552 93032 153604
rect 93084 153592 93090 153604
rect 181714 153592 181720 153604
rect 93084 153564 181720 153592
rect 93084 153552 93090 153564
rect 181714 153552 181720 153564
rect 181772 153552 181778 153604
rect 182082 153552 182088 153604
rect 182140 153592 182146 153604
rect 190822 153592 190828 153604
rect 182140 153564 190828 153592
rect 182140 153552 182146 153564
rect 190822 153552 190828 153564
rect 190880 153552 190886 153604
rect 197265 153595 197323 153601
rect 197265 153561 197277 153595
rect 197311 153592 197323 153595
rect 197998 153592 198004 153604
rect 197311 153564 198004 153592
rect 197311 153561 197323 153564
rect 197265 153555 197323 153561
rect 197998 153552 198004 153564
rect 198056 153552 198062 153604
rect 248693 153595 248751 153601
rect 248693 153561 248705 153595
rect 248739 153592 248751 153595
rect 253290 153592 253296 153604
rect 248739 153564 253296 153592
rect 248739 153561 248751 153564
rect 248693 153555 248751 153561
rect 253290 153552 253296 153564
rect 253348 153552 253354 153604
rect 255866 153592 255872 153604
rect 253906 153564 255872 153592
rect 100846 153484 100852 153536
rect 100904 153524 100910 153536
rect 186958 153524 186964 153536
rect 100904 153496 186964 153524
rect 100904 153484 100910 153496
rect 186958 153484 186964 153496
rect 187016 153484 187022 153536
rect 195974 153484 195980 153536
rect 196032 153524 196038 153536
rect 211614 153524 211620 153536
rect 196032 153496 211620 153524
rect 196032 153484 196038 153496
rect 211614 153484 211620 153496
rect 211672 153484 211678 153536
rect 229186 153484 229192 153536
rect 229244 153524 229250 153536
rect 235074 153524 235080 153536
rect 229244 153496 235080 153524
rect 229244 153484 229250 153496
rect 235074 153484 235080 153496
rect 235132 153484 235138 153536
rect 251174 153484 251180 153536
rect 251232 153524 251238 153536
rect 253906 153524 253934 153564
rect 255866 153552 255872 153564
rect 255924 153552 255930 153604
rect 265066 153552 265072 153604
rect 265124 153592 265130 153604
rect 270494 153592 270500 153604
rect 265124 153564 270500 153592
rect 265124 153552 265130 153564
rect 270494 153552 270500 153564
rect 270552 153552 270558 153604
rect 280246 153552 280252 153604
rect 280304 153592 280310 153604
rect 281902 153592 281908 153604
rect 280304 153564 281908 153592
rect 280304 153552 280310 153564
rect 281902 153552 281908 153564
rect 281960 153552 281966 153604
rect 284386 153552 284392 153604
rect 284444 153592 284450 153604
rect 286410 153592 286416 153604
rect 284444 153564 286416 153592
rect 284444 153552 284450 153564
rect 286410 153552 286416 153564
rect 286468 153552 286474 153604
rect 288342 153552 288348 153604
rect 288400 153592 288406 153604
rect 297542 153592 297548 153604
rect 288400 153564 297548 153592
rect 288400 153552 288406 153564
rect 297542 153552 297548 153564
rect 297600 153552 297606 153604
rect 322934 153552 322940 153604
rect 322992 153592 322998 153604
rect 328086 153592 328092 153604
rect 322992 153564 328092 153592
rect 322992 153552 322998 153564
rect 328086 153552 328092 153564
rect 328144 153552 328150 153604
rect 380066 153552 380072 153604
rect 380124 153592 380130 153604
rect 386322 153592 386328 153604
rect 380124 153564 386328 153592
rect 380124 153552 380130 153564
rect 386322 153552 386328 153564
rect 386380 153552 386386 153604
rect 389818 153552 389824 153604
rect 389876 153592 389882 153604
rect 401686 153592 401692 153604
rect 389876 153564 401692 153592
rect 389876 153552 389882 153564
rect 401686 153552 401692 153564
rect 401744 153552 401750 153604
rect 410702 153552 410708 153604
rect 410760 153592 410766 153604
rect 435174 153592 435180 153604
rect 410760 153564 435180 153592
rect 410760 153552 410766 153564
rect 435174 153552 435180 153564
rect 435232 153552 435238 153604
rect 458082 153552 458088 153604
rect 458140 153592 458146 153604
rect 506290 153592 506296 153604
rect 458140 153564 506296 153592
rect 458140 153552 458146 153564
rect 506290 153552 506296 153564
rect 506348 153552 506354 153604
rect 251232 153496 253934 153524
rect 251232 153484 251238 153496
rect 270310 153484 270316 153536
rect 270368 153524 270374 153536
rect 272794 153524 272800 153536
rect 270368 153496 272800 153524
rect 270368 153484 270374 153496
rect 272794 153484 272800 153496
rect 272852 153484 272858 153536
rect 298002 153484 298008 153536
rect 298060 153524 298066 153536
rect 302234 153524 302240 153536
rect 298060 153496 302240 153524
rect 298060 153484 298066 153496
rect 302234 153484 302240 153496
rect 302292 153484 302298 153536
rect 317322 153484 317328 153536
rect 317380 153524 317386 153536
rect 320910 153524 320916 153536
rect 317380 153496 320916 153524
rect 317380 153484 317386 153496
rect 320910 153484 320916 153496
rect 320968 153484 320974 153536
rect 321554 153484 321560 153536
rect 321612 153524 321618 153536
rect 327442 153524 327448 153536
rect 321612 153496 327448 153524
rect 321612 153484 321618 153496
rect 327442 153484 327448 153496
rect 327500 153484 327506 153536
rect 329742 153484 329748 153536
rect 329800 153524 329806 153536
rect 331950 153524 331956 153536
rect 329800 153496 331956 153524
rect 329800 153484 329806 153496
rect 331950 153484 331956 153496
rect 332008 153484 332014 153536
rect 333974 153484 333980 153536
rect 334032 153524 334038 153536
rect 335906 153524 335912 153536
rect 334032 153496 335912 153524
rect 334032 153484 334038 153496
rect 335906 153484 335912 153496
rect 335964 153484 335970 153536
rect 338574 153484 338580 153536
rect 338632 153524 338638 153536
rect 341702 153524 341708 153536
rect 338632 153496 341708 153524
rect 338632 153484 338638 153496
rect 341702 153484 341708 153496
rect 341760 153484 341766 153536
rect 370958 153484 370964 153536
rect 371016 153524 371022 153536
rect 375742 153524 375748 153536
rect 371016 153496 375748 153524
rect 371016 153484 371022 153496
rect 375742 153484 375748 153496
rect 375800 153484 375806 153536
rect 378778 153484 378784 153536
rect 378836 153524 378842 153536
rect 384574 153524 384580 153536
rect 378836 153496 384580 153524
rect 378836 153484 378842 153496
rect 384574 153484 384580 153496
rect 384632 153484 384638 153536
rect 393774 153484 393780 153536
rect 393832 153524 393838 153536
rect 405826 153524 405832 153536
rect 393832 153496 405832 153524
rect 393832 153484 393838 153496
rect 405826 153484 405832 153496
rect 405884 153484 405890 153536
rect 477034 153484 477040 153536
rect 477092 153524 477098 153536
rect 482738 153524 482744 153536
rect 477092 153496 482744 153524
rect 477092 153484 477098 153496
rect 482738 153484 482744 153496
rect 482796 153484 482802 153536
rect 502242 153484 502248 153536
rect 502300 153524 502306 153536
rect 549162 153524 549168 153536
rect 502300 153496 549168 153524
rect 502300 153484 502306 153496
rect 549162 153484 549168 153496
rect 549220 153484 549226 153536
rect 102778 153416 102784 153468
rect 102836 153456 102842 153468
rect 188246 153456 188252 153468
rect 102836 153428 188252 153456
rect 102836 153416 102842 153428
rect 188246 153416 188252 153428
rect 188304 153416 188310 153468
rect 193122 153416 193128 153468
rect 193180 153456 193186 153468
rect 203150 153456 203156 153468
rect 193180 153428 203156 153456
rect 193180 153416 193186 153428
rect 203150 153416 203156 153428
rect 203208 153416 203214 153468
rect 242986 153416 242992 153468
rect 243044 153456 243050 153468
rect 245654 153456 245660 153468
rect 243044 153428 245660 153456
rect 243044 153416 243050 153428
rect 245654 153416 245660 153428
rect 245712 153416 245718 153468
rect 277394 153416 277400 153468
rect 277452 153456 277458 153468
rect 278774 153456 278780 153468
rect 277452 153428 278780 153456
rect 277452 153416 277458 153428
rect 278774 153416 278780 153428
rect 278832 153416 278838 153468
rect 323026 153416 323032 153468
rect 323084 153456 323090 153468
rect 327074 153456 327080 153468
rect 323084 153428 327080 153456
rect 323084 153416 323090 153428
rect 327074 153416 327080 153428
rect 327132 153416 327138 153468
rect 333882 153416 333888 153468
rect 333940 153456 333946 153468
rect 334618 153456 334624 153468
rect 333940 153428 334624 153456
rect 333940 153416 333946 153428
rect 334618 153416 334624 153428
rect 334676 153416 334682 153468
rect 365162 153416 365168 153468
rect 365220 153456 365226 153468
rect 366910 153456 366916 153468
rect 365220 153428 366916 153456
rect 365220 153416 365226 153428
rect 366910 153416 366916 153428
rect 366968 153416 366974 153468
rect 370314 153416 370320 153468
rect 370372 153456 370378 153468
rect 374730 153456 374736 153468
rect 370372 153428 374736 153456
rect 370372 153416 370378 153428
rect 374730 153416 374736 153428
rect 374788 153416 374794 153468
rect 378042 153416 378048 153468
rect 378100 153456 378106 153468
rect 382274 153456 382280 153468
rect 378100 153428 382280 153456
rect 378100 153416 378106 153428
rect 382274 153416 382280 153428
rect 382332 153416 382338 153468
rect 392486 153416 392492 153468
rect 392544 153456 392550 153468
rect 404630 153456 404636 153468
rect 392544 153428 404636 153456
rect 392544 153416 392550 153428
rect 404630 153416 404636 153428
rect 404688 153416 404694 153468
rect 455230 153416 455236 153468
rect 455288 153456 455294 153468
rect 502150 153456 502156 153468
rect 455288 153428 502156 153456
rect 455288 153416 455294 153428
rect 502150 153416 502156 153428
rect 502208 153416 502214 153468
rect 109586 153348 109592 153400
rect 109644 153388 109650 153400
rect 109644 153360 113174 153388
rect 109644 153348 109650 153360
rect 112438 153280 112444 153332
rect 112496 153320 112502 153332
rect 113146 153320 113174 153360
rect 114462 153348 114468 153400
rect 114520 153388 114526 153400
rect 196066 153388 196072 153400
rect 114520 153360 196072 153388
rect 114520 153348 114526 153360
rect 196066 153348 196072 153360
rect 196124 153348 196130 153400
rect 259362 153348 259368 153400
rect 259420 153388 259426 153400
rect 260466 153388 260472 153400
rect 259420 153360 260472 153388
rect 259420 153348 259426 153360
rect 260466 153348 260472 153360
rect 260524 153348 260530 153400
rect 297910 153348 297916 153400
rect 297968 153388 297974 153400
rect 304626 153388 304632 153400
rect 297968 153360 304632 153388
rect 297968 153348 297974 153360
rect 304626 153348 304632 153360
rect 304684 153348 304690 153400
rect 307662 153348 307668 153400
rect 307720 153388 307726 153400
rect 310514 153388 310520 153400
rect 307720 153360 310520 153388
rect 307720 153348 307726 153360
rect 310514 153348 310520 153360
rect 310572 153348 310578 153400
rect 323210 153348 323216 153400
rect 323268 153388 323274 153400
rect 326154 153388 326160 153400
rect 323268 153360 326160 153388
rect 323268 153348 323274 153360
rect 326154 153348 326160 153360
rect 326212 153348 326218 153400
rect 332318 153348 332324 153400
rect 332376 153388 332382 153400
rect 333974 153388 333980 153400
rect 332376 153360 333980 153388
rect 332376 153348 332382 153360
rect 333974 153348 333980 153360
rect 334032 153348 334038 153400
rect 336550 153348 336556 153400
rect 336608 153388 336614 153400
rect 340414 153388 340420 153400
rect 336608 153360 340420 153388
rect 336608 153348 336614 153360
rect 340414 153348 340420 153360
rect 340472 153348 340478 153400
rect 342530 153348 342536 153400
rect 342588 153388 342594 153400
rect 345198 153388 345204 153400
rect 342588 153360 345204 153388
rect 342588 153348 342594 153360
rect 345198 153348 345204 153360
rect 345256 153348 345262 153400
rect 379422 153348 379428 153400
rect 379480 153388 379486 153400
rect 384758 153388 384764 153400
rect 379480 153360 384764 153388
rect 379480 153348 379486 153360
rect 384758 153348 384764 153360
rect 384816 153348 384822 153400
rect 391842 153348 391848 153400
rect 391900 153388 391906 153400
rect 404170 153388 404176 153400
rect 391900 153360 404176 153388
rect 391900 153348 391906 153360
rect 404170 153348 404176 153360
rect 404228 153348 404234 153400
rect 456242 153348 456248 153400
rect 456300 153388 456306 153400
rect 503346 153388 503352 153400
rect 456300 153360 503352 153388
rect 456300 153348 456306 153360
rect 503346 153348 503352 153360
rect 503404 153348 503410 153400
rect 192754 153320 192760 153332
rect 112496 153292 112668 153320
rect 113146 153292 192760 153320
rect 112496 153280 112502 153292
rect 12802 153212 12808 153264
rect 12860 153252 12866 153264
rect 26694 153252 26700 153264
rect 12860 153224 26700 153252
rect 12860 153212 12866 153224
rect 26694 153212 26700 153224
rect 26752 153212 26758 153264
rect 46750 153212 46756 153264
rect 46808 153252 46814 153264
rect 92198 153252 92204 153264
rect 46808 153224 92204 153252
rect 46808 153212 46814 153224
rect 92198 153212 92204 153224
rect 92256 153212 92262 153264
rect 108942 153212 108948 153264
rect 109000 153252 109006 153264
rect 112530 153252 112536 153264
rect 109000 153224 112536 153252
rect 109000 153212 109006 153224
rect 112530 153212 112536 153224
rect 112588 153212 112594 153264
rect 112640 153252 112668 153292
rect 192754 153280 192760 153292
rect 192812 153280 192818 153332
rect 245562 153280 245568 153332
rect 245620 153320 245626 153332
rect 250714 153320 250720 153332
rect 245620 153292 250720 153320
rect 245620 153280 245626 153292
rect 250714 153280 250720 153292
rect 250772 153280 250778 153332
rect 263778 153280 263784 153332
rect 263836 153320 263842 153332
rect 268194 153320 268200 153332
rect 263836 153292 268200 153320
rect 263836 153280 263842 153292
rect 268194 153280 268200 153292
rect 268252 153280 268258 153332
rect 271690 153280 271696 153332
rect 271748 153320 271754 153332
rect 277946 153320 277952 153332
rect 271748 153292 277952 153320
rect 271748 153280 271754 153292
rect 277946 153280 277952 153292
rect 278004 153280 278010 153332
rect 303798 153280 303804 153332
rect 303856 153320 303862 153332
rect 307938 153320 307944 153332
rect 303856 153292 307944 153320
rect 303856 153280 303862 153292
rect 307938 153280 307944 153292
rect 307996 153280 308002 153332
rect 314746 153280 314752 153332
rect 314804 153320 314810 153332
rect 318334 153320 318340 153332
rect 314804 153292 318340 153320
rect 314804 153280 314810 153292
rect 318334 153280 318340 153292
rect 318392 153280 318398 153332
rect 343634 153280 343640 153332
rect 343692 153320 343698 153332
rect 345658 153320 345664 153332
rect 343692 153292 345664 153320
rect 343692 153280 343698 153292
rect 345658 153280 345664 153292
rect 345716 153280 345722 153332
rect 364150 153280 364156 153332
rect 364208 153320 364214 153332
rect 365254 153320 365260 153332
rect 364208 153292 365260 153320
rect 364208 153280 364214 153292
rect 365254 153280 365260 153292
rect 365312 153280 365318 153332
rect 371602 153280 371608 153332
rect 371660 153320 371666 153332
rect 376662 153320 376668 153332
rect 371660 153292 376668 153320
rect 371660 153280 371666 153292
rect 376662 153280 376668 153292
rect 376720 153280 376726 153332
rect 387242 153280 387248 153332
rect 387300 153320 387306 153332
rect 400030 153320 400036 153332
rect 387300 153292 400036 153320
rect 387300 153280 387306 153292
rect 400030 153280 400036 153292
rect 400088 153280 400094 153332
rect 417142 153280 417148 153332
rect 417200 153320 417206 153332
rect 417970 153320 417976 153332
rect 417200 153292 417976 153320
rect 417200 153280 417206 153292
rect 417970 153280 417976 153292
rect 418028 153280 418034 153332
rect 514662 153280 514668 153332
rect 514720 153320 514726 153332
rect 520550 153320 520556 153332
rect 514720 153292 520556 153320
rect 514720 153280 514726 153292
rect 520550 153280 520556 153292
rect 520608 153280 520614 153332
rect 117774 153252 117780 153264
rect 112640 153224 117780 153252
rect 117774 153212 117780 153224
rect 117832 153212 117838 153264
rect 117958 153212 117964 153264
rect 118016 153252 118022 153264
rect 130378 153252 130384 153264
rect 118016 153224 130384 153252
rect 118016 153212 118022 153224
rect 130378 153212 130384 153224
rect 130436 153212 130442 153264
rect 130473 153255 130531 153261
rect 130473 153221 130485 153255
rect 130519 153252 130531 153255
rect 132954 153252 132960 153264
rect 130519 153224 132960 153252
rect 130519 153221 130531 153224
rect 130473 153215 130531 153221
rect 132954 153212 132960 153224
rect 133012 153212 133018 153264
rect 133782 153212 133788 153264
rect 133840 153252 133846 153264
rect 138106 153252 138112 153264
rect 133840 153224 138112 153252
rect 133840 153212 133846 153224
rect 138106 153212 138112 153224
rect 138164 153212 138170 153264
rect 138201 153255 138259 153261
rect 138201 153221 138213 153255
rect 138247 153252 138259 153255
rect 184290 153252 184296 153264
rect 138247 153224 184296 153252
rect 138247 153221 138259 153224
rect 138201 153215 138259 153221
rect 184290 153212 184296 153224
rect 184348 153212 184354 153264
rect 189074 153212 189080 153264
rect 189132 153252 189138 153264
rect 203886 153252 203892 153264
rect 189132 153224 203892 153252
rect 189132 153212 189138 153224
rect 203886 153212 203892 153224
rect 203944 153212 203950 153264
rect 225046 153212 225052 153264
rect 225104 153252 225110 153264
rect 229830 153252 229836 153264
rect 225104 153224 229836 153252
rect 225104 153212 225110 153224
rect 229830 153212 229836 153224
rect 229888 153212 229894 153264
rect 249794 153212 249800 153264
rect 249852 153252 249858 153264
rect 254578 153252 254584 153264
rect 249852 153224 254584 153252
rect 249852 153212 249858 153224
rect 254578 153212 254584 153224
rect 254636 153212 254642 153264
rect 256694 153212 256700 153264
rect 256752 153252 256758 153264
rect 258074 153252 258080 153264
rect 256752 153224 258080 153252
rect 256752 153212 256758 153224
rect 258074 153212 258080 153224
rect 258132 153212 258138 153264
rect 285674 153212 285680 153264
rect 285732 153252 285738 153264
rect 287238 153252 287244 153264
rect 285732 153224 287244 153252
rect 285732 153212 285738 153224
rect 287238 153212 287244 153224
rect 287296 153212 287302 153264
rect 313366 153212 313372 153264
rect 313424 153252 313430 153264
rect 316034 153252 316040 153264
rect 313424 153224 316040 153252
rect 313424 153212 313430 153224
rect 316034 153212 316040 153224
rect 316092 153212 316098 153264
rect 318702 153212 318708 153264
rect 318760 153252 318766 153264
rect 322198 153252 322204 153264
rect 318760 153224 322204 153252
rect 318760 153212 318766 153224
rect 322198 153212 322204 153224
rect 322256 153212 322262 153264
rect 324406 153212 324412 153264
rect 324464 153252 324470 153264
rect 325786 153252 325792 153264
rect 324464 153224 325792 153252
rect 324464 153212 324470 153224
rect 325786 153212 325792 153224
rect 325844 153212 325850 153264
rect 334066 153212 334072 153264
rect 334124 153252 334130 153264
rect 335446 153252 335452 153264
rect 334124 153224 335452 153252
rect 334124 153212 334130 153224
rect 335446 153212 335452 153224
rect 335504 153212 335510 153264
rect 353386 153212 353392 153264
rect 353444 153252 353450 153264
rect 354858 153252 354864 153264
rect 353444 153224 354864 153252
rect 353444 153212 353450 153224
rect 354858 153212 354864 153224
rect 354916 153212 354922 153264
rect 363874 153212 363880 153264
rect 363932 153252 363938 153264
rect 364978 153252 364984 153264
rect 363932 153224 364984 153252
rect 363932 153212 363938 153224
rect 364978 153212 364984 153224
rect 365036 153212 365042 153264
rect 380710 153212 380716 153264
rect 380768 153252 380774 153264
rect 385494 153252 385500 153264
rect 380768 153224 385500 153252
rect 380768 153212 380774 153224
rect 385494 153212 385500 153224
rect 385552 153212 385558 153264
rect 412450 153212 412456 153264
rect 412508 153252 412514 153264
rect 413830 153252 413836 153264
rect 412508 153224 413836 153252
rect 412508 153212 412514 153224
rect 413830 153212 413836 153224
rect 413888 153212 413894 153264
rect 473078 153212 473084 153264
rect 473136 153252 473142 153264
rect 476114 153252 476120 153264
rect 473136 153224 476120 153252
rect 473136 153212 473142 153224
rect 476114 153212 476120 153224
rect 476172 153212 476178 153264
rect 516042 153212 516048 153264
rect 516100 153252 516106 153264
rect 520642 153252 520648 153264
rect 516100 153224 520648 153252
rect 516100 153212 516106 153224
rect 520642 153212 520648 153224
rect 520700 153212 520706 153264
rect 72602 153144 72608 153196
rect 72660 153184 72666 153196
rect 168374 153184 168380 153196
rect 72660 153156 168380 153184
rect 72660 153144 72666 153156
rect 168374 153144 168380 153156
rect 168432 153144 168438 153196
rect 170030 153144 170036 153196
rect 170088 153184 170094 153196
rect 233234 153184 233240 153196
rect 170088 153156 233240 153184
rect 170088 153144 170094 153156
rect 233234 153144 233240 153156
rect 233292 153144 233298 153196
rect 468570 153144 468576 153196
rect 468628 153184 468634 153196
rect 521930 153184 521936 153196
rect 468628 153156 521936 153184
rect 468628 153144 468634 153156
rect 521930 153144 521936 153156
rect 521988 153144 521994 153196
rect 60826 153076 60832 153128
rect 60884 153116 60890 153128
rect 160278 153116 160284 153128
rect 60884 153088 160284 153116
rect 60884 153076 60890 153088
rect 160278 153076 160284 153088
rect 160336 153076 160342 153128
rect 162302 153076 162308 153128
rect 162360 153116 162366 153128
rect 162360 153088 166672 153116
rect 162360 153076 162366 153088
rect 54018 153008 54024 153060
rect 54076 153048 54082 153060
rect 155954 153048 155960 153060
rect 54076 153020 155960 153048
rect 54076 153008 54082 153020
rect 155954 153008 155960 153020
rect 156012 153008 156018 153060
rect 156414 153008 156420 153060
rect 156472 153048 156478 153060
rect 166644 153048 166672 153088
rect 168098 153076 168104 153128
rect 168156 153116 168162 153128
rect 231854 153116 231860 153128
rect 168156 153088 231860 153116
rect 168156 153076 168162 153088
rect 231854 153076 231860 153088
rect 231912 153076 231918 153128
rect 431494 153076 431500 153128
rect 431552 153116 431558 153128
rect 466362 153116 466368 153128
rect 431552 153088 466368 153116
rect 431552 153076 431558 153088
rect 466362 153076 466368 153088
rect 466420 153076 466426 153128
rect 472434 153076 472440 153128
rect 472492 153116 472498 153128
rect 527726 153116 527732 153128
rect 472492 153088 527732 153116
rect 472492 153076 472498 153088
rect 527726 153076 527732 153088
rect 527784 153076 527790 153128
rect 227898 153048 227904 153060
rect 156472 153020 166304 153048
rect 166644 153020 227904 153048
rect 156472 153008 156478 153020
rect 49142 152940 49148 152992
rect 49200 152980 49206 152992
rect 152458 152980 152464 152992
rect 49200 152952 152464 152980
rect 49200 152940 49206 152952
rect 152458 152940 152464 152952
rect 152516 152940 152522 152992
rect 24854 152872 24860 152924
rect 24912 152912 24918 152924
rect 128998 152912 129004 152924
rect 24912 152884 129004 152912
rect 24912 152872 24918 152884
rect 128998 152872 129004 152884
rect 129056 152872 129062 152924
rect 142706 152872 142712 152924
rect 142764 152912 142770 152924
rect 149057 152915 149115 152921
rect 149057 152912 149069 152915
rect 142764 152884 149069 152912
rect 142764 152872 142770 152884
rect 149057 152881 149069 152884
rect 149103 152881 149115 152915
rect 149057 152875 149115 152881
rect 149146 152872 149152 152924
rect 149204 152912 149210 152924
rect 166077 152915 166135 152921
rect 166077 152912 166089 152915
rect 149204 152884 166089 152912
rect 149204 152872 149210 152884
rect 166077 152881 166089 152884
rect 166123 152881 166135 152915
rect 166276 152912 166304 153020
rect 227898 153008 227904 153020
rect 227956 153008 227962 153060
rect 259730 153008 259736 153060
rect 259788 153048 259794 153060
rect 292942 153048 292948 153060
rect 259788 153020 292948 153048
rect 259788 153008 259794 153020
rect 292942 153008 292948 153020
rect 293000 153008 293006 153060
rect 434070 153008 434076 153060
rect 434128 153048 434134 153060
rect 470226 153048 470232 153060
rect 434128 153020 470232 153048
rect 434128 153008 434134 153020
rect 470226 153008 470232 153020
rect 470284 153008 470290 153060
rect 476022 153008 476028 153060
rect 476080 153048 476086 153060
rect 533614 153048 533620 153060
rect 476080 153020 533620 153048
rect 476080 153008 476086 153020
rect 533614 153008 533620 153020
rect 533672 153008 533678 153060
rect 166353 152983 166411 152989
rect 166353 152949 166365 152983
rect 166399 152980 166411 152983
rect 215570 152980 215576 152992
rect 166399 152952 215576 152980
rect 166399 152949 166411 152952
rect 166353 152943 166411 152949
rect 215570 152940 215576 152952
rect 215628 152940 215634 152992
rect 255774 152940 255780 152992
rect 255832 152980 255838 152992
rect 290366 152980 290372 152992
rect 255832 152952 290372 152980
rect 255832 152940 255838 152952
rect 290366 152940 290372 152952
rect 290424 152940 290430 152992
rect 439958 152940 439964 152992
rect 440016 152980 440022 152992
rect 479058 152980 479064 152992
rect 440016 152952 479064 152980
rect 440016 152940 440022 152952
rect 479058 152940 479064 152952
rect 479116 152940 479122 152992
rect 480070 152940 480076 152992
rect 480128 152980 480134 152992
rect 539502 152980 539508 152992
rect 480128 152952 539508 152980
rect 480128 152940 480134 152952
rect 539502 152940 539508 152952
rect 539560 152940 539566 152992
rect 224034 152912 224040 152924
rect 166276 152884 224040 152912
rect 166077 152875 166135 152881
rect 224034 152872 224040 152884
rect 224092 152872 224098 152924
rect 248138 152872 248144 152924
rect 248196 152912 248202 152924
rect 285122 152912 285128 152924
rect 248196 152884 285128 152912
rect 248196 152872 248202 152884
rect 285122 152872 285128 152884
rect 285180 152872 285186 152924
rect 441706 152872 441712 152924
rect 441764 152912 441770 152924
rect 481910 152912 481916 152924
rect 441764 152884 481916 152912
rect 441764 152872 441770 152884
rect 481910 152872 481916 152884
rect 481968 152872 481974 152924
rect 484210 152872 484216 152924
rect 484268 152912 484274 152924
rect 545298 152912 545304 152924
rect 484268 152884 545304 152912
rect 484268 152872 484274 152884
rect 545298 152872 545304 152884
rect 545356 152872 545362 152924
rect 45278 152804 45284 152856
rect 45336 152844 45342 152856
rect 149882 152844 149888 152856
rect 45336 152816 149888 152844
rect 45336 152804 45342 152816
rect 149882 152804 149888 152816
rect 149940 152804 149946 152856
rect 154482 152804 154488 152856
rect 154540 152844 154546 152856
rect 222746 152844 222752 152856
rect 154540 152816 222752 152844
rect 154540 152804 154546 152816
rect 222746 152804 222752 152816
rect 222804 152804 222810 152856
rect 240318 152804 240324 152856
rect 240376 152844 240382 152856
rect 280154 152844 280160 152856
rect 240376 152816 280160 152844
rect 240376 152804 240382 152816
rect 280154 152804 280160 152816
rect 280212 152804 280218 152856
rect 444282 152804 444288 152856
rect 444340 152844 444346 152856
rect 485866 152844 485872 152856
rect 444340 152816 485872 152844
rect 444340 152804 444346 152816
rect 485866 152804 485872 152816
rect 485924 152804 485930 152856
rect 488074 152804 488080 152856
rect 488132 152844 488138 152856
rect 551186 152844 551192 152856
rect 488132 152816 551192 152844
rect 488132 152804 488138 152816
rect 551186 152804 551192 152816
rect 551244 152804 551250 152856
rect 46198 152736 46204 152788
rect 46256 152776 46262 152788
rect 150526 152776 150532 152788
rect 46256 152748 150532 152776
rect 46256 152736 46262 152748
rect 150526 152736 150532 152748
rect 150584 152736 150590 152788
rect 151538 152736 151544 152788
rect 151596 152776 151602 152788
rect 220814 152776 220820 152788
rect 151596 152748 220820 152776
rect 151596 152736 151602 152748
rect 220814 152736 220820 152748
rect 220872 152736 220878 152788
rect 232406 152736 232412 152788
rect 232464 152776 232470 152788
rect 274726 152776 274732 152788
rect 232464 152748 274732 152776
rect 232464 152736 232470 152748
rect 274726 152736 274732 152748
rect 274784 152736 274790 152788
rect 447042 152736 447048 152788
rect 447100 152776 447106 152788
rect 489270 152776 489276 152788
rect 447100 152748 489276 152776
rect 447100 152736 447106 152748
rect 489270 152736 489276 152748
rect 489328 152736 489334 152788
rect 489362 152736 489368 152788
rect 489420 152776 489426 152788
rect 553118 152776 553124 152788
rect 489420 152748 553124 152776
rect 489420 152736 489426 152748
rect 553118 152736 553124 152748
rect 553176 152736 553182 152788
rect 41322 152668 41328 152720
rect 41380 152708 41386 152720
rect 147214 152708 147220 152720
rect 41380 152680 147220 152708
rect 41380 152668 41386 152680
rect 147214 152668 147220 152680
rect 147272 152668 147278 152720
rect 217502 152708 217508 152720
rect 149256 152680 217508 152708
rect 31662 152600 31668 152652
rect 31720 152640 31726 152652
rect 139486 152640 139492 152652
rect 31720 152612 139492 152640
rect 31720 152600 31726 152612
rect 139486 152600 139492 152612
rect 139544 152600 139550 152652
rect 146662 152600 146668 152652
rect 146720 152640 146726 152652
rect 149256 152640 149284 152680
rect 217502 152668 217508 152680
rect 217560 152668 217566 152720
rect 224586 152668 224592 152720
rect 224644 152708 224650 152720
rect 269574 152708 269580 152720
rect 224644 152680 269580 152708
rect 224644 152668 224650 152680
rect 269574 152668 269580 152680
rect 269632 152668 269638 152720
rect 448422 152668 448428 152720
rect 448480 152708 448486 152720
rect 491662 152708 491668 152720
rect 448480 152680 491668 152708
rect 448480 152668 448486 152680
rect 491662 152668 491668 152680
rect 491720 152668 491726 152720
rect 491938 152668 491944 152720
rect 491996 152708 492002 152720
rect 556982 152708 556988 152720
rect 491996 152680 556988 152708
rect 491996 152668 492002 152680
rect 556982 152668 556988 152680
rect 557040 152668 557046 152720
rect 146720 152612 149284 152640
rect 149333 152643 149391 152649
rect 146720 152600 146726 152612
rect 149333 152609 149345 152643
rect 149379 152640 149391 152643
rect 214926 152640 214932 152652
rect 149379 152612 214932 152640
rect 149379 152609 149391 152612
rect 149333 152603 149391 152609
rect 214926 152600 214932 152612
rect 214984 152600 214990 152652
rect 220722 152600 220728 152652
rect 220780 152640 220786 152652
rect 266906 152640 266912 152652
rect 220780 152612 266912 152640
rect 220780 152600 220786 152612
rect 266906 152600 266912 152612
rect 266964 152600 266970 152652
rect 451642 152600 451648 152652
rect 451700 152640 451706 152652
rect 451700 152612 495756 152640
rect 451700 152600 451706 152612
rect 21910 152532 21916 152584
rect 21968 152572 21974 152584
rect 134242 152572 134248 152584
rect 21968 152544 134248 152572
rect 21968 152532 21974 152544
rect 134242 152532 134248 152544
rect 134300 152532 134306 152584
rect 138934 152532 138940 152584
rect 138992 152572 138998 152584
rect 212534 152572 212540 152584
rect 138992 152544 212540 152572
rect 138992 152532 138998 152544
rect 212534 152532 212540 152544
rect 212592 152532 212598 152584
rect 216950 152532 216956 152584
rect 217008 152572 217014 152584
rect 264330 152572 264336 152584
rect 217008 152544 264336 152572
rect 217008 152532 217014 152544
rect 264330 152532 264336 152544
rect 264388 152532 264394 152584
rect 450906 152532 450912 152584
rect 450964 152572 450970 152584
rect 495618 152572 495624 152584
rect 450964 152544 495624 152572
rect 450964 152532 450970 152544
rect 495618 152532 495624 152544
rect 495676 152532 495682 152584
rect 495728 152572 495756 152612
rect 495894 152600 495900 152652
rect 495952 152640 495958 152652
rect 562870 152640 562876 152652
rect 495952 152612 562876 152640
rect 495952 152600 495958 152612
rect 562870 152600 562876 152612
rect 562928 152600 562934 152652
rect 496446 152572 496452 152584
rect 495728 152544 496452 152572
rect 496446 152532 496452 152544
rect 496504 152532 496510 152584
rect 498102 152532 498108 152584
rect 498160 152572 498166 152584
rect 566734 152572 566740 152584
rect 498160 152544 566740 152572
rect 498160 152532 498166 152544
rect 566734 152532 566740 152544
rect 566792 152532 566798 152584
rect 7282 152464 7288 152516
rect 7340 152504 7346 152516
rect 124490 152504 124496 152516
rect 7340 152476 124496 152504
rect 7340 152464 7346 152476
rect 124490 152464 124496 152476
rect 124548 152464 124554 152516
rect 135898 152464 135904 152516
rect 135956 152504 135962 152516
rect 210326 152504 210332 152516
rect 135956 152476 210332 152504
rect 135956 152464 135962 152476
rect 210326 152464 210332 152476
rect 210384 152464 210390 152516
rect 214834 152464 214840 152516
rect 214892 152504 214898 152516
rect 263042 152504 263048 152516
rect 214892 152476 263048 152504
rect 214892 152464 214898 152476
rect 263042 152464 263048 152476
rect 263100 152464 263106 152516
rect 271414 152464 271420 152516
rect 271472 152504 271478 152516
rect 300854 152504 300860 152516
rect 271472 152476 300860 152504
rect 271472 152464 271478 152476
rect 300854 152464 300860 152476
rect 300912 152464 300918 152516
rect 423582 152464 423588 152516
rect 423640 152504 423646 152516
rect 454678 152504 454684 152516
rect 423640 152476 454684 152504
rect 423640 152464 423646 152476
rect 454678 152464 454684 152476
rect 454736 152464 454742 152516
rect 458818 152464 458824 152516
rect 458876 152504 458882 152516
rect 507302 152504 507308 152516
rect 458876 152476 507308 152504
rect 458876 152464 458882 152476
rect 507302 152464 507308 152476
rect 507360 152464 507366 152516
rect 510154 152464 510160 152516
rect 510212 152504 510218 152516
rect 578421 152507 578479 152513
rect 578421 152504 578433 152507
rect 510212 152476 578433 152504
rect 510212 152464 510218 152476
rect 578421 152473 578433 152476
rect 578467 152473 578479 152507
rect 578421 152467 578479 152473
rect 61838 152396 61844 152448
rect 61896 152436 61902 152448
rect 160922 152436 160928 152448
rect 61896 152408 160928 152436
rect 61896 152396 61902 152408
rect 160922 152396 160928 152408
rect 160980 152396 160986 152448
rect 165522 152396 165528 152448
rect 165580 152436 165586 152448
rect 228542 152436 228548 152448
rect 165580 152408 228548 152436
rect 165580 152396 165586 152408
rect 228542 152396 228548 152408
rect 228600 152396 228606 152448
rect 439314 152396 439320 152448
rect 439372 152436 439378 152448
rect 478046 152436 478052 152448
rect 439372 152408 478052 152436
rect 439372 152396 439378 152408
rect 478046 152396 478052 152408
rect 478104 152396 478110 152448
rect 482738 152396 482744 152448
rect 482796 152436 482802 152448
rect 534626 152436 534632 152448
rect 482796 152408 534632 152436
rect 482796 152396 482802 152408
rect 534626 152396 534632 152408
rect 534684 152396 534690 152448
rect 69658 152328 69664 152380
rect 69716 152368 69722 152380
rect 166074 152368 166080 152380
rect 69716 152340 166080 152368
rect 69716 152328 69722 152340
rect 166074 152328 166080 152340
rect 166132 152328 166138 152380
rect 172514 152328 172520 152380
rect 172572 152368 172578 152380
rect 233786 152368 233792 152380
rect 172572 152340 233792 152368
rect 172572 152328 172578 152340
rect 233786 152328 233792 152340
rect 233844 152328 233850 152380
rect 476114 152328 476120 152380
rect 476172 152368 476178 152380
rect 528738 152368 528744 152380
rect 476172 152340 528744 152368
rect 476172 152328 476178 152340
rect 528738 152328 528744 152340
rect 528796 152328 528802 152380
rect 77478 152260 77484 152312
rect 77536 152300 77542 152312
rect 171410 152300 171416 152312
rect 77536 152272 171416 152300
rect 77536 152260 77542 152272
rect 171410 152260 171416 152272
rect 171468 152260 171474 152312
rect 181806 152260 181812 152312
rect 181864 152300 181870 152312
rect 240962 152300 240968 152312
rect 181864 152272 240968 152300
rect 181864 152260 181870 152272
rect 240962 152260 240968 152272
rect 241020 152260 241026 152312
rect 462682 152260 462688 152312
rect 462740 152300 462746 152312
rect 513098 152300 513104 152312
rect 462740 152272 513104 152300
rect 462740 152260 462746 152272
rect 513098 152260 513104 152272
rect 513156 152260 513162 152312
rect 80330 152192 80336 152244
rect 80388 152232 80394 152244
rect 173572 152232 173578 152244
rect 80388 152204 173578 152232
rect 80388 152192 80394 152204
rect 173572 152192 173578 152204
rect 173630 152192 173636 152244
rect 185762 152192 185768 152244
rect 185820 152232 185826 152244
rect 243860 152232 243866 152244
rect 185820 152204 243866 152232
rect 185820 152192 185826 152204
rect 243860 152192 243866 152204
rect 243918 152192 243924 152244
rect 453896 152192 453902 152244
rect 453954 152232 453960 152244
rect 500494 152232 500500 152244
rect 453954 152204 500500 152232
rect 453954 152192 453960 152204
rect 500494 152192 500500 152204
rect 500552 152192 500558 152244
rect 85206 152124 85212 152176
rect 85264 152164 85270 152176
rect 176884 152164 176890 152176
rect 85264 152136 176890 152164
rect 85264 152124 85270 152136
rect 176884 152124 176890 152136
rect 176942 152124 176948 152176
rect 187602 152124 187608 152176
rect 187660 152164 187666 152176
rect 245148 152164 245154 152176
rect 187660 152136 245154 152164
rect 187660 152124 187666 152136
rect 245148 152124 245154 152136
rect 245206 152124 245212 152176
rect 452608 152124 452614 152176
rect 452666 152164 452672 152176
rect 498562 152164 498568 152176
rect 452666 152136 498568 152164
rect 452666 152124 452672 152136
rect 498562 152124 498568 152136
rect 498620 152124 498626 152176
rect 88150 152056 88156 152108
rect 88208 152096 88214 152108
rect 178816 152096 178822 152108
rect 88208 152068 178822 152096
rect 88208 152056 88214 152068
rect 178816 152056 178822 152068
rect 178874 152056 178880 152108
rect 187786 152056 187792 152108
rect 187844 152096 187850 152108
rect 191101 152099 191159 152105
rect 187844 152068 191052 152096
rect 187844 152056 187850 152068
rect 95970 151988 95976 152040
rect 96028 152028 96034 152040
rect 183646 152028 183652 152040
rect 96028 152000 183652 152028
rect 96028 151988 96034 152000
rect 183646 151988 183652 152000
rect 183704 151988 183710 152040
rect 43806 151960 43812 151972
rect 43767 151932 43812 151960
rect 43806 151920 43812 151932
rect 43864 151920 43870 151972
rect 57514 151960 57520 151972
rect 57475 151932 57520 151960
rect 57514 151920 57520 151932
rect 57572 151920 57578 151972
rect 60826 151960 60832 151972
rect 60787 151932 60832 151960
rect 60826 151920 60832 151932
rect 60884 151920 60890 151972
rect 64414 151960 64420 151972
rect 64375 151932 64420 151960
rect 64414 151920 64420 151932
rect 64472 151920 64478 151972
rect 67358 151960 67364 151972
rect 67319 151932 67364 151960
rect 67358 151920 67364 151932
rect 67416 151920 67422 151972
rect 74534 151960 74540 151972
rect 74495 151932 74540 151960
rect 74534 151920 74540 151932
rect 74592 151920 74598 151972
rect 78122 151960 78128 151972
rect 78083 151932 78128 151960
rect 78122 151920 78128 151932
rect 78180 151920 78186 151972
rect 85022 151960 85028 151972
rect 84983 151932 85028 151960
rect 85022 151920 85028 151932
rect 85080 151920 85086 151972
rect 91002 151960 91008 151972
rect 90963 151932 91008 151960
rect 91002 151920 91008 151932
rect 91060 151920 91066 151972
rect 95142 151960 95148 151972
rect 95103 151932 95148 151960
rect 95142 151920 95148 151932
rect 95200 151920 95206 151972
rect 105630 151960 105636 151972
rect 105591 151932 105636 151960
rect 105630 151920 105636 151932
rect 105688 151920 105694 151972
rect 115474 151920 115480 151972
rect 115532 151960 115538 151972
rect 190917 151963 190975 151969
rect 190917 151960 190929 151963
rect 115532 151932 190929 151960
rect 115532 151920 115538 151932
rect 190917 151929 190929 151932
rect 190963 151929 190975 151963
rect 191024 151960 191052 152068
rect 191101 152065 191113 152099
rect 191147 152096 191159 152099
rect 197032 152096 197038 152108
rect 191147 152068 197038 152096
rect 191147 152065 191159 152068
rect 191101 152059 191159 152065
rect 197032 152056 197038 152068
rect 197090 152056 197096 152108
rect 201218 152056 201224 152108
rect 201276 152096 201282 152108
rect 254256 152096 254262 152108
rect 201276 152068 254262 152096
rect 201276 152056 201282 152068
rect 254256 152056 254262 152068
rect 254314 152056 254320 152108
rect 449388 152056 449394 152108
rect 449446 152096 449452 152108
rect 493686 152096 493692 152108
rect 449446 152068 493692 152096
rect 449446 152056 449452 152068
rect 493686 152056 493692 152068
rect 493744 152056 493750 152108
rect 200114 152028 200120 152040
rect 192128 152000 200120 152028
rect 192021 151963 192079 151969
rect 192021 151960 192033 151963
rect 191024 151932 192033 151960
rect 190917 151923 190975 151929
rect 192021 151929 192033 151932
rect 192067 151929 192079 151963
rect 192021 151923 192079 151929
rect 3234 151852 3240 151904
rect 3292 151892 3298 151904
rect 115106 151892 115112 151904
rect 3292 151864 115112 151892
rect 3292 151852 3298 151864
rect 115106 151852 115112 151864
rect 115164 151852 115170 151904
rect 120442 151852 120448 151904
rect 120500 151892 120506 151904
rect 192128 151892 192156 152000
rect 200114 151988 200120 152000
rect 200172 151988 200178 152040
rect 205082 151988 205088 152040
rect 205140 152028 205146 152040
rect 256694 152028 256700 152040
rect 205140 152000 256700 152028
rect 205140 151988 205146 152000
rect 256694 151988 256700 152000
rect 256752 151988 256758 152040
rect 443822 151988 443828 152040
rect 443880 152028 443886 152040
rect 484946 152028 484952 152040
rect 443880 152000 484952 152028
rect 443880 151988 443886 152000
rect 484946 151988 484952 152000
rect 485004 151988 485010 152040
rect 238938 151960 238944 151972
rect 195348 151932 238944 151960
rect 120500 151864 192156 151892
rect 192205 151895 192263 151901
rect 120500 151852 120506 151864
rect 192205 151861 192217 151895
rect 192251 151892 192263 151895
rect 195348 151892 195376 151932
rect 238938 151920 238944 151932
rect 238996 151920 239002 151972
rect 192251 151864 195376 151892
rect 192251 151861 192263 151864
rect 192205 151855 192263 151861
rect 196526 151852 196532 151904
rect 196584 151892 196590 151904
rect 246942 151892 246948 151904
rect 196584 151864 246948 151892
rect 196584 151852 196590 151864
rect 246942 151852 246948 151864
rect 247000 151852 247006 151904
rect 503622 151852 503628 151904
rect 503680 151892 503686 151904
rect 520274 151892 520280 151904
rect 503680 151864 520280 151892
rect 503680 151852 503686 151864
rect 520274 151852 520280 151864
rect 520332 151852 520338 151904
rect 3510 151784 3516 151836
rect 3568 151824 3574 151836
rect 117038 151824 117044 151836
rect 3568 151796 117044 151824
rect 3568 151784 3574 151796
rect 117038 151784 117044 151796
rect 117096 151784 117102 151836
rect 127526 151784 127532 151836
rect 127584 151824 127590 151836
rect 204530 151824 204536 151836
rect 127584 151796 204536 151824
rect 127584 151784 127590 151796
rect 204530 151784 204536 151796
rect 204588 151784 204594 151836
rect 211062 151784 211068 151836
rect 211120 151824 211126 151836
rect 252002 151824 252008 151836
rect 211120 151796 252008 151824
rect 211120 151784 211126 151796
rect 252002 151784 252008 151796
rect 252060 151784 252066 151836
rect 505002 151784 505008 151836
rect 505060 151824 505066 151836
rect 525058 151824 525064 151836
rect 505060 151796 525064 151824
rect 505060 151784 505066 151796
rect 525058 151784 525064 151796
rect 525116 151784 525122 151836
rect 2958 151716 2964 151768
rect 3016 151756 3022 151768
rect 114186 151756 114192 151768
rect 3016 151728 114192 151756
rect 3016 151716 3022 151728
rect 114186 151716 114192 151728
rect 114244 151716 114250 151768
rect 3142 151648 3148 151700
rect 3200 151688 3206 151700
rect 115658 151688 115664 151700
rect 3200 151660 115664 151688
rect 3200 151648 3206 151660
rect 115658 151648 115664 151660
rect 115716 151648 115722 151700
rect 3234 151580 3240 151632
rect 3292 151620 3298 151632
rect 112898 151620 112904 151632
rect 3292 151592 112904 151620
rect 3292 151580 3298 151592
rect 112898 151580 112904 151592
rect 112956 151580 112962 151632
rect 16298 151552 16304 151564
rect 16259 151524 16304 151552
rect 16298 151512 16304 151524
rect 16356 151512 16362 151564
rect 26694 151512 26700 151564
rect 26752 151552 26758 151564
rect 118602 151552 118608 151564
rect 26752 151524 118608 151552
rect 26752 151512 26758 151524
rect 118602 151512 118608 151524
rect 118660 151512 118666 151564
rect 507762 151552 507768 151564
rect 489886 151524 507768 151552
rect 5074 151444 5080 151496
rect 5132 151484 5138 151496
rect 112806 151484 112812 151496
rect 5132 151456 112812 151484
rect 5132 151444 5138 151456
rect 112806 151444 112812 151456
rect 112864 151444 112870 151496
rect 3786 151376 3792 151428
rect 3844 151416 3850 151428
rect 112530 151416 112536 151428
rect 3844 151388 112536 151416
rect 3844 151376 3850 151388
rect 112530 151376 112536 151388
rect 112588 151376 112594 151428
rect 177206 151416 177212 151428
rect 177167 151388 177212 151416
rect 177206 151376 177212 151388
rect 177264 151376 177270 151428
rect 3602 151308 3608 151360
rect 3660 151348 3666 151360
rect 112990 151348 112996 151360
rect 3660 151320 112996 151348
rect 3660 151308 3666 151320
rect 112990 151308 112996 151320
rect 113048 151308 113054 151360
rect 116946 151308 116952 151360
rect 117004 151348 117010 151360
rect 489886 151348 489914 151524
rect 507762 151512 507768 151524
rect 507820 151512 507826 151564
rect 505646 151444 505652 151496
rect 505704 151484 505710 151496
rect 505704 151456 513236 151484
rect 505704 151444 505710 151456
rect 506934 151416 506940 151428
rect 117004 151320 489914 151348
rect 503410 151388 506940 151416
rect 117004 151308 117010 151320
rect 91005 151283 91063 151289
rect 91005 151249 91017 151283
rect 91051 151280 91063 151283
rect 177209 151283 177267 151289
rect 177209 151280 177221 151283
rect 91051 151252 177221 151280
rect 91051 151249 91063 151252
rect 91005 151243 91063 151249
rect 177209 151249 177221 151252
rect 177255 151249 177267 151283
rect 177209 151243 177267 151249
rect 64417 151215 64475 151221
rect 64417 151181 64429 151215
rect 64463 151212 64475 151215
rect 118050 151212 118056 151224
rect 64463 151184 118056 151212
rect 64463 151181 64475 151184
rect 64417 151175 64475 151181
rect 118050 151172 118056 151184
rect 118108 151172 118114 151224
rect 119706 151172 119712 151224
rect 119764 151212 119770 151224
rect 503410 151212 503438 151388
rect 506934 151376 506940 151388
rect 506992 151376 506998 151428
rect 503714 151308 503720 151360
rect 503772 151308 503778 151360
rect 510154 151348 510160 151360
rect 509206 151320 510160 151348
rect 119764 151184 503438 151212
rect 119764 151172 119770 151184
rect 113910 151104 113916 151156
rect 113968 151144 113974 151156
rect 503732 151144 503760 151308
rect 113968 151116 503760 151144
rect 113968 151104 113974 151116
rect 60829 151079 60887 151085
rect 60829 151045 60841 151079
rect 60875 151076 60887 151079
rect 114278 151076 114284 151088
rect 60875 151048 114284 151076
rect 60875 151045 60887 151048
rect 60829 151039 60887 151045
rect 114278 151036 114284 151048
rect 114336 151036 114342 151088
rect 119430 151036 119436 151088
rect 119488 151076 119494 151088
rect 509206 151076 509234 151320
rect 510154 151308 510160 151320
rect 510212 151308 510218 151360
rect 513208 151348 513236 151456
rect 513282 151444 513288 151496
rect 513340 151484 513346 151496
rect 520734 151484 520740 151496
rect 513340 151456 520740 151484
rect 513340 151444 513346 151456
rect 520734 151444 520740 151456
rect 520792 151444 520798 151496
rect 517974 151376 517980 151428
rect 518032 151416 518038 151428
rect 520366 151416 520372 151428
rect 518032 151388 520372 151416
rect 518032 151376 518038 151388
rect 520366 151376 520372 151388
rect 520424 151376 520430 151428
rect 513208 151320 518894 151348
rect 518866 151144 518894 151320
rect 519262 151308 519268 151360
rect 519320 151348 519326 151360
rect 520458 151348 520464 151360
rect 519320 151320 520464 151348
rect 519320 151308 519326 151320
rect 520458 151308 520464 151320
rect 520516 151308 520522 151360
rect 527818 151144 527824 151156
rect 518866 151116 527824 151144
rect 527818 151104 527824 151116
rect 527876 151104 527882 151156
rect 119488 151048 509234 151076
rect 119488 151036 119494 151048
rect 57517 151011 57575 151017
rect 57517 150977 57529 151011
rect 57563 151008 57575 151011
rect 117130 151008 117136 151020
rect 57563 150980 117136 151008
rect 57563 150977 57575 150980
rect 57517 150971 57575 150977
rect 117130 150968 117136 150980
rect 117188 150968 117194 151020
rect 105633 150943 105691 150949
rect 105633 150909 105645 150943
rect 105679 150940 105691 150943
rect 519722 150940 519728 150952
rect 105679 150912 519728 150940
rect 105679 150909 105691 150912
rect 105633 150903 105691 150909
rect 519722 150900 519728 150912
rect 519780 150900 519786 150952
rect 95145 150875 95203 150881
rect 95145 150841 95157 150875
rect 95191 150872 95203 150875
rect 522114 150872 522120 150884
rect 95191 150844 522120 150872
rect 95191 150841 95203 150844
rect 95145 150835 95203 150841
rect 522114 150832 522120 150844
rect 522172 150832 522178 150884
rect 85025 150807 85083 150813
rect 85025 150773 85037 150807
rect 85071 150804 85083 150807
rect 522206 150804 522212 150816
rect 85071 150776 522212 150804
rect 85071 150773 85083 150776
rect 85025 150767 85083 150773
rect 522206 150764 522212 150776
rect 522264 150764 522270 150816
rect 78125 150739 78183 150745
rect 78125 150705 78137 150739
rect 78171 150736 78183 150739
rect 520826 150736 520832 150748
rect 78171 150708 520832 150736
rect 78171 150705 78183 150708
rect 78125 150699 78183 150705
rect 520826 150696 520832 150708
rect 520884 150696 520890 150748
rect 74537 150671 74595 150677
rect 74537 150637 74549 150671
rect 74583 150668 74595 150671
rect 521930 150668 521936 150680
rect 74583 150640 521936 150668
rect 74583 150637 74595 150640
rect 74537 150631 74595 150637
rect 521930 150628 521936 150640
rect 521988 150628 521994 150680
rect 67361 150603 67419 150609
rect 67361 150569 67373 150603
rect 67407 150600 67419 150603
rect 521746 150600 521752 150612
rect 67407 150572 521752 150600
rect 67407 150569 67419 150572
rect 67361 150563 67419 150569
rect 521746 150560 521752 150572
rect 521804 150560 521810 150612
rect 43809 150535 43867 150541
rect 43809 150501 43821 150535
rect 43855 150532 43867 150535
rect 116854 150532 116860 150544
rect 43855 150504 116860 150532
rect 43855 150501 43867 150504
rect 43809 150495 43867 150501
rect 116854 150492 116860 150504
rect 116912 150492 116918 150544
rect 4062 150424 4068 150476
rect 4120 150464 4126 150476
rect 5534 150464 5540 150476
rect 4120 150436 5540 150464
rect 4120 150424 4126 150436
rect 5534 150424 5540 150436
rect 5592 150424 5598 150476
rect 16301 150467 16359 150473
rect 16301 150433 16313 150467
rect 16347 150464 16359 150467
rect 117774 150464 117780 150476
rect 16347 150436 117780 150464
rect 16347 150433 16359 150436
rect 16301 150427 16359 150433
rect 117774 150424 117780 150436
rect 117832 150424 117838 150476
rect 3694 150356 3700 150408
rect 3752 150396 3758 150408
rect 112438 150396 112444 150408
rect 3752 150368 112444 150396
rect 3752 150356 3758 150368
rect 112438 150356 112444 150368
rect 112496 150356 112502 150408
rect 3878 150288 3884 150340
rect 3936 150328 3942 150340
rect 114094 150328 114100 150340
rect 3936 150300 114100 150328
rect 3936 150288 3942 150300
rect 114094 150288 114100 150300
rect 114152 150288 114158 150340
rect 3970 150220 3976 150272
rect 4028 150260 4034 150272
rect 118418 150260 118424 150272
rect 4028 150232 118424 150260
rect 4028 150220 4034 150232
rect 118418 150220 118424 150232
rect 118476 150220 118482 150272
rect 112898 149336 112904 149388
rect 112956 149376 112962 149388
rect 114002 149376 114008 149388
rect 112956 149348 114008 149376
rect 112956 149336 112962 149348
rect 114002 149336 114008 149348
rect 114060 149336 114066 149388
rect 3418 149064 3424 149116
rect 3476 149104 3482 149116
rect 5074 149104 5080 149116
rect 3476 149076 5080 149104
rect 3476 149064 3482 149076
rect 5074 149064 5080 149076
rect 5132 149064 5138 149116
rect 115290 147636 115296 147688
rect 115348 147676 115354 147688
rect 117682 147676 117688 147688
rect 115348 147648 117688 147676
rect 115348 147636 115354 147648
rect 117682 147636 117688 147648
rect 117740 147636 117746 147688
rect 3234 146684 3240 146736
rect 3292 146724 3298 146736
rect 3418 146724 3424 146736
rect 3292 146696 3424 146724
rect 3292 146684 3298 146696
rect 3418 146684 3424 146696
rect 3476 146684 3482 146736
rect 112622 146208 112628 146260
rect 112680 146248 112686 146260
rect 117314 146248 117320 146260
rect 112680 146220 117320 146248
rect 112680 146208 112686 146220
rect 117314 146208 117320 146220
rect 117372 146208 117378 146260
rect 115382 142536 115388 142588
rect 115440 142576 115446 142588
rect 117314 142576 117320 142588
rect 115440 142548 117320 142576
rect 115440 142536 115446 142548
rect 117314 142536 117320 142548
rect 117372 142536 117378 142588
rect 115474 140768 115480 140820
rect 115532 140808 115538 140820
rect 117314 140808 117320 140820
rect 115532 140780 117320 140808
rect 115532 140768 115538 140780
rect 117314 140768 117320 140780
rect 117372 140768 117378 140820
rect 115566 137980 115572 138032
rect 115624 138020 115630 138032
rect 117682 138020 117688 138032
rect 115624 137992 117688 138020
rect 115624 137980 115630 137992
rect 117682 137980 117688 137992
rect 117740 137980 117746 138032
rect 115106 133832 115112 133884
rect 115164 133872 115170 133884
rect 117866 133872 117872 133884
rect 115164 133844 117872 133872
rect 115164 133832 115170 133844
rect 117866 133832 117872 133844
rect 117924 133832 117930 133884
rect 114278 133764 114284 133816
rect 114336 133804 114342 133816
rect 117314 133804 117320 133816
rect 114336 133776 117320 133804
rect 114336 133764 114342 133776
rect 117314 133764 117320 133776
rect 117372 133764 117378 133816
rect 116486 115948 116492 116000
rect 116544 115988 116550 116000
rect 117498 115988 117504 116000
rect 116544 115960 117504 115988
rect 116544 115948 116550 115960
rect 117498 115948 117504 115960
rect 117556 115948 117562 116000
rect 112714 113976 112720 114028
rect 112772 114016 112778 114028
rect 115842 114016 115848 114028
rect 112772 113988 115848 114016
rect 112772 113976 112778 113988
rect 115842 113976 115848 113988
rect 115900 113976 115906 114028
rect 112622 94324 112628 94376
rect 112680 94364 112686 94376
rect 115106 94364 115112 94376
rect 112680 94336 115112 94364
rect 112680 94324 112686 94336
rect 115106 94324 115112 94336
rect 115164 94324 115170 94376
rect 115750 88272 115756 88324
rect 115808 88312 115814 88324
rect 117682 88312 117688 88324
rect 115808 88284 117688 88312
rect 115808 88272 115814 88284
rect 117682 88272 117688 88284
rect 117740 88272 117746 88324
rect 115842 81812 115848 81864
rect 115900 81852 115906 81864
rect 117866 81852 117872 81864
rect 115900 81824 117872 81852
rect 115900 81812 115906 81824
rect 117866 81812 117872 81824
rect 117924 81812 117930 81864
rect 114186 81336 114192 81388
rect 114244 81376 114250 81388
rect 117314 81376 117320 81388
rect 114244 81348 117320 81376
rect 114244 81336 114250 81348
rect 117314 81336 117320 81348
rect 117372 81336 117378 81388
rect 115106 79296 115112 79348
rect 115164 79336 115170 79348
rect 117774 79336 117780 79348
rect 115164 79308 117780 79336
rect 115164 79296 115170 79308
rect 117774 79296 117780 79308
rect 117832 79296 117838 79348
rect 115658 78616 115664 78668
rect 115716 78656 115722 78668
rect 117682 78656 117688 78668
rect 115716 78628 117688 78656
rect 115716 78616 115722 78628
rect 117682 78616 117688 78628
rect 117740 78616 117746 78668
rect 112530 74536 112536 74588
rect 112588 74576 112594 74588
rect 114554 74576 114560 74588
rect 112588 74548 114560 74576
rect 112588 74536 112594 74548
rect 114554 74536 114560 74548
rect 114612 74536 114618 74588
rect 114094 71680 114100 71732
rect 114152 71720 114158 71732
rect 117314 71720 117320 71732
rect 114152 71692 117320 71720
rect 114152 71680 114158 71692
rect 117314 71680 117320 71692
rect 117372 71680 117378 71732
rect 114554 68960 114560 69012
rect 114612 69000 114618 69012
rect 117314 69000 117320 69012
rect 114612 68972 117320 69000
rect 114612 68960 114618 68972
rect 117314 68960 117320 68972
rect 117372 68960 117378 69012
rect 116394 67532 116400 67584
rect 116452 67572 116458 67584
rect 119430 67572 119436 67584
rect 116452 67544 119436 67572
rect 116452 67532 116458 67544
rect 119430 67532 119436 67544
rect 119488 67532 119494 67584
rect 112438 66172 112444 66224
rect 112496 66212 112502 66224
rect 117314 66212 117320 66224
rect 112496 66184 117320 66212
rect 112496 66172 112502 66184
rect 117314 66172 117320 66184
rect 117372 66172 117378 66224
rect 114002 61616 114008 61668
rect 114060 61656 114066 61668
rect 117314 61656 117320 61668
rect 114060 61628 117320 61656
rect 114060 61616 114066 61628
rect 117314 61616 117320 61628
rect 117372 61616 117378 61668
rect 2774 56856 2780 56908
rect 2832 56896 2838 56908
rect 4798 56896 4804 56908
rect 2832 56868 4804 56896
rect 2832 56856 2838 56868
rect 4798 56856 4804 56868
rect 4856 56856 4862 56908
rect 114002 55564 114008 55616
rect 114060 55604 114066 55616
rect 117314 55604 117320 55616
rect 114060 55576 117320 55604
rect 114060 55564 114066 55576
rect 117314 55564 117320 55576
rect 117372 55564 117378 55616
rect 115658 52436 115664 52488
rect 115716 52476 115722 52488
rect 117314 52476 117320 52488
rect 115716 52448 117320 52476
rect 115716 52436 115722 52448
rect 117314 52436 117320 52448
rect 117372 52436 117378 52488
rect 117314 48328 117320 48340
rect 115952 48300 117320 48328
rect 114094 48220 114100 48272
rect 114152 48260 114158 48272
rect 115952 48260 115980 48300
rect 117314 48288 117320 48300
rect 117372 48288 117378 48340
rect 114152 48232 115980 48260
rect 114152 48220 114158 48232
rect 115750 46112 115756 46164
rect 115808 46152 115814 46164
rect 117222 46152 117228 46164
rect 115808 46124 117228 46152
rect 115808 46112 115814 46124
rect 117222 46112 117228 46124
rect 117280 46112 117286 46164
rect 117866 44180 117872 44192
rect 114664 44152 117872 44180
rect 114186 44072 114192 44124
rect 114244 44112 114250 44124
rect 114664 44112 114692 44152
rect 117866 44140 117872 44152
rect 117924 44140 117930 44192
rect 114244 44084 114692 44112
rect 114244 44072 114250 44084
rect 117314 40100 117320 40112
rect 114572 40072 117320 40100
rect 3786 39992 3792 40044
rect 3844 40032 3850 40044
rect 4890 40032 4896 40044
rect 3844 40004 4896 40032
rect 3844 39992 3850 40004
rect 4890 39992 4896 40004
rect 4948 39992 4954 40044
rect 114278 39992 114284 40044
rect 114336 40032 114342 40044
rect 114572 40032 114600 40072
rect 117314 40060 117320 40072
rect 117372 40060 117378 40112
rect 114336 40004 114600 40032
rect 114336 39992 114342 40004
rect 112530 38632 112536 38684
rect 112588 38672 112594 38684
rect 117314 38672 117320 38684
rect 112588 38644 117320 38672
rect 112588 38632 112594 38644
rect 117314 38632 117320 38644
rect 117372 38632 117378 38684
rect 114554 37000 114560 37052
rect 114612 37040 114618 37052
rect 117222 37040 117228 37052
rect 114612 37012 117228 37040
rect 114612 37000 114618 37012
rect 117222 37000 117228 37012
rect 117280 37000 117286 37052
rect 114646 36184 114652 36236
rect 114704 36224 114710 36236
rect 117314 36224 117320 36236
rect 114704 36196 117320 36224
rect 114704 36184 114710 36196
rect 117314 36184 117320 36196
rect 117372 36184 117378 36236
rect 522574 34416 522580 34468
rect 522632 34456 522638 34468
rect 548518 34456 548524 34468
rect 522632 34428 548524 34456
rect 522632 34416 522638 34428
rect 548518 34416 548524 34428
rect 548576 34416 548582 34468
rect 113726 31764 113732 31816
rect 113784 31804 113790 31816
rect 117314 31804 117320 31816
rect 113784 31776 117320 31804
rect 113784 31764 113790 31776
rect 117314 31764 117320 31776
rect 117372 31764 117378 31816
rect 3694 30268 3700 30320
rect 3752 30308 3758 30320
rect 4982 30308 4988 30320
rect 3752 30280 4988 30308
rect 3752 30268 3758 30280
rect 4982 30268 4988 30280
rect 5040 30268 5046 30320
rect 113634 28976 113640 29028
rect 113692 29016 113698 29028
rect 117314 29016 117320 29028
rect 113692 28988 117320 29016
rect 113692 28976 113698 28988
rect 117314 28976 117320 28988
rect 117372 28976 117378 29028
rect 112622 27616 112628 27668
rect 112680 27656 112686 27668
rect 114462 27656 114468 27668
rect 112680 27628 114468 27656
rect 112680 27616 112686 27628
rect 114462 27616 114468 27628
rect 114520 27616 114526 27668
rect 113726 27480 113732 27532
rect 113784 27520 113790 27532
rect 114462 27520 114468 27532
rect 113784 27492 114468 27520
rect 113784 27480 113790 27492
rect 114462 27480 114468 27492
rect 114520 27480 114526 27532
rect 3602 24828 3608 24880
rect 3660 24868 3666 24880
rect 5074 24868 5080 24880
rect 3660 24840 5080 24868
rect 3660 24828 3666 24840
rect 5074 24828 5080 24840
rect 5132 24828 5138 24880
rect 3878 21360 3884 21412
rect 3936 21400 3942 21412
rect 5166 21400 5172 21412
rect 3936 21372 5172 21400
rect 3936 21360 3942 21372
rect 5166 21360 5172 21372
rect 5224 21360 5230 21412
rect 3326 17892 3332 17944
rect 3384 17932 3390 17944
rect 5258 17932 5264 17944
rect 3384 17904 5264 17932
rect 3384 17892 3390 17904
rect 5258 17892 5264 17904
rect 5316 17892 5322 17944
rect 115842 16872 115848 16924
rect 115900 16912 115906 16924
rect 117498 16912 117504 16924
rect 115900 16884 117504 16912
rect 115900 16872 115906 16884
rect 117498 16872 117504 16884
rect 117556 16872 117562 16924
rect 522666 15104 522672 15156
rect 522724 15144 522730 15156
rect 573358 15144 573364 15156
rect 522724 15116 573364 15144
rect 522724 15104 522730 15116
rect 573358 15104 573364 15116
rect 573416 15104 573422 15156
rect 113634 13812 113640 13864
rect 113692 13852 113698 13864
rect 117314 13852 117320 13864
rect 113692 13824 117320 13852
rect 113692 13812 113698 13824
rect 117314 13812 117320 13824
rect 117372 13812 117378 13864
rect 3234 13540 3240 13592
rect 3292 13580 3298 13592
rect 5442 13580 5448 13592
rect 3292 13552 5448 13580
rect 3292 13540 3298 13552
rect 5442 13540 5448 13552
rect 5500 13540 5506 13592
rect 521654 12928 521660 12980
rect 521712 12968 521718 12980
rect 521838 12968 521844 12980
rect 521712 12940 521844 12968
rect 521712 12928 521718 12940
rect 521838 12928 521844 12940
rect 521896 12928 521902 12980
rect 3970 12860 3976 12912
rect 4028 12900 4034 12912
rect 5350 12900 5356 12912
rect 4028 12872 5356 12900
rect 4028 12860 4034 12872
rect 5350 12860 5356 12872
rect 5408 12860 5414 12912
rect 117682 11704 117688 11756
rect 117740 11744 117746 11756
rect 117958 11744 117964 11756
rect 117740 11716 117964 11744
rect 117740 11704 117746 11716
rect 117958 11704 117964 11716
rect 118016 11704 118022 11756
rect 115106 9664 115112 9716
rect 115164 9704 115170 9716
rect 117314 9704 117320 9716
rect 115164 9676 117320 9704
rect 115164 9664 115170 9676
rect 117314 9664 117320 9676
rect 117372 9664 117378 9716
rect 3326 8916 3332 8968
rect 3384 8956 3390 8968
rect 3602 8956 3608 8968
rect 3384 8928 3608 8956
rect 3384 8916 3390 8928
rect 3602 8916 3608 8928
rect 3660 8916 3666 8968
rect 3602 8780 3608 8832
rect 3660 8820 3666 8832
rect 4062 8820 4068 8832
rect 3660 8792 4068 8820
rect 3660 8780 3666 8792
rect 4062 8780 4068 8792
rect 4120 8780 4126 8832
rect 116026 8304 116032 8356
rect 116084 8344 116090 8356
rect 118970 8344 118976 8356
rect 116084 8316 118976 8344
rect 116084 8304 116090 8316
rect 118970 8304 118976 8316
rect 119028 8304 119034 8356
rect 114554 7148 114560 7200
rect 114612 7188 114618 7200
rect 117314 7188 117320 7200
rect 114612 7160 117320 7188
rect 114612 7148 114618 7160
rect 117314 7148 117320 7160
rect 117372 7148 117378 7200
rect 112438 5924 112444 5976
rect 112496 5964 112502 5976
rect 112714 5964 112720 5976
rect 112496 5936 112720 5964
rect 112496 5924 112502 5936
rect 112714 5924 112720 5936
rect 112772 5924 112778 5976
rect 2958 5856 2964 5908
rect 3016 5896 3022 5908
rect 118510 5896 118516 5908
rect 3016 5868 118516 5896
rect 3016 5856 3022 5868
rect 118510 5856 118516 5868
rect 118568 5856 118574 5908
rect 2866 5788 2872 5840
rect 2924 5828 2930 5840
rect 117866 5828 117872 5840
rect 2924 5800 117872 5828
rect 2924 5788 2930 5800
rect 117866 5788 117872 5800
rect 117924 5788 117930 5840
rect 2774 5720 2780 5772
rect 2832 5760 2838 5772
rect 117130 5760 117136 5772
rect 2832 5732 117136 5760
rect 2832 5720 2838 5732
rect 117130 5720 117136 5732
rect 117188 5720 117194 5772
rect 3786 5652 3792 5704
rect 3844 5692 3850 5704
rect 117774 5692 117780 5704
rect 3844 5664 117780 5692
rect 3844 5652 3850 5664
rect 117774 5652 117780 5664
rect 117832 5652 117838 5704
rect 3142 5584 3148 5636
rect 3200 5624 3206 5636
rect 114462 5624 114468 5636
rect 3200 5596 114468 5624
rect 3200 5584 3206 5596
rect 114462 5584 114468 5596
rect 114520 5584 114526 5636
rect 3050 5516 3056 5568
rect 3108 5556 3114 5568
rect 113726 5556 113732 5568
rect 3108 5528 113732 5556
rect 3108 5516 3114 5528
rect 113726 5516 113732 5528
rect 113784 5516 113790 5568
rect 3970 5448 3976 5500
rect 4028 5488 4034 5500
rect 117222 5488 117228 5500
rect 4028 5460 117228 5488
rect 4028 5448 4034 5460
rect 117222 5448 117228 5460
rect 117280 5448 117286 5500
rect 3418 5380 3424 5432
rect 3476 5420 3482 5432
rect 108393 5423 108451 5429
rect 3476 5392 108344 5420
rect 3476 5380 3482 5392
rect 3694 5312 3700 5364
rect 3752 5352 3758 5364
rect 108209 5355 108267 5361
rect 108209 5352 108221 5355
rect 3752 5324 108221 5352
rect 3752 5312 3758 5324
rect 108209 5321 108221 5324
rect 108255 5321 108267 5355
rect 108316 5352 108344 5392
rect 108393 5389 108405 5423
rect 108439 5420 108451 5423
rect 112438 5420 112444 5432
rect 108439 5392 112444 5420
rect 108439 5389 108451 5392
rect 108393 5383 108451 5389
rect 112438 5380 112444 5392
rect 112496 5380 112502 5432
rect 112622 5380 112628 5432
rect 112680 5420 112686 5432
rect 115290 5420 115296 5432
rect 112680 5392 115296 5420
rect 112680 5380 112686 5392
rect 115290 5380 115296 5392
rect 115348 5380 115354 5432
rect 115658 5352 115664 5364
rect 108316 5324 115664 5352
rect 108209 5315 108267 5321
rect 115658 5312 115664 5324
rect 115716 5312 115722 5364
rect 116578 5312 116584 5364
rect 116636 5352 116642 5364
rect 116946 5352 116952 5364
rect 116636 5324 116952 5352
rect 116636 5312 116642 5324
rect 116946 5312 116952 5324
rect 117004 5312 117010 5364
rect 3234 5244 3240 5296
rect 3292 5284 3298 5296
rect 114554 5284 114560 5296
rect 3292 5256 114560 5284
rect 3292 5244 3298 5256
rect 114554 5244 114560 5256
rect 114612 5244 114618 5296
rect 4062 5176 4068 5228
rect 4120 5216 4126 5228
rect 115106 5216 115112 5228
rect 4120 5188 115112 5216
rect 4120 5176 4126 5188
rect 115106 5176 115112 5188
rect 115164 5176 115170 5228
rect 3510 5108 3516 5160
rect 3568 5148 3574 5160
rect 114370 5148 114376 5160
rect 3568 5120 114376 5148
rect 3568 5108 3574 5120
rect 114370 5108 114376 5120
rect 114428 5108 114434 5160
rect 116670 5108 116676 5160
rect 116728 5148 116734 5160
rect 168837 5151 168895 5157
rect 168837 5148 168849 5151
rect 116728 5120 168849 5148
rect 116728 5108 116734 5120
rect 168837 5117 168849 5120
rect 168883 5117 168895 5151
rect 168837 5111 168895 5117
rect 474461 5151 474519 5157
rect 474461 5117 474473 5151
rect 474507 5148 474519 5151
rect 571978 5148 571984 5160
rect 474507 5120 571984 5148
rect 474507 5117 474519 5120
rect 474461 5111 474519 5117
rect 571978 5108 571984 5120
rect 572036 5108 572042 5160
rect 4982 5040 4988 5092
rect 5040 5080 5046 5092
rect 108209 5083 108267 5089
rect 108209 5080 108221 5083
rect 5040 5052 108221 5080
rect 5040 5040 5046 5052
rect 108209 5049 108221 5052
rect 108255 5049 108267 5083
rect 108209 5043 108267 5049
rect 108301 5083 108359 5089
rect 108301 5049 108313 5083
rect 108347 5080 108359 5083
rect 114002 5080 114008 5092
rect 108347 5052 114008 5080
rect 108347 5049 108359 5052
rect 108301 5043 108359 5049
rect 114002 5040 114008 5052
rect 114060 5040 114066 5092
rect 118878 5040 118884 5092
rect 118936 5080 118942 5092
rect 518621 5083 518679 5089
rect 518621 5080 518633 5083
rect 118936 5052 518633 5080
rect 118936 5040 118942 5052
rect 518621 5049 518633 5052
rect 518667 5049 518679 5083
rect 518621 5043 518679 5049
rect 86865 5015 86923 5021
rect 86865 4981 86877 5015
rect 86911 5012 86923 5015
rect 521746 5012 521752 5024
rect 86911 4984 521752 5012
rect 86911 4981 86923 4984
rect 86865 4975 86923 4981
rect 521746 4972 521752 4984
rect 521804 4972 521810 5024
rect 3326 4904 3332 4956
rect 3384 4944 3390 4956
rect 113634 4944 113640 4956
rect 3384 4916 113640 4944
rect 3384 4904 3390 4916
rect 113634 4904 113640 4916
rect 113692 4904 113698 4956
rect 118694 4904 118700 4956
rect 118752 4944 118758 4956
rect 566550 4944 566556 4956
rect 118752 4916 566556 4944
rect 118752 4904 118758 4916
rect 566550 4904 566556 4916
rect 566608 4904 566614 4956
rect 65981 4879 66039 4885
rect 65981 4845 65993 4879
rect 66027 4876 66039 4879
rect 520826 4876 520832 4888
rect 66027 4848 520832 4876
rect 66027 4845 66039 4848
rect 65981 4839 66039 4845
rect 520826 4836 520832 4848
rect 520884 4836 520890 4888
rect 4890 4768 4896 4820
rect 4948 4808 4954 4820
rect 108301 4811 108359 4817
rect 108301 4808 108313 4811
rect 4948 4780 108313 4808
rect 4948 4768 4954 4780
rect 108301 4777 108313 4780
rect 108347 4777 108359 4811
rect 108301 4771 108359 4777
rect 108393 4811 108451 4817
rect 108393 4777 108405 4811
rect 108439 4808 108451 4811
rect 115842 4808 115848 4820
rect 108439 4780 115848 4808
rect 108439 4777 108451 4780
rect 108393 4771 108451 4777
rect 115842 4768 115848 4780
rect 115900 4768 115906 4820
rect 118786 4768 118792 4820
rect 118844 4808 118850 4820
rect 577222 4808 577228 4820
rect 118844 4780 577228 4808
rect 118844 4768 118850 4780
rect 577222 4768 577228 4780
rect 577280 4768 577286 4820
rect 5074 4700 5080 4752
rect 5132 4740 5138 4752
rect 114094 4740 114100 4752
rect 5132 4712 114100 4740
rect 5132 4700 5138 4712
rect 114094 4700 114100 4712
rect 114152 4700 114158 4752
rect 5166 4632 5172 4684
rect 5224 4672 5230 4684
rect 114186 4672 114192 4684
rect 5224 4644 114192 4672
rect 5224 4632 5230 4644
rect 114186 4632 114192 4644
rect 114244 4632 114250 4684
rect 168834 4672 168840 4684
rect 168795 4644 168840 4672
rect 168834 4632 168840 4644
rect 168892 4632 168898 4684
rect 474458 4672 474464 4684
rect 474419 4644 474464 4672
rect 474458 4632 474464 4644
rect 474516 4632 474522 4684
rect 518618 4672 518624 4684
rect 518579 4644 518624 4672
rect 518618 4632 518624 4644
rect 518676 4632 518682 4684
rect 519630 4632 519636 4684
rect 519688 4672 519694 4684
rect 522390 4672 522396 4684
rect 519688 4644 522396 4672
rect 519688 4632 519694 4644
rect 522390 4632 522396 4644
rect 522448 4632 522454 4684
rect 5350 4564 5356 4616
rect 5408 4604 5414 4616
rect 114278 4604 114284 4616
rect 5408 4576 114284 4604
rect 5408 4564 5414 4576
rect 114278 4564 114284 4576
rect 114336 4564 114342 4616
rect 5258 4496 5264 4548
rect 5316 4536 5322 4548
rect 108209 4539 108267 4545
rect 5316 4508 108068 4536
rect 5316 4496 5322 4508
rect 5442 4428 5448 4480
rect 5500 4468 5506 4480
rect 107933 4471 107991 4477
rect 107933 4468 107945 4471
rect 5500 4440 107945 4468
rect 5500 4428 5506 4440
rect 107933 4437 107945 4440
rect 107979 4437 107991 4471
rect 108040 4468 108068 4508
rect 108209 4505 108221 4539
rect 108255 4536 108267 4539
rect 115750 4536 115756 4548
rect 108255 4508 115756 4536
rect 108255 4505 108267 4508
rect 108209 4499 108267 4505
rect 115750 4496 115756 4508
rect 115808 4496 115814 4548
rect 112714 4468 112720 4480
rect 108040 4440 112720 4468
rect 107933 4431 107991 4437
rect 112714 4428 112720 4440
rect 112772 4428 112778 4480
rect 42610 4360 42616 4412
rect 42668 4400 42674 4412
rect 118326 4400 118332 4412
rect 42668 4372 118332 4400
rect 42668 4360 42674 4372
rect 118326 4360 118332 4372
rect 118384 4360 118390 4412
rect 62666 4292 62672 4344
rect 62724 4332 62730 4344
rect 116762 4332 116768 4344
rect 62724 4304 116768 4332
rect 62724 4292 62730 4304
rect 116762 4292 116768 4304
rect 116820 4292 116826 4344
rect 65978 4264 65984 4276
rect 65939 4236 65984 4264
rect 65978 4224 65984 4236
rect 66036 4224 66042 4276
rect 66162 4224 66168 4276
rect 66220 4264 66226 4276
rect 118050 4264 118056 4276
rect 66220 4236 118056 4264
rect 66220 4224 66226 4236
rect 118050 4224 118056 4236
rect 118108 4224 118114 4276
rect 2958 4156 2964 4208
rect 3016 4196 3022 4208
rect 117314 4196 117320 4208
rect 3016 4168 117320 4196
rect 3016 4156 3022 4168
rect 117314 4156 117320 4168
rect 117372 4156 117378 4208
rect 520090 4156 520096 4208
rect 520148 4196 520154 4208
rect 522114 4196 522120 4208
rect 520148 4168 522120 4196
rect 520148 4156 520154 4168
rect 522114 4156 522120 4168
rect 522172 4156 522178 4208
rect 7834 4088 7840 4140
rect 7892 4128 7898 4140
rect 124674 4128 124680 4140
rect 7892 4100 124680 4128
rect 7892 4088 7898 4100
rect 124674 4088 124680 4100
rect 124732 4088 124738 4140
rect 125134 4088 125140 4140
rect 125192 4128 125198 4140
rect 125192 4100 127756 4128
rect 125192 4088 125198 4100
rect 45094 4020 45100 4072
rect 45152 4060 45158 4072
rect 116854 4060 116860 4072
rect 45152 4032 116860 4060
rect 45152 4020 45158 4032
rect 116854 4020 116860 4032
rect 116912 4020 116918 4072
rect 117038 4020 117044 4072
rect 117096 4060 117102 4072
rect 125505 4063 125563 4069
rect 117096 4032 122834 4060
rect 117096 4020 117102 4032
rect 86862 3992 86868 4004
rect 86823 3964 86868 3992
rect 86862 3952 86868 3964
rect 86920 3952 86926 4004
rect 107933 3995 107991 4001
rect 107933 3961 107945 3995
rect 107979 3992 107991 3995
rect 114189 3995 114247 4001
rect 114189 3992 114201 3995
rect 107979 3964 114201 3992
rect 107979 3961 107991 3964
rect 107933 3955 107991 3961
rect 114189 3961 114201 3964
rect 114235 3961 114247 3995
rect 114189 3955 114247 3961
rect 114278 3952 114284 4004
rect 114336 3992 114342 4004
rect 121641 3995 121699 4001
rect 121641 3992 121653 3995
rect 114336 3964 121653 3992
rect 114336 3952 114342 3964
rect 121641 3961 121653 3964
rect 121687 3961 121699 3995
rect 122806 3992 122834 4032
rect 125505 4029 125517 4063
rect 125551 4060 125563 4063
rect 127621 4063 127679 4069
rect 127621 4060 127633 4063
rect 125551 4032 127633 4060
rect 125551 4029 125563 4032
rect 125505 4023 125563 4029
rect 127621 4029 127633 4032
rect 127667 4029 127679 4063
rect 127728 4060 127756 4100
rect 130286 4088 130292 4140
rect 130344 4128 130350 4140
rect 198734 4128 198740 4140
rect 130344 4100 198740 4128
rect 130344 4088 130350 4100
rect 198734 4088 198740 4100
rect 198792 4088 198798 4140
rect 404262 4088 404268 4140
rect 404320 4128 404326 4140
rect 454310 4128 454316 4140
rect 404320 4100 454316 4128
rect 404320 4088 404326 4100
rect 454310 4088 454316 4100
rect 454368 4088 454374 4140
rect 527818 4088 527824 4140
rect 527876 4128 527882 4140
rect 529290 4128 529296 4140
rect 527876 4100 529296 4128
rect 527876 4088 527882 4100
rect 529290 4088 529296 4100
rect 529348 4088 529354 4140
rect 195238 4060 195244 4072
rect 127728 4032 195244 4060
rect 127621 4023 127679 4029
rect 195238 4020 195244 4032
rect 195296 4020 195302 4072
rect 215386 4020 215392 4072
rect 215444 4060 215450 4072
rect 252554 4060 252560 4072
rect 215444 4032 252560 4060
rect 215444 4020 215450 4032
rect 252554 4020 252560 4032
rect 252612 4020 252618 4072
rect 407666 4020 407672 4072
rect 407724 4060 407730 4072
rect 460106 4060 460112 4072
rect 407724 4032 460112 4060
rect 407724 4020 407730 4032
rect 460106 4020 460112 4032
rect 460164 4020 460170 4072
rect 461486 4020 461492 4072
rect 461544 4060 461550 4072
rect 545298 4060 545304 4072
rect 461544 4032 545304 4060
rect 461544 4020 461550 4032
rect 545298 4020 545304 4032
rect 545356 4020 545362 4072
rect 470870 3992 470876 4004
rect 122806 3964 470876 3992
rect 121641 3955 121699 3961
rect 470870 3952 470876 3964
rect 470928 3952 470934 4004
rect 77018 3884 77024 3936
rect 77076 3924 77082 3936
rect 164970 3924 164976 3936
rect 77076 3896 164976 3924
rect 77076 3884 77082 3896
rect 164970 3884 164976 3896
rect 165028 3884 165034 3936
rect 219112 3924 219118 3936
rect 165172 3896 219118 3924
rect 82354 3816 82360 3868
rect 82412 3856 82418 3868
rect 165065 3859 165123 3865
rect 165065 3856 165077 3859
rect 82412 3828 165077 3856
rect 82412 3816 82418 3828
rect 165065 3825 165077 3828
rect 165111 3825 165123 3859
rect 165065 3819 165123 3825
rect 66438 3748 66444 3800
rect 66496 3788 66502 3800
rect 158254 3788 158260 3800
rect 66496 3760 158260 3788
rect 66496 3748 66502 3760
rect 158254 3748 158260 3760
rect 158312 3748 158318 3800
rect 162210 3748 162216 3800
rect 162268 3788 162274 3800
rect 165172 3788 165200 3896
rect 219112 3884 219118 3896
rect 219170 3884 219176 3936
rect 311158 3884 311164 3936
rect 311216 3924 311222 3936
rect 313228 3924 313234 3936
rect 311216 3896 313234 3924
rect 311216 3884 311222 3896
rect 313228 3884 313234 3896
rect 313286 3884 313292 3936
rect 414060 3884 414066 3936
rect 414118 3924 414124 3936
rect 470778 3924 470784 3936
rect 414118 3896 470784 3924
rect 414118 3884 414124 3896
rect 470778 3884 470784 3896
rect 470836 3884 470842 3936
rect 165249 3859 165307 3865
rect 165249 3825 165261 3859
rect 165295 3856 165307 3859
rect 168282 3856 168288 3868
rect 165295 3828 168288 3856
rect 165295 3825 165307 3828
rect 165249 3819 165307 3825
rect 168282 3816 168288 3828
rect 168340 3816 168346 3868
rect 178126 3816 178132 3868
rect 178184 3856 178190 3868
rect 229094 3856 229100 3868
rect 178184 3828 229100 3856
rect 178184 3816 178190 3828
rect 229094 3816 229100 3828
rect 229152 3816 229158 3868
rect 417786 3816 417792 3868
rect 417844 3856 417850 3868
rect 476114 3856 476120 3868
rect 417844 3828 476120 3856
rect 417844 3816 417850 3828
rect 476114 3816 476120 3828
rect 476172 3816 476178 3868
rect 162268 3760 165200 3788
rect 162268 3748 162274 3760
rect 167454 3748 167460 3800
rect 167512 3788 167518 3800
rect 222194 3788 222200 3800
rect 167512 3760 222200 3788
rect 167512 3748 167518 3760
rect 222194 3748 222200 3760
rect 222252 3748 222258 3800
rect 420730 3748 420736 3800
rect 420788 3788 420794 3800
rect 481450 3788 481456 3800
rect 420788 3760 481456 3788
rect 420788 3748 420794 3760
rect 481450 3748 481456 3760
rect 481508 3748 481514 3800
rect 61102 3680 61108 3732
rect 61160 3720 61166 3732
rect 154942 3720 154948 3732
rect 61160 3692 154948 3720
rect 61160 3680 61166 3692
rect 154942 3680 154948 3692
rect 155000 3680 155006 3732
rect 212074 3720 212080 3732
rect 156616 3692 212080 3720
rect 55766 3612 55772 3664
rect 55824 3652 55830 3664
rect 146938 3652 146944 3664
rect 55824 3624 146944 3652
rect 55824 3612 55830 3624
rect 146938 3612 146944 3624
rect 146996 3612 147002 3664
rect 151538 3612 151544 3664
rect 151596 3652 151602 3664
rect 156616 3652 156644 3692
rect 212074 3680 212080 3692
rect 212132 3680 212138 3732
rect 241974 3680 241980 3732
rect 242032 3720 242038 3732
rect 269206 3720 269212 3732
rect 242032 3692 269212 3720
rect 242032 3680 242038 3692
rect 269206 3680 269212 3692
rect 269264 3680 269270 3732
rect 411070 3680 411076 3732
rect 411128 3720 411134 3732
rect 465442 3720 465448 3732
rect 411128 3692 465448 3720
rect 411128 3680 411134 3692
rect 465442 3680 465448 3692
rect 465500 3680 465506 3732
rect 151596 3624 156644 3652
rect 156693 3655 156751 3661
rect 151596 3612 151602 3624
rect 156693 3621 156705 3655
rect 156739 3652 156751 3655
rect 208670 3652 208676 3664
rect 156739 3624 208676 3652
rect 156739 3621 156751 3624
rect 156693 3615 156751 3621
rect 208670 3612 208676 3624
rect 208728 3612 208734 3664
rect 226058 3612 226064 3664
rect 226116 3652 226122 3664
rect 259454 3652 259460 3664
rect 226116 3624 259460 3652
rect 226116 3612 226122 3624
rect 259454 3612 259460 3624
rect 259512 3612 259518 3664
rect 367002 3612 367008 3664
rect 367060 3652 367066 3664
rect 396258 3652 396264 3664
rect 367060 3624 396264 3652
rect 367060 3612 367066 3624
rect 396258 3612 396264 3624
rect 396316 3612 396322 3664
rect 400861 3655 400919 3661
rect 400861 3621 400873 3655
rect 400907 3652 400919 3655
rect 401594 3652 401600 3664
rect 400907 3624 401600 3652
rect 400907 3621 400919 3624
rect 400861 3615 400919 3621
rect 401594 3612 401600 3624
rect 401652 3612 401658 3664
rect 424502 3612 424508 3664
rect 424560 3652 424566 3664
rect 486694 3652 486700 3664
rect 424560 3624 486700 3652
rect 424560 3612 424566 3624
rect 486694 3612 486700 3624
rect 486752 3612 486758 3664
rect 50430 3544 50436 3596
rect 50488 3584 50494 3596
rect 141602 3584 141608 3596
rect 50488 3556 141608 3584
rect 50488 3544 50494 3556
rect 141602 3544 141608 3556
rect 141660 3544 141666 3596
rect 205634 3584 205640 3596
rect 141712 3556 205640 3584
rect 39758 3476 39764 3528
rect 39816 3516 39822 3528
rect 107933 3519 107991 3525
rect 107933 3516 107945 3519
rect 39816 3488 107945 3516
rect 39816 3476 39822 3488
rect 107933 3485 107945 3488
rect 107979 3485 107991 3519
rect 107933 3479 107991 3485
rect 108850 3476 108856 3528
rect 108908 3516 108914 3528
rect 113910 3516 113916 3528
rect 108908 3488 113916 3516
rect 108908 3476 108914 3488
rect 113910 3476 113916 3488
rect 113968 3476 113974 3528
rect 114189 3519 114247 3525
rect 114189 3485 114201 3519
rect 114235 3516 114247 3519
rect 114646 3516 114652 3528
rect 114235 3488 114652 3516
rect 114235 3485 114247 3488
rect 114189 3479 114247 3485
rect 114646 3476 114652 3488
rect 114704 3476 114710 3528
rect 114741 3519 114799 3525
rect 114741 3485 114753 3519
rect 114787 3516 114799 3519
rect 118234 3516 118240 3528
rect 114787 3488 118240 3516
rect 114787 3485 114799 3488
rect 114741 3479 114799 3485
rect 118234 3476 118240 3488
rect 118292 3476 118298 3528
rect 118970 3476 118976 3528
rect 119028 3516 119034 3528
rect 125505 3519 125563 3525
rect 125505 3516 125517 3519
rect 119028 3488 125517 3516
rect 119028 3476 119034 3488
rect 125505 3485 125517 3488
rect 125551 3485 125563 3519
rect 125505 3479 125563 3485
rect 125597 3519 125655 3525
rect 125597 3485 125609 3519
rect 125643 3516 125655 3519
rect 128354 3516 128360 3528
rect 125643 3488 128360 3516
rect 125643 3485 125655 3488
rect 125597 3479 125655 3485
rect 128354 3476 128360 3488
rect 128412 3476 128418 3528
rect 140866 3476 140872 3528
rect 140924 3516 140930 3528
rect 141712 3516 141740 3556
rect 205634 3544 205640 3556
rect 205692 3544 205698 3596
rect 373902 3544 373908 3596
rect 373960 3584 373966 3596
rect 406930 3584 406936 3596
rect 373960 3556 406936 3584
rect 373960 3544 373966 3556
rect 406930 3544 406936 3556
rect 406988 3544 406994 3596
rect 427722 3544 427728 3596
rect 427780 3584 427786 3596
rect 492030 3584 492036 3596
rect 427780 3556 492036 3584
rect 427780 3544 427786 3556
rect 492030 3544 492036 3556
rect 492088 3544 492094 3596
rect 508038 3544 508044 3596
rect 508096 3584 508102 3596
rect 520274 3584 520280 3596
rect 508096 3556 520280 3584
rect 508096 3544 508102 3556
rect 520274 3544 520280 3556
rect 520332 3544 520338 3596
rect 140924 3488 141740 3516
rect 141789 3519 141847 3525
rect 140924 3476 140930 3488
rect 141789 3485 141801 3519
rect 141835 3516 141847 3519
rect 201954 3516 201960 3528
rect 141835 3488 201960 3516
rect 141835 3485 141847 3488
rect 141789 3479 141847 3485
rect 201954 3476 201960 3488
rect 202012 3476 202018 3528
rect 213822 3476 213828 3528
rect 213880 3516 213886 3528
rect 521838 3516 521844 3528
rect 213880 3488 521844 3516
rect 213880 3476 213886 3488
rect 521838 3476 521844 3488
rect 521896 3476 521902 3528
rect 98362 3408 98368 3460
rect 98420 3448 98426 3460
rect 178494 3448 178500 3460
rect 98420 3420 178500 3448
rect 98420 3408 98426 3420
rect 178494 3408 178500 3420
rect 178552 3408 178558 3460
rect 522206 3448 522212 3460
rect 178604 3420 522212 3448
rect 93026 3340 93032 3392
rect 93084 3380 93090 3392
rect 175274 3380 175280 3392
rect 93084 3352 175280 3380
rect 93084 3340 93090 3352
rect 175274 3340 175280 3352
rect 175332 3340 175338 3392
rect 176654 3340 176660 3392
rect 176712 3380 176718 3392
rect 178604 3380 178632 3420
rect 522206 3408 522212 3420
rect 522264 3408 522270 3460
rect 525058 3408 525064 3460
rect 525116 3448 525122 3460
rect 539962 3448 539968 3460
rect 525116 3420 539968 3448
rect 525116 3408 525122 3420
rect 539962 3408 539968 3420
rect 540020 3408 540026 3460
rect 225506 3380 225512 3392
rect 176712 3352 178632 3380
rect 180766 3352 225512 3380
rect 176712 3340 176718 3352
rect 87690 3272 87696 3324
rect 87748 3312 87754 3324
rect 171778 3312 171784 3324
rect 87748 3284 171784 3312
rect 87748 3272 87754 3284
rect 171778 3272 171784 3284
rect 171836 3272 171842 3324
rect 172790 3272 172796 3324
rect 172848 3312 172854 3324
rect 180766 3312 180794 3352
rect 225506 3340 225512 3352
rect 225564 3340 225570 3392
rect 231302 3340 231308 3392
rect 231360 3380 231366 3392
rect 262490 3380 262496 3392
rect 231360 3352 262496 3380
rect 231360 3340 231366 3352
rect 262490 3340 262496 3352
rect 262548 3340 262554 3392
rect 360654 3340 360660 3392
rect 360712 3380 360718 3392
rect 385678 3380 385684 3392
rect 360712 3352 385684 3380
rect 360712 3340 360718 3352
rect 385678 3340 385684 3352
rect 385736 3340 385742 3392
rect 394234 3340 394240 3392
rect 394292 3380 394298 3392
rect 431957 3383 432015 3389
rect 431957 3380 431969 3383
rect 394292 3352 431969 3380
rect 394292 3340 394298 3352
rect 431957 3349 431969 3352
rect 432003 3349 432015 3383
rect 497366 3380 497372 3392
rect 431957 3343 432015 3349
rect 432064 3352 497372 3380
rect 172848 3284 180794 3312
rect 172848 3272 172854 3284
rect 210050 3272 210056 3324
rect 210108 3312 210114 3324
rect 249058 3312 249064 3324
rect 210108 3284 249064 3312
rect 210108 3272 210114 3284
rect 249058 3272 249064 3284
rect 249116 3272 249122 3324
rect 370682 3272 370688 3324
rect 370740 3312 370746 3324
rect 400861 3315 400919 3321
rect 400861 3312 400873 3315
rect 370740 3284 400873 3312
rect 370740 3272 370746 3284
rect 400861 3281 400873 3284
rect 400907 3281 400919 3315
rect 400861 3275 400919 3281
rect 400950 3272 400956 3324
rect 401008 3312 401014 3324
rect 417421 3315 417479 3321
rect 417421 3312 417433 3315
rect 401008 3284 417433 3312
rect 401008 3272 401014 3284
rect 417421 3281 417433 3284
rect 417467 3281 417479 3315
rect 417421 3275 417479 3281
rect 431218 3272 431224 3324
rect 431276 3312 431282 3324
rect 432064 3312 432092 3352
rect 497366 3340 497372 3352
rect 497424 3340 497430 3392
rect 502702 3312 502708 3324
rect 431276 3284 432092 3312
rect 437952 3284 502708 3312
rect 431276 3272 431282 3284
rect 29178 3204 29184 3256
rect 29236 3244 29242 3256
rect 138106 3244 138112 3256
rect 29236 3216 138112 3244
rect 29236 3204 29242 3216
rect 138106 3204 138112 3216
rect 138164 3204 138170 3256
rect 146202 3204 146208 3256
rect 146260 3244 146266 3256
rect 156693 3247 156751 3253
rect 156693 3244 156705 3247
rect 146260 3216 156705 3244
rect 146260 3204 146266 3216
rect 156693 3213 156705 3216
rect 156739 3213 156751 3247
rect 156693 3207 156751 3213
rect 188798 3204 188804 3256
rect 188856 3244 188862 3256
rect 235626 3244 235632 3256
rect 188856 3216 235632 3244
rect 188856 3204 188862 3216
rect 235626 3204 235632 3216
rect 235684 3204 235690 3256
rect 236638 3204 236644 3256
rect 236696 3244 236702 3256
rect 265894 3244 265900 3256
rect 236696 3216 265900 3244
rect 236696 3204 236702 3216
rect 265894 3204 265900 3216
rect 265952 3204 265958 3256
rect 353938 3204 353944 3256
rect 353996 3244 354002 3256
rect 375006 3244 375012 3256
rect 353996 3216 375012 3244
rect 353996 3204 354002 3216
rect 375006 3204 375012 3216
rect 375064 3204 375070 3256
rect 377398 3204 377404 3256
rect 377456 3244 377462 3256
rect 412266 3244 412272 3256
rect 377456 3216 412272 3244
rect 377456 3204 377462 3216
rect 412266 3204 412272 3216
rect 412324 3204 412330 3256
rect 434622 3204 434628 3256
rect 434680 3244 434686 3256
rect 437952 3244 437980 3284
rect 502702 3272 502708 3284
rect 502760 3272 502766 3324
rect 434680 3216 437980 3244
rect 434680 3204 434686 3216
rect 441246 3204 441252 3256
rect 441304 3244 441310 3256
rect 523954 3244 523960 3256
rect 441304 3216 523960 3244
rect 441304 3204 441310 3216
rect 523954 3204 523960 3216
rect 524012 3204 524018 3256
rect 23842 3136 23848 3188
rect 23900 3176 23906 3188
rect 134794 3176 134800 3188
rect 23900 3148 134800 3176
rect 23900 3136 23906 3148
rect 134794 3136 134800 3148
rect 134852 3136 134858 3188
rect 135530 3136 135536 3188
rect 135588 3176 135594 3188
rect 141789 3179 141847 3185
rect 141789 3176 141801 3179
rect 135588 3148 141801 3176
rect 135588 3136 135594 3148
rect 141789 3145 141801 3148
rect 141835 3145 141847 3179
rect 141789 3139 141847 3145
rect 183462 3136 183468 3188
rect 183520 3176 183526 3188
rect 232222 3176 232228 3188
rect 183520 3148 232228 3176
rect 183520 3136 183526 3148
rect 232222 3136 232228 3148
rect 232280 3136 232286 3188
rect 257982 3136 257988 3188
rect 258040 3176 258046 3188
rect 279326 3176 279332 3188
rect 258040 3148 279332 3176
rect 258040 3136 258046 3148
rect 279326 3136 279332 3148
rect 279384 3136 279390 3188
rect 384114 3136 384120 3188
rect 384172 3176 384178 3188
rect 422846 3176 422852 3188
rect 384172 3148 422852 3176
rect 384172 3136 384178 3148
rect 422846 3136 422852 3148
rect 422904 3136 422910 3188
rect 431957 3179 432015 3185
rect 431957 3145 431969 3179
rect 432003 3176 432015 3179
rect 438854 3176 438860 3188
rect 432003 3148 438860 3176
rect 432003 3145 432015 3148
rect 431957 3139 432015 3145
rect 438854 3136 438860 3148
rect 438912 3136 438918 3188
rect 444282 3136 444288 3188
rect 444340 3176 444346 3188
rect 534626 3176 534632 3188
rect 444340 3148 534632 3176
rect 444340 3136 444346 3148
rect 534626 3136 534632 3148
rect 534684 3136 534690 3188
rect 18506 3068 18512 3120
rect 18564 3108 18570 3120
rect 126977 3111 127035 3117
rect 18564 3080 126928 3108
rect 18564 3068 18570 3080
rect 13170 3000 13176 3052
rect 13228 3040 13234 3052
rect 125597 3043 125655 3049
rect 125597 3040 125609 3043
rect 13228 3012 125609 3040
rect 13228 3000 13234 3012
rect 125597 3009 125609 3012
rect 125643 3009 125655 3043
rect 126900 3040 126928 3080
rect 126977 3077 126989 3111
rect 127023 3108 127035 3111
rect 191926 3108 191932 3120
rect 127023 3080 191932 3108
rect 127023 3077 127035 3080
rect 126977 3071 127035 3077
rect 191926 3068 191932 3080
rect 191984 3068 191990 3120
rect 204714 3068 204720 3120
rect 204772 3108 204778 3120
rect 245654 3108 245660 3120
rect 204772 3080 245660 3108
rect 204772 3068 204778 3080
rect 245654 3068 245660 3080
rect 245712 3068 245718 3120
rect 247310 3068 247316 3120
rect 247368 3108 247374 3120
rect 272610 3108 272616 3120
rect 247368 3080 272616 3108
rect 247368 3068 247374 3080
rect 272610 3068 272616 3080
rect 272668 3068 272674 3120
rect 273898 3068 273904 3120
rect 273956 3108 273962 3120
rect 289354 3108 289360 3120
rect 273956 3080 289360 3108
rect 273956 3068 273962 3080
rect 289354 3068 289360 3080
rect 289412 3068 289418 3120
rect 347222 3068 347228 3120
rect 347280 3108 347286 3120
rect 364334 3108 364340 3120
rect 347280 3080 364340 3108
rect 347280 3068 347286 3080
rect 364334 3068 364340 3080
rect 364392 3068 364398 3120
rect 387518 3068 387524 3120
rect 387576 3108 387582 3120
rect 428182 3108 428188 3120
rect 387576 3080 428188 3108
rect 387576 3068 387582 3080
rect 428182 3068 428188 3080
rect 428240 3068 428246 3120
rect 448054 3068 448060 3120
rect 448112 3108 448118 3120
rect 555878 3108 555884 3120
rect 448112 3080 555884 3108
rect 448112 3068 448118 3080
rect 555878 3068 555884 3080
rect 555936 3068 555942 3120
rect 127253 3043 127311 3049
rect 127253 3040 127265 3043
rect 126900 3012 127265 3040
rect 125597 3003 125655 3009
rect 127253 3009 127265 3012
rect 127299 3009 127311 3043
rect 127253 3003 127311 3009
rect 127437 3043 127495 3049
rect 127437 3009 127449 3043
rect 127483 3040 127495 3043
rect 188522 3040 188528 3052
rect 127483 3012 188528 3040
rect 127483 3009 127495 3012
rect 127437 3003 127495 3009
rect 188522 3000 188528 3012
rect 188580 3000 188586 3052
rect 199378 3000 199384 3052
rect 199436 3040 199442 3052
rect 242342 3040 242348 3052
rect 199436 3012 242348 3040
rect 199436 3000 199442 3012
rect 242342 3000 242348 3012
rect 242400 3000 242406 3052
rect 252646 3000 252652 3052
rect 252704 3040 252710 3052
rect 276014 3040 276020 3052
rect 252704 3012 276020 3040
rect 252704 3000 252710 3012
rect 276014 3000 276020 3012
rect 276072 3000 276078 3052
rect 279234 3000 279240 3052
rect 279292 3040 279298 3052
rect 292758 3040 292764 3052
rect 279292 3012 292764 3040
rect 279292 3000 279298 3012
rect 292758 3000 292764 3012
rect 292816 3000 292822 3052
rect 295150 3000 295156 3052
rect 295208 3040 295214 3052
rect 302878 3040 302884 3052
rect 295208 3012 302884 3040
rect 295208 3000 295214 3012
rect 302878 3000 302884 3012
rect 302936 3000 302942 3052
rect 357250 3000 357256 3052
rect 357308 3040 357314 3052
rect 380342 3040 380348 3052
rect 357308 3012 380348 3040
rect 357308 3000 357314 3012
rect 380342 3000 380348 3012
rect 380400 3000 380406 3052
rect 390922 3000 390928 3052
rect 390980 3040 390986 3052
rect 433518 3040 433524 3052
rect 390980 3012 433524 3040
rect 390980 3000 390986 3012
rect 433518 3000 433524 3012
rect 433576 3000 433582 3052
rect 451182 3000 451188 3052
rect 451240 3040 451246 3052
rect 561214 3040 561220 3052
rect 451240 3012 561220 3040
rect 451240 3000 451246 3012
rect 561214 3000 561220 3012
rect 561272 3000 561278 3052
rect 103606 2932 103612 2984
rect 103664 2972 103670 2984
rect 181806 2972 181812 2984
rect 103664 2944 181812 2972
rect 103664 2932 103670 2944
rect 181806 2932 181812 2944
rect 181864 2932 181870 2984
rect 194134 2932 194140 2984
rect 194192 2972 194198 2984
rect 238938 2972 238944 2984
rect 194192 2944 238944 2972
rect 194192 2932 194198 2944
rect 238938 2932 238944 2944
rect 238996 2932 239002 2984
rect 263226 2932 263232 2984
rect 263284 2972 263290 2984
rect 282914 2972 282920 2984
rect 263284 2944 282920 2972
rect 263284 2932 263290 2944
rect 282914 2932 282920 2944
rect 282972 2932 282978 2984
rect 289906 2932 289912 2984
rect 289964 2972 289970 2984
rect 299474 2972 299480 2984
rect 289964 2944 299480 2972
rect 289964 2932 289970 2944
rect 299474 2932 299480 2944
rect 299532 2932 299538 2984
rect 363966 2932 363972 2984
rect 364024 2972 364030 2984
rect 390830 2972 390836 2984
rect 364024 2944 390836 2972
rect 364024 2932 364030 2944
rect 390830 2932 390836 2944
rect 390888 2932 390894 2984
rect 397270 2932 397276 2984
rect 397328 2972 397334 2984
rect 444190 2972 444196 2984
rect 397328 2944 444196 2972
rect 397328 2932 397334 2944
rect 444190 2932 444196 2944
rect 444248 2932 444254 2984
rect 454770 2932 454776 2984
rect 454828 2972 454834 2984
rect 571886 2972 571892 2984
rect 454828 2944 571892 2972
rect 454828 2932 454834 2944
rect 571886 2932 571892 2944
rect 571944 2932 571950 2984
rect 49326 2864 49332 2916
rect 49384 2904 49390 2916
rect 114465 2907 114523 2913
rect 114465 2904 114477 2907
rect 49384 2876 114477 2904
rect 49384 2864 49390 2876
rect 114465 2873 114477 2876
rect 114511 2873 114523 2907
rect 114465 2867 114523 2873
rect 114554 2864 114560 2916
rect 114612 2904 114618 2916
rect 115474 2904 115480 2916
rect 114612 2876 115480 2904
rect 114612 2864 114618 2876
rect 115474 2864 115480 2876
rect 115532 2864 115538 2916
rect 119614 2864 119620 2916
rect 119672 2904 119678 2916
rect 121641 2907 121699 2913
rect 119672 2876 121592 2904
rect 119672 2864 119678 2876
rect 2590 2796 2596 2848
rect 2648 2836 2654 2848
rect 121454 2836 121460 2848
rect 2648 2808 121460 2836
rect 2648 2796 2654 2808
rect 121454 2796 121460 2808
rect 121512 2796 121518 2848
rect 121564 2836 121592 2876
rect 121641 2873 121653 2907
rect 121687 2904 121699 2907
rect 127437 2907 127495 2913
rect 127437 2904 127449 2907
rect 121687 2876 127449 2904
rect 121687 2873 121699 2876
rect 121641 2867 121699 2873
rect 127437 2873 127449 2876
rect 127483 2873 127495 2907
rect 127437 2867 127495 2873
rect 127621 2907 127679 2913
rect 127621 2873 127633 2907
rect 127667 2904 127679 2907
rect 464154 2904 464160 2916
rect 127667 2876 464160 2904
rect 127667 2873 127679 2876
rect 127621 2867 127679 2873
rect 464154 2864 464160 2876
rect 464212 2864 464218 2916
rect 126977 2839 127035 2845
rect 126977 2836 126989 2839
rect 121564 2808 126989 2836
rect 126977 2805 126989 2808
rect 127023 2805 127035 2839
rect 126977 2799 127035 2805
rect 127253 2839 127311 2845
rect 127253 2805 127265 2839
rect 127299 2836 127311 2839
rect 131390 2836 131396 2848
rect 127299 2808 131396 2836
rect 127299 2805 127311 2808
rect 127253 2799 127311 2805
rect 131390 2796 131396 2808
rect 131448 2796 131454 2848
rect 156874 2796 156880 2848
rect 156932 2836 156938 2848
rect 215478 2836 215484 2848
rect 156932 2808 215484 2836
rect 156932 2796 156938 2808
rect 215478 2796 215484 2808
rect 215536 2796 215542 2848
rect 220722 2796 220728 2848
rect 220780 2836 220786 2848
rect 255774 2836 255780 2848
rect 220780 2808 255780 2836
rect 220780 2796 220786 2808
rect 255774 2796 255780 2808
rect 255832 2796 255838 2848
rect 268562 2796 268568 2848
rect 268620 2836 268626 2848
rect 268620 2808 281856 2836
rect 268620 2796 268626 2808
rect 55950 2728 55956 2780
rect 56008 2768 56014 2780
rect 66162 2768 66168 2780
rect 56008 2740 66168 2768
rect 56008 2728 56014 2740
rect 66162 2728 66168 2740
rect 66220 2728 66226 2780
rect 85942 2728 85948 2780
rect 86000 2768 86006 2780
rect 86000 2740 103514 2768
rect 86000 2728 86006 2740
rect 103486 2700 103514 2740
rect 108942 2728 108948 2780
rect 109000 2768 109006 2780
rect 115382 2768 115388 2780
rect 109000 2740 115388 2768
rect 109000 2728 109006 2740
rect 115382 2728 115388 2740
rect 115440 2728 115446 2780
rect 116854 2728 116860 2780
rect 116912 2768 116918 2780
rect 144914 2768 144920 2780
rect 116912 2740 144920 2768
rect 116912 2728 116918 2740
rect 144914 2728 144920 2740
rect 144972 2728 144978 2780
rect 146938 2728 146944 2780
rect 146996 2768 147002 2780
rect 151814 2768 151820 2780
rect 146996 2740 151820 2768
rect 146996 2728 147002 2740
rect 151814 2728 151820 2740
rect 151872 2728 151878 2780
rect 281828 2768 281856 2808
rect 284570 2796 284576 2848
rect 284628 2836 284634 2848
rect 284628 2808 294000 2836
rect 284628 2796 284634 2808
rect 286042 2768 286048 2780
rect 281828 2740 286048 2768
rect 286042 2728 286048 2740
rect 286100 2728 286106 2780
rect 293972 2768 294000 2808
rect 300486 2796 300492 2848
rect 300544 2836 300550 2848
rect 300544 2808 303660 2836
rect 300544 2796 300550 2808
rect 296070 2768 296076 2780
rect 293972 2740 296076 2768
rect 296070 2728 296076 2740
rect 296128 2728 296134 2780
rect 303632 2768 303660 2808
rect 305822 2796 305828 2848
rect 305880 2836 305886 2848
rect 309594 2836 309600 2848
rect 305880 2808 309600 2836
rect 305880 2796 305886 2808
rect 309594 2796 309600 2808
rect 309652 2796 309658 2848
rect 320174 2796 320180 2848
rect 320232 2836 320238 2848
rect 321830 2836 321836 2848
rect 320232 2808 321836 2836
rect 320232 2796 320238 2808
rect 321830 2796 321836 2808
rect 321888 2796 321894 2848
rect 325666 2808 327028 2836
rect 306374 2768 306380 2780
rect 303632 2740 306380 2768
rect 306374 2728 306380 2740
rect 306432 2728 306438 2780
rect 323670 2728 323676 2780
rect 323728 2768 323734 2780
rect 325666 2768 325694 2808
rect 323728 2740 325694 2768
rect 323728 2728 323734 2740
rect 114554 2700 114560 2712
rect 103486 2672 114560 2700
rect 114554 2660 114560 2672
rect 114612 2660 114618 2712
rect 114646 2660 114652 2712
rect 114704 2700 114710 2712
rect 141510 2700 141516 2712
rect 114704 2672 141516 2700
rect 114704 2660 114710 2672
rect 141510 2660 141516 2672
rect 141568 2660 141574 2712
rect 141602 2660 141608 2712
rect 141660 2700 141666 2712
rect 148226 2700 148232 2712
rect 141660 2672 148232 2700
rect 141660 2660 141666 2672
rect 148226 2660 148232 2672
rect 148284 2660 148290 2712
rect 327000 2700 327028 2808
rect 327074 2796 327080 2848
rect 327132 2836 327138 2848
rect 332410 2836 332416 2848
rect 327132 2808 332416 2836
rect 327132 2796 327138 2808
rect 332410 2796 332416 2808
rect 332468 2796 332474 2848
rect 337746 2836 337752 2848
rect 332520 2808 337752 2836
rect 330386 2728 330392 2780
rect 330444 2768 330450 2780
rect 332520 2768 332548 2808
rect 337746 2796 337752 2808
rect 337804 2796 337810 2848
rect 350442 2796 350448 2848
rect 350500 2836 350506 2848
rect 369670 2836 369676 2848
rect 350500 2808 369676 2836
rect 350500 2796 350506 2808
rect 369670 2796 369676 2808
rect 369728 2796 369734 2848
rect 380802 2796 380808 2848
rect 380860 2836 380866 2848
rect 417421 2839 417479 2845
rect 380860 2808 417372 2836
rect 380860 2796 380866 2808
rect 330444 2740 332548 2768
rect 417344 2768 417372 2808
rect 417421 2805 417433 2839
rect 417467 2836 417479 2839
rect 449526 2836 449532 2848
rect 417467 2808 449532 2836
rect 417467 2805 417479 2808
rect 417421 2799 417479 2805
rect 449526 2796 449532 2808
rect 449584 2796 449590 2848
rect 458174 2796 458180 2848
rect 458232 2836 458238 2848
rect 513374 2836 513380 2848
rect 458232 2808 513380 2836
rect 458232 2796 458238 2808
rect 513374 2796 513380 2808
rect 513432 2796 513438 2848
rect 417602 2768 417608 2780
rect 417344 2740 417608 2768
rect 330444 2728 330450 2740
rect 417602 2728 417608 2740
rect 417660 2728 417666 2780
rect 426342 2728 426348 2780
rect 426400 2768 426406 2780
rect 467834 2768 467840 2780
rect 426400 2740 467840 2768
rect 426400 2728 426406 2740
rect 467834 2728 467840 2740
rect 467892 2728 467898 2780
rect 327074 2700 327080 2712
rect 327000 2672 327080 2700
rect 327074 2660 327080 2672
rect 327132 2660 327138 2712
rect 337102 2660 337108 2712
rect 337160 2700 337166 2712
rect 348418 2700 348424 2712
rect 337160 2672 348424 2700
rect 337160 2660 337166 2672
rect 348418 2660 348424 2672
rect 348476 2660 348482 2712
rect 437934 2660 437940 2712
rect 437992 2700 437998 2712
rect 458174 2700 458180 2712
rect 437992 2672 458180 2700
rect 437992 2660 437998 2672
rect 458174 2660 458180 2672
rect 458232 2660 458238 2712
rect 35802 2592 35808 2644
rect 35860 2632 35866 2644
rect 519630 2632 519636 2644
rect 35860 2604 519636 2632
rect 35860 2592 35866 2604
rect 519630 2592 519636 2604
rect 519688 2592 519694 2644
rect 15930 2524 15936 2576
rect 15988 2564 15994 2576
rect 477678 2564 477684 2576
rect 15988 2536 477684 2564
rect 15988 2524 15994 2536
rect 477678 2524 477684 2536
rect 477736 2524 477742 2576
rect 25958 2456 25964 2508
rect 26016 2496 26022 2508
rect 487706 2496 487712 2508
rect 26016 2468 487712 2496
rect 26016 2456 26022 2468
rect 487706 2456 487712 2468
rect 487764 2456 487770 2508
rect 1302 2388 1308 2440
rect 1360 2428 1366 2440
rect 58618 2428 58624 2440
rect 1360 2400 58624 2428
rect 1360 2388 1366 2400
rect 58618 2388 58624 2400
rect 58676 2388 58682 2440
rect 68922 2388 68928 2440
rect 68980 2428 68986 2440
rect 86862 2428 86868 2440
rect 68980 2400 86868 2428
rect 68980 2388 68986 2400
rect 86862 2388 86868 2400
rect 86920 2388 86926 2440
rect 92382 2388 92388 2440
rect 92440 2428 92446 2440
rect 520366 2428 520372 2440
rect 92440 2400 520372 2428
rect 92440 2388 92446 2400
rect 520366 2388 520372 2400
rect 520424 2388 520430 2440
rect 79318 2320 79324 2372
rect 79376 2360 79382 2372
rect 504542 2360 504548 2372
rect 79376 2332 504548 2360
rect 79376 2320 79382 2332
rect 504542 2320 504548 2332
rect 504600 2320 504606 2372
rect 99282 2252 99288 2304
rect 99340 2292 99346 2304
rect 520458 2292 520464 2304
rect 99340 2264 520464 2292
rect 99340 2252 99346 2264
rect 520458 2252 520464 2264
rect 520516 2252 520522 2304
rect 89346 2184 89352 2236
rect 89404 2224 89410 2236
rect 507854 2224 507860 2236
rect 89404 2196 507860 2224
rect 89404 2184 89410 2196
rect 507854 2184 507860 2196
rect 507912 2184 507918 2236
rect 95970 2116 95976 2168
rect 96028 2156 96034 2168
rect 511258 2156 511264 2168
rect 96028 2128 511264 2156
rect 96028 2116 96034 2128
rect 511258 2116 511264 2128
rect 511316 2116 511322 2168
rect 102686 2048 102692 2100
rect 102744 2088 102750 2100
rect 517974 2088 517980 2100
rect 102744 2060 517980 2088
rect 102744 2048 102750 2060
rect 517974 2048 517980 2060
rect 518032 2048 518038 2100
rect 115198 1980 115204 2032
rect 115256 2020 115262 2032
rect 514754 2020 514760 2032
rect 115256 1992 514760 2020
rect 115256 1980 115262 1992
rect 514754 1980 514760 1992
rect 514812 1980 514818 2032
rect 82630 1912 82636 1964
rect 82688 1952 82694 1964
rect 115566 1952 115572 1964
rect 82688 1924 115572 1952
rect 82688 1912 82694 1924
rect 115566 1912 115572 1924
rect 115624 1912 115630 1964
rect 116486 1912 116492 1964
rect 116544 1952 116550 1964
rect 501138 1952 501144 1964
rect 116544 1924 501144 1952
rect 116544 1912 116550 1924
rect 501138 1912 501144 1924
rect 501196 1912 501202 1964
rect 113818 1844 113824 1896
rect 113876 1884 113882 1896
rect 491294 1884 491300 1896
rect 113876 1856 491300 1884
rect 113876 1844 113882 1856
rect 491294 1844 491300 1856
rect 491352 1844 491358 1896
rect 22646 1776 22652 1828
rect 22704 1816 22710 1828
rect 116578 1816 116584 1828
rect 22704 1788 116584 1816
rect 22704 1776 22710 1788
rect 116578 1776 116584 1788
rect 116636 1776 116642 1828
rect 117682 1776 117688 1828
rect 117740 1816 117746 1828
rect 494422 1816 494428 1828
rect 117740 1788 494428 1816
rect 117740 1776 117746 1788
rect 494422 1776 494428 1788
rect 494480 1776 494486 1828
rect 118142 1708 118148 1760
rect 118200 1748 118206 1760
rect 484394 1748 484400 1760
rect 118200 1720 484400 1748
rect 118200 1708 118206 1720
rect 484394 1708 484400 1720
rect 484452 1708 484458 1760
rect 168834 1640 168840 1692
rect 168892 1680 168898 1692
rect 480990 1680 480996 1692
rect 168892 1652 480996 1680
rect 168892 1640 168898 1652
rect 480990 1640 480996 1652
rect 481048 1640 481054 1692
rect 9306 1572 9312 1624
rect 9364 1612 9370 1624
rect 176654 1612 176660 1624
rect 9364 1584 176660 1612
rect 9364 1572 9370 1584
rect 176654 1572 176660 1584
rect 176712 1572 176718 1624
rect 333698 1572 333704 1624
rect 333756 1612 333762 1624
rect 343082 1612 343088 1624
rect 333756 1584 343088 1612
rect 333756 1572 333762 1584
rect 343082 1572 343088 1584
rect 343140 1572 343146 1624
rect 343450 1572 343456 1624
rect 343508 1612 343514 1624
rect 358998 1612 359004 1624
rect 343508 1584 359004 1612
rect 343508 1572 343514 1584
rect 358998 1572 359004 1584
rect 359056 1572 359062 1624
rect 105998 1504 106004 1556
rect 106056 1544 106062 1556
rect 213822 1544 213828 1556
rect 106056 1516 213828 1544
rect 106056 1504 106062 1516
rect 213822 1504 213828 1516
rect 213880 1504 213886 1556
rect 340414 1504 340420 1556
rect 340472 1544 340478 1556
rect 353754 1544 353760 1556
rect 340472 1516 353760 1544
rect 340472 1504 340478 1516
rect 353754 1504 353760 1516
rect 353812 1504 353818 1556
rect 32582 1436 32588 1488
rect 32640 1476 32646 1488
rect 520734 1476 520740 1488
rect 32640 1448 520740 1476
rect 32640 1436 32646 1448
rect 520734 1436 520740 1448
rect 520792 1436 520798 1488
rect 19242 1368 19248 1420
rect 19300 1408 19306 1420
rect 520090 1408 520096 1420
rect 19300 1380 520096 1408
rect 19300 1368 19306 1380
rect 520090 1368 520096 1380
rect 520148 1368 520154 1420
rect 72602 1300 72608 1352
rect 72660 1340 72666 1352
rect 497826 1340 497832 1352
rect 72660 1312 497832 1340
rect 72660 1300 72666 1312
rect 497826 1300 497832 1312
rect 497884 1300 497890 1352
rect 71590 76 71596 128
rect 71648 116 71654 128
rect 161658 116 161664 128
rect 71648 88 161664 116
rect 71648 76 71654 88
rect 161658 76 161664 88
rect 161716 76 161722 128
rect 34606 8 34612 60
rect 34664 48 34670 60
rect 457438 48 457444 60
rect 34664 20 457444 48
rect 34664 8 34670 20
rect 457438 8 457444 20
rect 457496 8 457502 60
<< via1 >>
rect 26792 158856 26844 158908
rect 137468 158856 137520 158908
rect 15200 158788 15252 158840
rect 129740 158788 129792 158840
rect 22836 158720 22888 158772
rect 134892 158720 134944 158772
rect 11152 158652 11204 158704
rect 127072 158652 127124 158704
rect 82820 158584 82872 158636
rect 164240 158584 164292 158636
rect 70400 158516 70452 158568
rect 156328 158516 156380 158568
rect 75000 158448 75052 158500
rect 161664 158448 161716 158500
rect 67364 158380 67416 158432
rect 153752 158380 153804 158432
rect 51080 158312 51132 158364
rect 148692 158312 148744 158364
rect 34520 158244 34572 158296
rect 142804 158244 142856 158296
rect 12440 158176 12492 158228
rect 122840 158176 122892 158228
rect 18972 158108 19024 158160
rect 132592 158108 132644 158160
rect 112536 158040 112588 158092
rect 194784 158040 194836 158092
rect 94044 157972 94096 158024
rect 182364 157972 182416 158024
rect 82268 157904 82320 157956
rect 174544 157904 174596 157956
rect 58900 157836 58952 157888
rect 158996 157836 159048 157888
rect 47216 157768 47268 157820
rect 151176 157768 151228 157820
rect 38476 157700 38528 157752
rect 145288 157700 145340 157752
rect 148600 157700 148652 157752
rect 218888 157700 218940 157752
rect 30656 157632 30708 157684
rect 140136 157632 140188 157684
rect 140780 157632 140832 157684
rect 214104 157632 214156 157684
rect 129096 157564 129148 157616
rect 205824 157564 205876 157616
rect 113548 157496 113600 157548
rect 195428 157496 195480 157548
rect 104716 157428 104768 157480
rect 189632 157428 189684 157480
rect 119436 157360 119488 157412
rect 511540 157360 511592 157412
rect 73528 157292 73580 157344
rect 168748 157292 168800 157344
rect 181076 157292 181128 157344
rect 189540 157292 189592 157344
rect 246120 157292 246172 157344
rect 426256 157292 426308 157344
rect 458548 157292 458600 157344
rect 475016 157292 475068 157344
rect 68652 157224 68704 157276
rect 165620 157224 165672 157276
rect 170680 157224 170732 157276
rect 65708 157156 65760 157208
rect 163504 157156 163556 157208
rect 167092 157156 167144 157208
rect 175924 157224 175976 157276
rect 237012 157224 237064 157276
rect 428924 157224 428976 157276
rect 462504 157224 462556 157276
rect 473728 157224 473780 157276
rect 176016 157156 176068 157208
rect 177856 157156 177908 157208
rect 238392 157156 238444 157208
rect 436652 157156 436704 157208
rect 474188 157156 474240 157208
rect 57980 157088 58032 157140
rect 158444 157088 158496 157140
rect 163044 157088 163096 157140
rect 173900 157088 173952 157140
rect 236000 157088 236052 157140
rect 251916 157088 251968 157140
rect 287796 157088 287848 157140
rect 438032 157088 438084 157140
rect 476120 157088 476172 157140
rect 56968 157020 57020 157072
rect 157708 157020 157760 157072
rect 160100 157020 160152 157072
rect 166172 157020 166224 157072
rect 230572 157020 230624 157072
rect 244096 157020 244148 157072
rect 282552 157020 282604 157072
rect 437388 157020 437440 157072
rect 475108 157020 475160 157072
rect 477316 157224 477368 157276
rect 529756 157292 529808 157344
rect 531688 157224 531740 157276
rect 535552 157156 535604 157208
rect 478788 157088 478840 157140
rect 537484 157088 537536 157140
rect 541440 157020 541492 157072
rect 53104 156952 53156 157004
rect 155040 156952 155092 157004
rect 158352 156952 158404 157004
rect 225328 156952 225380 157004
rect 236276 156952 236328 157004
rect 277492 156952 277544 157004
rect 442540 156952 442592 157004
rect 482928 156952 482980 157004
rect 483020 156952 483072 157004
rect 543372 156952 543424 157004
rect 42340 156884 42392 156936
rect 147956 156884 148008 156936
rect 150532 156884 150584 156936
rect 220084 156884 220136 156936
rect 228548 156884 228600 156936
rect 272156 156884 272208 156936
rect 442816 156884 442868 156936
rect 483940 156884 483992 156936
rect 485504 156884 485556 156936
rect 547236 156884 547288 156936
rect 25780 156816 25832 156868
rect 136824 156816 136876 156868
rect 139860 156816 139912 156868
rect 213000 156816 213052 156868
rect 218796 156816 218848 156868
rect 265624 156816 265676 156868
rect 445116 156816 445168 156868
rect 486792 156816 486844 156868
rect 486884 156816 486936 156868
rect 549168 156816 549220 156868
rect 17960 156748 18012 156800
rect 131672 156748 131724 156800
rect 134984 156748 135036 156800
rect 209872 156748 209924 156800
rect 218152 156748 218204 156800
rect 221740 156748 221792 156800
rect 267832 156748 267884 156800
rect 445668 156748 445720 156800
rect 487804 156748 487856 156800
rect 490656 156748 490708 156800
rect 555056 156748 555108 156800
rect 10140 156680 10192 156732
rect 126428 156680 126480 156732
rect 132040 156680 132092 156732
rect 207756 156680 207808 156732
rect 212908 156680 212960 156732
rect 261760 156680 261812 156732
rect 449072 156680 449124 156732
rect 492680 156680 492732 156732
rect 493324 156680 493376 156732
rect 558920 156680 558972 156732
rect 6276 156612 6328 156664
rect 123852 156612 123904 156664
rect 124220 156612 124272 156664
rect 202512 156612 202564 156664
rect 209044 156612 209096 156664
rect 259092 156612 259144 156664
rect 420736 156612 420788 156664
rect 450728 156612 450780 156664
rect 456708 156612 456760 156664
rect 504364 156612 504416 156664
rect 508780 156612 508832 156664
rect 577504 156612 577556 156664
rect 76472 156544 76524 156596
rect 223580 156544 223632 156596
rect 469864 156544 469916 156596
rect 523868 156544 523920 156596
rect 81348 156476 81400 156528
rect 84292 156408 84344 156460
rect 231124 156476 231176 156528
rect 466000 156476 466052 156528
rect 517980 156476 518032 156528
rect 173716 156408 173768 156460
rect 225972 156408 226024 156460
rect 440608 156408 440660 156460
rect 479984 156408 480036 156460
rect 480076 156408 480128 156460
rect 530676 156408 530728 156460
rect 92020 156340 92072 156392
rect 178776 156340 178828 156392
rect 180892 156340 180944 156392
rect 191564 156340 191616 156392
rect 193404 156340 193456 156392
rect 248696 156340 248748 156392
rect 481548 156340 481600 156392
rect 487160 156340 487212 156392
rect 538496 156340 538548 156392
rect 99840 156272 99892 156324
rect 186504 156272 186556 156324
rect 197360 156272 197412 156324
rect 251364 156272 251416 156324
rect 460664 156272 460716 156324
rect 510252 156272 510304 156324
rect 107660 156204 107712 156256
rect 180892 156204 180944 156256
rect 183468 156204 183520 156256
rect 236368 156204 236420 156256
rect 453580 156204 453632 156256
rect 499488 156204 499540 156256
rect 111524 156136 111576 156188
rect 116400 156068 116452 156120
rect 191748 156136 191800 156188
rect 241612 156136 241664 156188
rect 452292 156136 452344 156188
rect 497556 156136 497608 156188
rect 119344 156000 119396 156052
rect 194048 156068 194100 156120
rect 199384 156068 199436 156120
rect 244372 156068 244424 156120
rect 450360 156068 450412 156120
rect 494612 156068 494664 156120
rect 197452 156000 197504 156052
rect 205640 156000 205692 156052
rect 155868 155932 155920 155984
rect 12164 155864 12216 155916
rect 4344 155796 4396 155848
rect 12440 155796 12492 155848
rect 33600 155864 33652 155916
rect 34704 155864 34756 155916
rect 66720 155864 66772 155916
rect 82820 155864 82872 155916
rect 176844 155864 176896 155916
rect 179144 155864 179196 155916
rect 180800 155864 180852 155916
rect 183376 155864 183428 155916
rect 17868 155796 17920 155848
rect 43352 155796 43404 155848
rect 51080 155796 51132 155848
rect 63776 155796 63828 155848
rect 186412 155864 186464 155916
rect 186596 155864 186648 155916
rect 200212 155864 200264 155916
rect 202788 155864 202840 155916
rect 206100 155864 206152 155916
rect 257160 156000 257212 156052
rect 446496 156000 446548 156052
rect 488816 156000 488868 156052
rect 249340 155932 249392 155984
rect 215852 155864 215904 155916
rect 216588 155864 216640 155916
rect 55956 155728 56008 155780
rect 136916 155728 136968 155780
rect 143724 155728 143776 155780
rect 144644 155728 144696 155780
rect 144736 155728 144788 155780
rect 149612 155728 149664 155780
rect 153108 155728 153160 155780
rect 153476 155728 153528 155780
rect 155408 155728 155460 155780
rect 160100 155728 160152 155780
rect 160284 155728 160336 155780
rect 74540 155660 74592 155712
rect 167736 155660 167788 155712
rect 171048 155660 171100 155712
rect 172152 155728 172204 155780
rect 219716 155728 219768 155780
rect 222108 155728 222160 155780
rect 222660 155864 222712 155916
rect 258724 155864 258776 155916
rect 262128 155864 262180 155916
rect 229468 155796 229520 155848
rect 225052 155728 225104 155780
rect 225604 155728 225656 155780
rect 241152 155796 241204 155848
rect 280252 155864 280304 155916
rect 171968 155660 172020 155712
rect 233424 155660 233476 155712
rect 243176 155660 243228 155712
rect 281448 155796 281500 155848
rect 284116 155864 284168 155916
rect 291752 155864 291804 155916
rect 292856 155864 292908 155916
rect 447784 155932 447836 155984
rect 490748 155932 490800 155984
rect 313740 155864 313792 155916
rect 316224 155864 316276 155916
rect 328460 155864 328512 155916
rect 328920 155864 328972 155916
rect 334348 155864 334400 155916
rect 334808 155864 334860 155916
rect 340236 155864 340288 155916
rect 353300 155864 353352 155916
rect 355416 155864 355468 155916
rect 382372 155864 382424 155916
rect 385500 155864 385552 155916
rect 388444 155864 388496 155916
rect 393228 155864 393280 155916
rect 404176 155864 404228 155916
rect 406936 155864 406988 155916
rect 426348 155864 426400 155916
rect 284392 155796 284444 155848
rect 286968 155796 287020 155848
rect 311256 155796 311308 155848
rect 315304 155796 315356 155848
rect 329656 155796 329708 155848
rect 330852 155796 330904 155848
rect 336556 155796 336608 155848
rect 354220 155796 354272 155848
rect 355968 155796 356020 155848
rect 387340 155796 387392 155848
rect 391296 155796 391348 155848
rect 402244 155796 402296 155848
rect 422484 155796 422536 155848
rect 424968 155796 425020 155848
rect 425612 155796 425664 155848
rect 457628 155864 457680 155916
rect 466276 155864 466328 155916
rect 518992 155864 519044 155916
rect 546500 155864 546552 155916
rect 548248 155864 548300 155916
rect 428280 155796 428332 155848
rect 263784 155728 263836 155780
rect 264612 155728 264664 155780
rect 268476 155728 268528 155780
rect 39396 155592 39448 155644
rect 182732 155592 182784 155644
rect 191472 155592 191524 155644
rect 239220 155592 239272 155644
rect 241428 155592 241480 155644
rect 16028 155524 16080 155576
rect 117964 155524 118016 155576
rect 118332 155524 118384 155576
rect 187792 155524 187844 155576
rect 190552 155524 190604 155576
rect 195336 155524 195388 155576
rect 245108 155592 245160 155644
rect 242164 155524 242216 155576
rect 278228 155728 278280 155780
rect 305000 155728 305052 155780
rect 305552 155728 305604 155780
rect 323492 155728 323544 155780
rect 331864 155728 331916 155780
rect 337936 155728 337988 155780
rect 385500 155728 385552 155780
rect 390284 155728 390336 155780
rect 405832 155728 405884 155780
rect 409788 155728 409840 155780
rect 411352 155728 411404 155780
rect 412732 155728 412784 155780
rect 413284 155728 413336 155780
rect 414664 155728 414716 155780
rect 428372 155728 428424 155780
rect 456616 155796 456668 155848
rect 469128 155796 469180 155848
rect 522856 155796 522908 155848
rect 461492 155728 461544 155780
rect 471152 155728 471204 155780
rect 525800 155728 525852 155780
rect 282920 155660 282972 155712
rect 283104 155660 283156 155712
rect 305920 155660 305972 155712
rect 313372 155660 313424 155712
rect 314292 155660 314344 155712
rect 329380 155660 329432 155712
rect 404820 155660 404872 155712
rect 411260 155660 411312 155712
rect 413744 155660 413796 155712
rect 414112 155660 414164 155712
rect 416688 155660 416740 155712
rect 430304 155660 430356 155712
rect 430396 155660 430448 155712
rect 464436 155660 464488 155712
rect 475752 155660 475804 155712
rect 532608 155660 532660 155712
rect 250904 155592 250956 155644
rect 262772 155592 262824 155644
rect 295524 155592 295576 155644
rect 295800 155592 295852 155644
rect 317052 155592 317104 155644
rect 317236 155592 317288 155644
rect 331312 155592 331364 155644
rect 333796 155592 333848 155644
rect 338948 155592 339000 155644
rect 342536 155592 342588 155644
rect 348240 155592 348292 155644
rect 379704 155592 379756 155644
rect 382556 155592 382608 155644
rect 404084 155592 404136 155644
rect 425428 155592 425480 155644
rect 427636 155592 427688 155644
rect 249984 155524 250036 155576
rect 280160 155524 280212 155576
rect 290832 155524 290884 155576
rect 290924 155524 290976 155576
rect 311900 155524 311952 155576
rect 313280 155524 313332 155576
rect 328736 155524 328788 155576
rect 329932 155524 329984 155576
rect 335636 155524 335688 155576
rect 335728 155524 335780 155576
rect 340972 155524 341024 155576
rect 345480 155524 345532 155576
rect 347596 155524 347648 155576
rect 356244 155524 356296 155576
rect 357440 155524 357492 155576
rect 358176 155524 358228 155576
rect 358820 155524 358872 155576
rect 378140 155524 378192 155576
rect 380624 155524 380676 155576
rect 386328 155524 386380 155576
rect 389364 155524 389416 155576
rect 406752 155524 406804 155576
rect 429292 155524 429344 155576
rect 460480 155592 460532 155644
rect 478328 155592 478380 155644
rect 536564 155592 536616 155644
rect 571984 155592 572036 155644
rect 576492 155592 576544 155644
rect 430488 155524 430540 155576
rect 465356 155524 465408 155576
rect 480904 155524 480956 155576
rect 540428 155524 540480 155576
rect 573364 155524 573416 155576
rect 574560 155524 574612 155576
rect 27712 155456 27764 155508
rect 23848 155388 23900 155440
rect 125232 155388 125284 155440
rect 19892 155320 19944 155372
rect 126060 155320 126112 155372
rect 126152 155320 126204 155372
rect 132960 155456 133012 155508
rect 137836 155456 137888 155508
rect 147588 155456 147640 155508
rect 155868 155456 155920 155508
rect 135168 155388 135220 155440
rect 144736 155388 144788 155440
rect 144828 155388 144880 155440
rect 146760 155388 146812 155440
rect 158720 155456 158772 155508
rect 159272 155456 159324 155508
rect 163044 155456 163096 155508
rect 164148 155456 164200 155508
rect 229284 155456 229336 155508
rect 230480 155456 230532 155508
rect 233148 155456 233200 155508
rect 265072 155456 265124 155508
rect 265532 155456 265584 155508
rect 266452 155456 266504 155508
rect 266544 155456 266596 155508
rect 274364 155456 274416 155508
rect 162124 155388 162176 155440
rect 163228 155388 163280 155440
rect 165528 155388 165580 155440
rect 226524 155388 226576 155440
rect 226616 155388 226668 155440
rect 233240 155388 233292 155440
rect 234620 155388 234672 155440
rect 238300 155388 238352 155440
rect 133788 155320 133840 155372
rect 133972 155320 134024 155372
rect 209044 155320 209096 155372
rect 210976 155320 211028 155372
rect 253204 155320 253256 155372
rect 279148 155388 279200 155440
rect 279240 155388 279292 155440
rect 296720 155388 296772 155440
rect 296904 155456 296956 155508
rect 308404 155456 308456 155508
rect 308496 155456 308548 155508
rect 324412 155456 324464 155508
rect 325976 155456 326028 155508
rect 337200 155456 337252 155508
rect 337660 155456 337712 155508
rect 342536 155456 342588 155508
rect 344560 155456 344612 155508
rect 349528 155456 349580 155508
rect 380900 155456 380952 155508
rect 384488 155456 384540 155508
rect 384764 155456 384816 155508
rect 388352 155456 388404 155508
rect 404636 155456 404688 155508
rect 407856 155456 407908 155508
rect 408316 155456 408368 155508
rect 432236 155456 432288 155508
rect 433064 155456 433116 155508
rect 469312 155456 469364 155508
rect 484860 155456 484912 155508
rect 546316 155456 546368 155508
rect 277308 155320 277360 155372
rect 14096 155252 14148 155304
rect 24860 155252 24912 155304
rect 31668 155252 31720 155304
rect 480 155184 532 155236
rect 1308 155184 1360 155236
rect 8208 155184 8260 155236
rect 125048 155184 125100 155236
rect 138020 155252 138072 155304
rect 136732 155184 136784 155236
rect 140780 155184 140832 155236
rect 141792 155252 141844 155304
rect 213920 155252 213972 155304
rect 262404 155252 262456 155304
rect 270316 155252 270368 155304
rect 270408 155252 270460 155304
rect 300124 155252 300176 155304
rect 306472 155388 306524 155440
rect 324228 155388 324280 155440
rect 327908 155388 327960 155440
rect 338488 155388 338540 155440
rect 409696 155388 409748 155440
rect 434168 155388 434220 155440
rect 436008 155388 436060 155440
rect 473176 155388 473228 155440
rect 483572 155388 483624 155440
rect 544292 155388 544344 155440
rect 549168 155388 549220 155440
rect 572628 155388 572680 155440
rect 307484 155320 307536 155372
rect 324136 155320 324188 155372
rect 325056 155320 325108 155372
rect 336648 155320 336700 155372
rect 401600 155320 401652 155372
rect 404912 155320 404964 155372
rect 411168 155320 411220 155372
rect 436100 155320 436152 155372
rect 438676 155320 438728 155372
rect 477040 155320 477092 155372
rect 491208 155320 491260 155372
rect 556068 155320 556120 155372
rect 302516 155252 302568 155304
rect 302608 155252 302660 155304
rect 321652 155252 321704 155304
rect 326988 155252 327040 155304
rect 338028 155252 338080 155304
rect 414572 155252 414624 155304
rect 440976 155252 441028 155304
rect 441252 155252 441304 155304
rect 480996 155252 481048 155304
rect 488356 155252 488408 155304
rect 552112 155252 552164 155304
rect 554780 155252 554832 155304
rect 569684 155252 569736 155304
rect 208400 155184 208452 155236
rect 209964 155184 210016 155236
rect 259828 155184 259880 155236
rect 260656 155184 260708 155236
rect 263600 155184 263652 155236
rect 287980 155184 288032 155236
rect 296720 155184 296772 155236
rect 29644 155116 29696 155168
rect 31668 155116 31720 155168
rect 55036 155116 55088 155168
rect 70400 155116 70452 155168
rect 90088 155116 90140 155168
rect 168380 155116 168432 155168
rect 169024 155116 169076 155168
rect 172428 155116 172480 155168
rect 172980 155116 173032 155168
rect 229192 155116 229244 155168
rect 239588 155116 239640 155168
rect 269396 155116 269448 155168
rect 274640 155116 274692 155168
rect 275284 155116 275336 155168
rect 51172 155048 51224 155100
rect 67364 155048 67416 155100
rect 83280 155048 83332 155100
rect 187700 155048 187752 155100
rect 188528 155048 188580 155100
rect 242992 155048 243044 155100
rect 62856 154980 62908 155032
rect 75000 154980 75052 155032
rect 101772 154980 101824 155032
rect 182088 154980 182140 155032
rect 185492 154980 185544 155032
rect 193128 154980 193180 155032
rect 237196 154980 237248 155032
rect 237288 154980 237340 155032
rect 273352 155048 273404 155100
rect 298008 155116 298060 155168
rect 298744 155184 298796 155236
rect 318984 155184 319036 155236
rect 323032 155184 323084 155236
rect 334072 155184 334124 155236
rect 338672 155184 338724 155236
rect 343640 155184 343692 155236
rect 382280 155184 382332 155236
rect 386420 155184 386472 155236
rect 401508 155184 401560 155236
rect 421564 155184 421616 155236
rect 422208 155184 422260 155236
rect 452752 155184 452804 155236
rect 454868 155184 454920 155236
rect 501420 155184 501472 155236
rect 503076 155184 503128 155236
rect 573548 155184 573600 155236
rect 301596 155116 301648 155168
rect 317328 155116 317380 155168
rect 318156 155116 318208 155168
rect 329748 155116 329800 155168
rect 332784 155116 332836 155168
rect 338580 155116 338632 155168
rect 343548 155116 343600 155168
rect 349068 155116 349120 155168
rect 398564 155116 398616 155168
rect 417608 155116 417660 155168
rect 419448 155116 419500 155168
rect 448796 155116 448848 155168
rect 467196 155116 467248 155168
rect 520004 155116 520056 155168
rect 282092 155048 282144 155100
rect 300676 155048 300728 155100
rect 309324 155048 309376 155100
rect 309416 155048 309468 155100
rect 323216 155048 323268 155100
rect 398932 155048 398984 155100
rect 401048 155048 401100 155100
rect 266360 154980 266412 155032
rect 269488 154980 269540 155032
rect 292580 154980 292632 155032
rect 294696 154980 294748 155032
rect 294788 154980 294840 155032
rect 316408 154980 316460 155032
rect 321100 154980 321152 155032
rect 332324 154980 332376 155032
rect 355232 154980 355284 155032
rect 356704 154980 356756 155032
rect 400956 154980 401008 155032
rect 420552 155048 420604 155100
rect 423036 155048 423088 155100
rect 453672 155048 453724 155100
rect 463608 155048 463660 155100
rect 515128 155048 515180 155100
rect 401692 154980 401744 155032
rect 403992 154980 404044 155032
rect 87144 154912 87196 154964
rect 197360 154912 197412 154964
rect 207112 154912 207164 154964
rect 256700 154912 256752 154964
rect 257804 154912 257856 154964
rect 269396 154912 269448 154964
rect 271696 154912 271748 154964
rect 272340 154912 272392 154964
rect 71596 154844 71648 154896
rect 144828 154844 144880 154896
rect 195980 154844 196032 154896
rect 202236 154844 202288 154896
rect 259368 154844 259420 154896
rect 106648 154776 106700 154828
rect 117412 154776 117464 154828
rect 185584 154776 185636 154828
rect 196348 154776 196400 154828
rect 245568 154776 245620 154828
rect 248972 154776 249024 154828
rect 98920 154708 98972 154760
rect 164884 154708 164936 154760
rect 165160 154708 165212 154760
rect 179512 154708 179564 154760
rect 179788 154708 179840 154760
rect 185676 154708 185728 154760
rect 189080 154708 189132 154760
rect 194416 154708 194468 154760
rect 86224 154640 86276 154692
rect 91008 154640 91060 154692
rect 96896 154640 96948 154692
rect 184296 154640 184348 154692
rect 184664 154640 184716 154692
rect 196532 154640 196584 154692
rect 198280 154708 198332 154760
rect 211068 154708 211120 154760
rect 211988 154708 212040 154760
rect 255320 154708 255372 154760
rect 256792 154708 256844 154760
rect 276756 154912 276808 154964
rect 277216 154912 277268 154964
rect 297916 154912 297968 154964
rect 299664 154912 299716 154964
rect 319628 154912 319680 154964
rect 322112 154912 322164 154964
rect 333888 154912 333940 154964
rect 357164 154912 357216 154964
rect 357992 154912 358044 154964
rect 365260 154912 365312 154964
rect 365996 154912 366048 154964
rect 400312 154912 400364 154964
rect 402980 154912 403032 154964
rect 285680 154844 285732 154896
rect 286048 154844 286100 154896
rect 307668 154844 307720 154896
rect 311348 154844 311400 154896
rect 321560 154844 321612 154896
rect 276020 154776 276072 154828
rect 276296 154776 276348 154828
rect 289268 154776 289320 154828
rect 293868 154776 293920 154828
rect 308588 154776 308640 154828
rect 310428 154776 310480 154828
rect 323032 154776 323084 154828
rect 324044 154776 324096 154828
rect 333980 154776 334032 154828
rect 341616 154776 341668 154828
rect 347504 154776 347556 154828
rect 384580 154776 384632 154828
rect 387432 154776 387484 154828
rect 400220 154776 400272 154828
rect 402060 154776 402112 154828
rect 418620 154980 418672 155032
rect 420460 154980 420512 155032
rect 449808 154980 449860 155032
rect 462044 154980 462096 155032
rect 512184 154980 512236 155032
rect 281172 154708 281224 154760
rect 295340 154708 295392 154760
rect 297732 154708 297784 154760
rect 314752 154708 314804 154760
rect 319168 154708 319220 154760
rect 205640 154640 205692 154692
rect 214288 154640 214340 154692
rect 223672 154640 223724 154692
rect 269028 154640 269080 154692
rect 283288 154640 283340 154692
rect 285036 154640 285088 154692
rect 1308 154572 1360 154624
rect 106188 154572 106240 154624
rect 110604 154572 110656 154624
rect 67732 154504 67784 154556
rect 164792 154504 164844 154556
rect 59912 154436 59964 154488
rect 48228 154368 48280 154420
rect 152004 154368 152056 154420
rect 158720 154436 158772 154488
rect 175280 154572 175332 154624
rect 183468 154572 183520 154624
rect 183652 154572 183704 154624
rect 191748 154572 191800 154624
rect 242256 154572 242308 154624
rect 246028 154572 246080 154624
rect 179420 154504 179472 154556
rect 184940 154504 184992 154556
rect 186320 154504 186372 154556
rect 201500 154504 201552 154556
rect 202788 154504 202840 154556
rect 249800 154504 249852 154556
rect 271788 154572 271840 154624
rect 288348 154572 288400 154624
rect 288992 154572 289044 154624
rect 159640 154368 159692 154420
rect 171968 154368 172020 154420
rect 175280 154368 175332 154420
rect 184296 154436 184348 154488
rect 198740 154436 198792 154488
rect 203156 154436 203208 154488
rect 255320 154436 255372 154488
rect 261116 154436 261168 154488
rect 266360 154436 266412 154488
rect 275376 154436 275428 154488
rect 281540 154504 281592 154556
rect 282920 154504 282972 154556
rect 298836 154504 298888 154556
rect 284024 154436 284076 154488
rect 285680 154436 285732 154488
rect 303528 154640 303580 154692
rect 303620 154640 303672 154692
rect 318708 154640 318760 154692
rect 320180 154640 320232 154692
rect 303804 154572 303856 154624
rect 304540 154572 304592 154624
rect 311164 154572 311216 154624
rect 312360 154572 312412 154624
rect 322940 154572 322992 154624
rect 193404 154368 193456 154420
rect 199292 154368 199344 154420
rect 252652 154368 252704 154420
rect 253848 154368 253900 154420
rect 289084 154368 289136 154420
rect 300860 154436 300912 154488
rect 301412 154368 301464 154420
rect 44272 154300 44324 154352
rect 149244 154300 149296 154352
rect 40408 154232 40460 154284
rect 146576 154232 146628 154284
rect 149060 154232 149112 154284
rect 164884 154300 164936 154352
rect 185676 154300 185728 154352
rect 186412 154300 186464 154352
rect 192484 154300 192536 154352
rect 247408 154300 247460 154352
rect 249984 154300 250036 154352
rect 254860 154300 254912 154352
rect 289820 154300 289872 154352
rect 292580 154300 292632 154352
rect 299480 154300 299532 154352
rect 340604 154708 340656 154760
rect 339684 154640 339736 154692
rect 346308 154640 346360 154692
rect 336740 154572 336792 154624
rect 332600 154504 332652 154556
rect 344376 154504 344428 154556
rect 399484 154708 399536 154760
rect 407028 154708 407080 154760
rect 417792 154912 417844 154964
rect 445852 154912 445904 154964
rect 464620 154912 464672 154964
rect 516048 154912 516100 154964
rect 352288 154640 352340 154692
rect 353392 154640 353444 154692
rect 406108 154640 406160 154692
rect 413836 154776 413888 154828
rect 415216 154708 415268 154760
rect 441988 154844 442040 154896
rect 463332 154844 463384 154896
rect 514116 154844 514168 154896
rect 417976 154776 418028 154828
rect 444932 154776 444984 154828
rect 459468 154776 459520 154828
rect 508228 154776 508280 154828
rect 438124 154708 438176 154760
rect 460112 154708 460164 154760
rect 509240 154708 509292 154760
rect 411996 154640 412048 154692
rect 437112 154640 437164 154692
rect 461400 154640 461452 154692
rect 511172 154640 511224 154692
rect 346492 154572 346544 154624
rect 347044 154504 347096 154556
rect 333244 154436 333296 154488
rect 340972 154436 341024 154488
rect 343732 154436 343784 154488
rect 309876 154300 309928 154352
rect 35532 154164 35584 154216
rect 143540 154164 143592 154216
rect 144736 154164 144788 154216
rect 161848 154164 161900 154216
rect 32588 154096 32640 154148
rect 141424 154096 141476 154148
rect 144828 154096 144880 154148
rect 167460 154232 167512 154284
rect 168380 154232 168432 154284
rect 179788 154232 179840 154284
rect 183376 154232 183428 154284
rect 240232 154232 240284 154284
rect 247040 154232 247092 154284
rect 284484 154232 284536 154284
rect 289268 154232 289320 154284
rect 303988 154232 304040 154284
rect 305000 154232 305052 154284
rect 315028 154232 315080 154284
rect 348424 154572 348476 154624
rect 349344 154572 349396 154624
rect 350356 154572 350408 154624
rect 351368 154572 351420 154624
rect 354128 154504 354180 154556
rect 361488 154504 361540 154556
rect 362040 154504 362092 154556
rect 362592 154504 362644 154556
rect 363052 154504 363104 154556
rect 365628 154504 365680 154556
rect 367928 154572 367980 154624
rect 366456 154504 366508 154556
rect 368848 154572 368900 154624
rect 353484 154436 353536 154488
rect 362868 154436 362920 154488
rect 363972 154436 364024 154488
rect 367008 154436 367060 154488
rect 369860 154436 369912 154488
rect 352840 154368 352892 154420
rect 367744 154368 367796 154420
rect 370872 154572 370924 154624
rect 374920 154504 374972 154556
rect 381544 154572 381596 154624
rect 372988 154436 373040 154488
rect 378600 154436 378652 154488
rect 375196 154368 375248 154420
rect 379704 154368 379756 154420
rect 352104 154300 352156 154352
rect 368388 154300 368440 154352
rect 371792 154300 371844 154352
rect 376208 154300 376260 154352
rect 383476 154572 383528 154624
rect 403992 154572 404044 154624
rect 405924 154572 405976 154624
rect 409420 154572 409472 154624
rect 433248 154572 433300 154624
rect 457536 154572 457588 154624
rect 505376 154572 505428 154624
rect 578424 154615 578476 154624
rect 578424 154581 578433 154615
rect 578433 154581 578467 154615
rect 578467 154581 578476 154615
rect 578424 154572 578476 154581
rect 382096 154504 382148 154556
rect 392308 154504 392360 154556
rect 395988 154504 396040 154556
rect 411260 154504 411312 154556
rect 415860 154504 415912 154556
rect 443000 154504 443052 154556
rect 471796 154504 471848 154556
rect 526812 154504 526864 154556
rect 384028 154436 384080 154488
rect 395160 154436 395212 154488
rect 395712 154436 395764 154488
rect 411352 154436 411404 154488
rect 416504 154436 416556 154488
rect 443920 154436 443972 154488
rect 500408 154436 500460 154488
rect 554780 154436 554832 154488
rect 384672 154368 384724 154420
rect 396172 154368 396224 154420
rect 397000 154368 397052 154420
rect 413284 154368 413336 154420
rect 419172 154368 419224 154420
rect 447876 154368 447928 154420
rect 482192 154368 482244 154420
rect 542268 154368 542320 154420
rect 385960 154300 386012 154352
rect 398104 154300 398156 154352
rect 398288 154300 398340 154352
rect 414112 154300 414164 154352
rect 421748 154300 421800 154352
rect 451740 154300 451792 154352
rect 486148 154300 486200 154352
rect 546500 154300 546552 154352
rect 548524 154300 548576 154352
rect 575572 154300 575624 154352
rect 350816 154232 350868 154284
rect 369676 154232 369728 154284
rect 373724 154232 373776 154284
rect 384948 154232 385000 154284
rect 397184 154232 397236 154284
rect 397276 154232 397328 154284
rect 415676 154232 415728 154284
rect 424324 154232 424376 154284
rect 455604 154232 455656 154284
rect 487068 154232 487120 154284
rect 550180 154232 550232 154284
rect 162124 154164 162176 154216
rect 178040 154164 178092 154216
rect 179144 154164 179196 154216
rect 237656 154164 237708 154216
rect 241428 154164 241480 154216
rect 279332 154164 279384 154216
rect 285680 154164 285732 154216
rect 290832 154164 290884 154216
rect 306656 154164 306708 154216
rect 308404 154164 308456 154216
rect 317696 154164 317748 154216
rect 347596 154164 347648 154216
rect 350172 154164 350224 154216
rect 372344 154164 372396 154216
rect 377680 154164 377732 154216
rect 386236 154164 386288 154216
rect 398748 154164 398800 154216
rect 400128 154164 400180 154216
rect 419540 154164 419592 154216
rect 426900 154164 426952 154216
rect 459560 154164 459612 154216
rect 489644 154164 489696 154216
rect 554044 154164 554096 154216
rect 167000 154096 167052 154148
rect 172428 154096 172480 154148
rect 232504 154096 232556 154148
rect 235356 154096 235408 154148
rect 28724 154028 28776 154080
rect 138848 154028 138900 154080
rect 140780 154028 140832 154080
rect 156972 154028 157024 154080
rect 157340 154028 157392 154080
rect 224960 154028 225012 154080
rect 233148 154028 233200 154080
rect 273444 154028 273496 154080
rect 276020 154096 276072 154148
rect 285772 154096 285824 154148
rect 291752 154096 291804 154148
rect 309232 154096 309284 154148
rect 309324 154096 309376 154148
rect 320272 154096 320324 154148
rect 381452 154096 381504 154148
rect 387340 154096 387392 154148
rect 390468 154096 390520 154148
rect 401600 154096 401652 154148
rect 403532 154096 403584 154148
rect 424416 154096 424468 154148
rect 429568 154096 429620 154148
rect 463424 154096 463476 154148
rect 474464 154096 474516 154148
rect 480076 154096 480128 154148
rect 492588 154096 492640 154148
rect 558000 154096 558052 154148
rect 276664 154028 276716 154080
rect 276756 154028 276808 154080
rect 291200 154028 291252 154080
rect 291844 154028 291896 154080
rect 314660 154028 314712 154080
rect 387708 154028 387760 154080
rect 398932 154028 398984 154080
rect 402704 154028 402756 154080
rect 423496 154028 423548 154080
rect 431776 154028 431828 154080
rect 467288 154028 467340 154080
rect 495256 154028 495308 154080
rect 561588 154028 561640 154080
rect 20904 153960 20956 154012
rect 133880 153960 133932 154012
rect 135168 153960 135220 154012
rect 138020 153960 138072 154012
rect 145932 153960 145984 154012
rect 153108 153960 153160 154012
rect 219624 153960 219676 154012
rect 227536 153960 227588 154012
rect 271512 153960 271564 154012
rect 274640 153960 274692 154012
rect 288440 153960 288492 154012
rect 289912 153960 289964 154012
rect 313280 153960 313332 154012
rect 369032 153960 369084 154012
rect 372804 153960 372856 154012
rect 373908 153960 373960 154012
rect 378140 153960 378192 154012
rect 388536 153960 388588 154012
rect 400220 153960 400272 154012
rect 405464 153960 405516 154012
rect 427360 153960 427412 154012
rect 432788 153960 432840 154012
rect 468300 153960 468352 154012
rect 497832 153960 497884 154012
rect 565728 153960 565780 154012
rect 13084 153892 13136 153944
rect 128360 153892 128412 153944
rect 9220 153824 9272 153876
rect 125784 153824 125836 153876
rect 126060 153824 126112 153876
rect 135536 153892 135588 153944
rect 136732 153892 136784 153944
rect 140780 153892 140832 153944
rect 140872 153892 140924 153944
rect 144000 153892 144052 153944
rect 145656 153892 145708 153944
rect 216864 153892 216916 153944
rect 222108 153892 222160 153944
rect 266360 153892 266412 153944
rect 266452 153892 266504 153944
rect 296996 153892 297048 153944
rect 300860 153892 300912 153944
rect 312452 153892 312504 153944
rect 328460 153892 328512 153944
rect 330668 153892 330720 153944
rect 334348 153892 334400 153944
rect 339132 153892 339184 153944
rect 340236 153892 340288 153944
rect 342996 153892 343048 153944
rect 377496 153892 377548 153944
rect 382372 153892 382424 153944
rect 383292 153892 383344 153944
rect 394240 153892 394292 153944
rect 394424 153892 394476 153944
rect 410800 153892 410852 153944
rect 435364 153892 435416 153944
rect 472164 153892 472216 153944
rect 499120 153892 499172 153944
rect 567752 153892 567804 153944
rect 130108 153824 130160 153876
rect 206468 153824 206520 153876
rect 208032 153824 208084 153876
rect 258448 153824 258500 153876
rect 262128 153824 262180 153876
rect 292580 153824 292632 153876
rect 295340 153824 295392 153876
rect 307300 153824 307352 153876
rect 311164 153824 311216 153876
rect 323124 153824 323176 153876
rect 373632 153824 373684 153876
rect 379428 153824 379480 153876
rect 391204 153824 391256 153876
rect 403992 153824 404044 153876
rect 408040 153824 408092 153876
rect 431224 153824 431276 153876
rect 434628 153824 434680 153876
rect 471244 153824 471296 153876
rect 479616 153824 479668 153876
rect 487160 153824 487212 153876
rect 501696 153824 501748 153876
rect 571248 153824 571300 153876
rect 78404 153756 78456 153808
rect 79416 153688 79468 153740
rect 172612 153756 172664 153808
rect 179512 153756 179564 153808
rect 167736 153688 167788 153740
rect 169392 153688 169444 153740
rect 94964 153620 95016 153672
rect 183008 153688 183060 153740
rect 187700 153756 187752 153808
rect 216220 153756 216272 153808
rect 216588 153756 216640 153808
rect 263692 153756 263744 153808
rect 271788 153756 271840 153808
rect 283196 153756 283248 153808
rect 283288 153756 283340 153808
rect 296168 153756 296220 153808
rect 305276 153756 305328 153808
rect 337936 153756 337988 153808
rect 341064 153756 341116 153808
rect 347780 153756 347832 153808
rect 351460 153756 351512 153808
rect 382740 153756 382792 153808
rect 388444 153756 388496 153808
rect 395068 153756 395120 153808
rect 411812 153756 411864 153808
rect 418528 153756 418580 153808
rect 446864 153756 446916 153808
rect 470324 153756 470376 153808
rect 524880 153756 524932 153808
rect 185584 153688 185636 153740
rect 197360 153688 197412 153740
rect 222200 153688 222252 153740
rect 233240 153688 233292 153740
rect 270868 153688 270920 153740
rect 271972 153688 272024 153740
rect 274088 153688 274140 153740
rect 279148 153688 279200 153740
rect 293592 153688 293644 153740
rect 335636 153688 335688 153740
rect 339776 153688 339828 153740
rect 393044 153688 393096 153740
rect 408868 153688 408920 153740
rect 413284 153688 413336 153740
rect 439044 153688 439096 153740
rect 467748 153688 467800 153740
rect 520924 153688 520976 153740
rect 187700 153620 187752 153672
rect 211160 153620 211212 153672
rect 237380 153620 237432 153672
rect 242900 153620 242952 153672
rect 248052 153620 248104 153672
rect 255320 153620 255372 153672
rect 262220 153620 262272 153672
rect 264980 153620 265032 153672
rect 280620 153620 280672 153672
rect 281540 153620 281592 153672
rect 291660 153620 291712 153672
rect 292764 153620 292816 153672
rect 294236 153620 294288 153672
rect 324136 153620 324188 153672
rect 324872 153620 324924 153672
rect 338948 153620 339000 153672
rect 342352 153620 342404 153672
rect 376484 153620 376536 153672
rect 380900 153620 380952 153672
rect 389088 153620 389140 153672
rect 400312 153620 400364 153672
rect 413928 153620 413980 153672
rect 440056 153620 440108 153672
rect 464988 153620 465040 153672
rect 517060 153620 517112 153672
rect 93032 153552 93084 153604
rect 181720 153552 181772 153604
rect 182088 153552 182140 153604
rect 190828 153552 190880 153604
rect 198004 153552 198056 153604
rect 253296 153552 253348 153604
rect 100852 153484 100904 153536
rect 186964 153484 187016 153536
rect 195980 153484 196032 153536
rect 211620 153484 211672 153536
rect 229192 153484 229244 153536
rect 235080 153484 235132 153536
rect 251180 153484 251232 153536
rect 255872 153552 255924 153604
rect 265072 153552 265124 153604
rect 270500 153552 270552 153604
rect 280252 153552 280304 153604
rect 281908 153552 281960 153604
rect 284392 153552 284444 153604
rect 286416 153552 286468 153604
rect 288348 153552 288400 153604
rect 297548 153552 297600 153604
rect 322940 153552 322992 153604
rect 328092 153552 328144 153604
rect 380072 153552 380124 153604
rect 386328 153552 386380 153604
rect 389824 153552 389876 153604
rect 401692 153552 401744 153604
rect 410708 153552 410760 153604
rect 435180 153552 435232 153604
rect 458088 153552 458140 153604
rect 506296 153552 506348 153604
rect 270316 153484 270368 153536
rect 272800 153484 272852 153536
rect 298008 153484 298060 153536
rect 302240 153484 302292 153536
rect 317328 153484 317380 153536
rect 320916 153484 320968 153536
rect 321560 153484 321612 153536
rect 327448 153484 327500 153536
rect 329748 153484 329800 153536
rect 331956 153484 332008 153536
rect 333980 153484 334032 153536
rect 335912 153484 335964 153536
rect 338580 153484 338632 153536
rect 341708 153484 341760 153536
rect 370964 153484 371016 153536
rect 375748 153484 375800 153536
rect 378784 153484 378836 153536
rect 384580 153484 384632 153536
rect 393780 153484 393832 153536
rect 405832 153484 405884 153536
rect 477040 153484 477092 153536
rect 482744 153484 482796 153536
rect 502248 153484 502300 153536
rect 549168 153484 549220 153536
rect 102784 153416 102836 153468
rect 188252 153416 188304 153468
rect 193128 153416 193180 153468
rect 203156 153416 203208 153468
rect 242992 153416 243044 153468
rect 245660 153416 245712 153468
rect 277400 153416 277452 153468
rect 278780 153416 278832 153468
rect 323032 153416 323084 153468
rect 327080 153416 327132 153468
rect 333888 153416 333940 153468
rect 334624 153416 334676 153468
rect 365168 153416 365220 153468
rect 366916 153416 366968 153468
rect 370320 153416 370372 153468
rect 374736 153416 374788 153468
rect 378048 153416 378100 153468
rect 382280 153416 382332 153468
rect 392492 153416 392544 153468
rect 404636 153416 404688 153468
rect 455236 153416 455288 153468
rect 502156 153416 502208 153468
rect 109592 153348 109644 153400
rect 112444 153280 112496 153332
rect 114468 153348 114520 153400
rect 196072 153348 196124 153400
rect 259368 153348 259420 153400
rect 260472 153348 260524 153400
rect 297916 153348 297968 153400
rect 304632 153348 304684 153400
rect 307668 153348 307720 153400
rect 310520 153348 310572 153400
rect 323216 153348 323268 153400
rect 326160 153348 326212 153400
rect 332324 153348 332376 153400
rect 333980 153348 334032 153400
rect 336556 153348 336608 153400
rect 340420 153348 340472 153400
rect 342536 153348 342588 153400
rect 345204 153348 345256 153400
rect 379428 153348 379480 153400
rect 384764 153348 384816 153400
rect 391848 153348 391900 153400
rect 404176 153348 404228 153400
rect 456248 153348 456300 153400
rect 503352 153348 503404 153400
rect 12808 153212 12860 153264
rect 26700 153212 26752 153264
rect 46756 153212 46808 153264
rect 92204 153212 92256 153264
rect 108948 153212 109000 153264
rect 112536 153212 112588 153264
rect 192760 153280 192812 153332
rect 245568 153280 245620 153332
rect 250720 153280 250772 153332
rect 263784 153280 263836 153332
rect 268200 153280 268252 153332
rect 271696 153280 271748 153332
rect 277952 153280 278004 153332
rect 303804 153280 303856 153332
rect 307944 153280 307996 153332
rect 314752 153280 314804 153332
rect 318340 153280 318392 153332
rect 343640 153280 343692 153332
rect 345664 153280 345716 153332
rect 364156 153280 364208 153332
rect 365260 153280 365312 153332
rect 371608 153280 371660 153332
rect 376668 153280 376720 153332
rect 387248 153280 387300 153332
rect 400036 153280 400088 153332
rect 417148 153280 417200 153332
rect 417976 153280 418028 153332
rect 514668 153280 514720 153332
rect 520556 153280 520608 153332
rect 117780 153212 117832 153264
rect 117964 153212 118016 153264
rect 130384 153212 130436 153264
rect 132960 153212 133012 153264
rect 133788 153212 133840 153264
rect 138112 153212 138164 153264
rect 184296 153212 184348 153264
rect 189080 153212 189132 153264
rect 203892 153212 203944 153264
rect 225052 153212 225104 153264
rect 229836 153212 229888 153264
rect 249800 153212 249852 153264
rect 254584 153212 254636 153264
rect 256700 153212 256752 153264
rect 258080 153212 258132 153264
rect 285680 153212 285732 153264
rect 287244 153212 287296 153264
rect 313372 153212 313424 153264
rect 316040 153212 316092 153264
rect 318708 153212 318760 153264
rect 322204 153212 322256 153264
rect 324412 153212 324464 153264
rect 325792 153212 325844 153264
rect 334072 153212 334124 153264
rect 335452 153212 335504 153264
rect 353392 153212 353444 153264
rect 354864 153212 354916 153264
rect 363880 153212 363932 153264
rect 364984 153212 365036 153264
rect 380716 153212 380768 153264
rect 385500 153212 385552 153264
rect 412456 153212 412508 153264
rect 413836 153212 413888 153264
rect 473084 153212 473136 153264
rect 476120 153212 476172 153264
rect 516048 153212 516100 153264
rect 520648 153212 520700 153264
rect 72608 153144 72660 153196
rect 168380 153144 168432 153196
rect 170036 153144 170088 153196
rect 233240 153144 233292 153196
rect 468576 153144 468628 153196
rect 521936 153144 521988 153196
rect 60832 153076 60884 153128
rect 160284 153076 160336 153128
rect 162308 153076 162360 153128
rect 54024 153008 54076 153060
rect 155960 153008 156012 153060
rect 156420 153008 156472 153060
rect 168104 153076 168156 153128
rect 231860 153076 231912 153128
rect 431500 153076 431552 153128
rect 466368 153076 466420 153128
rect 472440 153076 472492 153128
rect 527732 153076 527784 153128
rect 49148 152940 49200 152992
rect 152464 152940 152516 152992
rect 24860 152872 24912 152924
rect 129004 152872 129056 152924
rect 142712 152872 142764 152924
rect 149152 152872 149204 152924
rect 227904 153008 227956 153060
rect 259736 153008 259788 153060
rect 292948 153008 293000 153060
rect 434076 153008 434128 153060
rect 470232 153008 470284 153060
rect 476028 153008 476080 153060
rect 533620 153008 533672 153060
rect 215576 152940 215628 152992
rect 255780 152940 255832 152992
rect 290372 152940 290424 152992
rect 439964 152940 440016 152992
rect 479064 152940 479116 152992
rect 480076 152940 480128 152992
rect 539508 152940 539560 152992
rect 224040 152872 224092 152924
rect 248144 152872 248196 152924
rect 285128 152872 285180 152924
rect 441712 152872 441764 152924
rect 481916 152872 481968 152924
rect 484216 152872 484268 152924
rect 545304 152872 545356 152924
rect 45284 152804 45336 152856
rect 149888 152804 149940 152856
rect 154488 152804 154540 152856
rect 222752 152804 222804 152856
rect 240324 152804 240376 152856
rect 280160 152804 280212 152856
rect 444288 152804 444340 152856
rect 485872 152804 485924 152856
rect 488080 152804 488132 152856
rect 551192 152804 551244 152856
rect 46204 152736 46256 152788
rect 150532 152736 150584 152788
rect 151544 152736 151596 152788
rect 220820 152736 220872 152788
rect 232412 152736 232464 152788
rect 274732 152736 274784 152788
rect 447048 152736 447100 152788
rect 489276 152736 489328 152788
rect 489368 152736 489420 152788
rect 553124 152736 553176 152788
rect 41328 152668 41380 152720
rect 147220 152668 147272 152720
rect 31668 152600 31720 152652
rect 139492 152600 139544 152652
rect 146668 152600 146720 152652
rect 217508 152668 217560 152720
rect 224592 152668 224644 152720
rect 269580 152668 269632 152720
rect 448428 152668 448480 152720
rect 491668 152668 491720 152720
rect 491944 152668 491996 152720
rect 556988 152668 557040 152720
rect 214932 152600 214984 152652
rect 220728 152600 220780 152652
rect 266912 152600 266964 152652
rect 451648 152600 451700 152652
rect 21916 152532 21968 152584
rect 134248 152532 134300 152584
rect 138940 152532 138992 152584
rect 212540 152532 212592 152584
rect 216956 152532 217008 152584
rect 264336 152532 264388 152584
rect 450912 152532 450964 152584
rect 495624 152532 495676 152584
rect 495900 152600 495952 152652
rect 562876 152600 562928 152652
rect 496452 152532 496504 152584
rect 498108 152532 498160 152584
rect 566740 152532 566792 152584
rect 7288 152464 7340 152516
rect 124496 152464 124548 152516
rect 135904 152464 135956 152516
rect 210332 152464 210384 152516
rect 214840 152464 214892 152516
rect 263048 152464 263100 152516
rect 271420 152464 271472 152516
rect 300860 152464 300912 152516
rect 423588 152464 423640 152516
rect 454684 152464 454736 152516
rect 458824 152464 458876 152516
rect 507308 152464 507360 152516
rect 510160 152464 510212 152516
rect 61844 152396 61896 152448
rect 160928 152396 160980 152448
rect 165528 152396 165580 152448
rect 228548 152396 228600 152448
rect 439320 152396 439372 152448
rect 478052 152396 478104 152448
rect 482744 152396 482796 152448
rect 534632 152396 534684 152448
rect 69664 152328 69716 152380
rect 166080 152328 166132 152380
rect 172520 152328 172572 152380
rect 233792 152328 233844 152380
rect 476120 152328 476172 152380
rect 528744 152328 528796 152380
rect 77484 152260 77536 152312
rect 171416 152260 171468 152312
rect 181812 152260 181864 152312
rect 240968 152260 241020 152312
rect 462688 152260 462740 152312
rect 513104 152260 513156 152312
rect 80336 152192 80388 152244
rect 173578 152192 173630 152244
rect 185768 152192 185820 152244
rect 243866 152192 243918 152244
rect 453902 152192 453954 152244
rect 500500 152192 500552 152244
rect 85212 152124 85264 152176
rect 176890 152124 176942 152176
rect 187608 152124 187660 152176
rect 245154 152124 245206 152176
rect 452614 152124 452666 152176
rect 498568 152124 498620 152176
rect 88156 152056 88208 152108
rect 178822 152056 178874 152108
rect 187792 152056 187844 152108
rect 95976 151988 96028 152040
rect 183652 151988 183704 152040
rect 43812 151963 43864 151972
rect 43812 151929 43821 151963
rect 43821 151929 43855 151963
rect 43855 151929 43864 151963
rect 43812 151920 43864 151929
rect 57520 151963 57572 151972
rect 57520 151929 57529 151963
rect 57529 151929 57563 151963
rect 57563 151929 57572 151963
rect 57520 151920 57572 151929
rect 60832 151963 60884 151972
rect 60832 151929 60841 151963
rect 60841 151929 60875 151963
rect 60875 151929 60884 151963
rect 60832 151920 60884 151929
rect 64420 151963 64472 151972
rect 64420 151929 64429 151963
rect 64429 151929 64463 151963
rect 64463 151929 64472 151963
rect 64420 151920 64472 151929
rect 67364 151963 67416 151972
rect 67364 151929 67373 151963
rect 67373 151929 67407 151963
rect 67407 151929 67416 151963
rect 67364 151920 67416 151929
rect 74540 151963 74592 151972
rect 74540 151929 74549 151963
rect 74549 151929 74583 151963
rect 74583 151929 74592 151963
rect 74540 151920 74592 151929
rect 78128 151963 78180 151972
rect 78128 151929 78137 151963
rect 78137 151929 78171 151963
rect 78171 151929 78180 151963
rect 78128 151920 78180 151929
rect 85028 151963 85080 151972
rect 85028 151929 85037 151963
rect 85037 151929 85071 151963
rect 85071 151929 85080 151963
rect 85028 151920 85080 151929
rect 91008 151963 91060 151972
rect 91008 151929 91017 151963
rect 91017 151929 91051 151963
rect 91051 151929 91060 151963
rect 91008 151920 91060 151929
rect 95148 151963 95200 151972
rect 95148 151929 95157 151963
rect 95157 151929 95191 151963
rect 95191 151929 95200 151963
rect 95148 151920 95200 151929
rect 105636 151963 105688 151972
rect 105636 151929 105645 151963
rect 105645 151929 105679 151963
rect 105679 151929 105688 151963
rect 105636 151920 105688 151929
rect 115480 151920 115532 151972
rect 197038 152056 197090 152108
rect 201224 152056 201276 152108
rect 254262 152056 254314 152108
rect 449394 152056 449446 152108
rect 493692 152056 493744 152108
rect 3240 151852 3292 151904
rect 115112 151852 115164 151904
rect 120448 151852 120500 151904
rect 200120 151988 200172 152040
rect 205088 151988 205140 152040
rect 256700 151988 256752 152040
rect 443828 151988 443880 152040
rect 484952 151988 485004 152040
rect 238944 151920 238996 151972
rect 196532 151852 196584 151904
rect 246948 151852 247000 151904
rect 503628 151852 503680 151904
rect 520280 151852 520332 151904
rect 3516 151784 3568 151836
rect 117044 151784 117096 151836
rect 127532 151784 127584 151836
rect 204536 151784 204588 151836
rect 211068 151784 211120 151836
rect 252008 151784 252060 151836
rect 505008 151784 505060 151836
rect 525064 151784 525116 151836
rect 2964 151716 3016 151768
rect 114192 151716 114244 151768
rect 3148 151648 3200 151700
rect 115664 151648 115716 151700
rect 3240 151580 3292 151632
rect 112904 151580 112956 151632
rect 16304 151555 16356 151564
rect 16304 151521 16313 151555
rect 16313 151521 16347 151555
rect 16347 151521 16356 151555
rect 16304 151512 16356 151521
rect 26700 151512 26752 151564
rect 118608 151512 118660 151564
rect 5080 151444 5132 151496
rect 112812 151444 112864 151496
rect 3792 151376 3844 151428
rect 112536 151376 112588 151428
rect 177212 151419 177264 151428
rect 177212 151385 177221 151419
rect 177221 151385 177255 151419
rect 177255 151385 177264 151419
rect 177212 151376 177264 151385
rect 3608 151308 3660 151360
rect 112996 151308 113048 151360
rect 116952 151308 117004 151360
rect 507768 151512 507820 151564
rect 505652 151444 505704 151496
rect 118056 151172 118108 151224
rect 119712 151172 119764 151224
rect 506940 151376 506992 151428
rect 503720 151308 503772 151360
rect 113916 151104 113968 151156
rect 114284 151036 114336 151088
rect 119436 151036 119488 151088
rect 510160 151308 510212 151360
rect 513288 151444 513340 151496
rect 520740 151444 520792 151496
rect 517980 151376 518032 151428
rect 520372 151376 520424 151428
rect 519268 151308 519320 151360
rect 520464 151308 520516 151360
rect 527824 151104 527876 151156
rect 117136 150968 117188 151020
rect 519728 150900 519780 150952
rect 522120 150832 522172 150884
rect 522212 150764 522264 150816
rect 520832 150696 520884 150748
rect 521936 150628 521988 150680
rect 521752 150560 521804 150612
rect 116860 150492 116912 150544
rect 4068 150424 4120 150476
rect 5540 150424 5592 150476
rect 117780 150424 117832 150476
rect 3700 150356 3752 150408
rect 112444 150356 112496 150408
rect 3884 150288 3936 150340
rect 114100 150288 114152 150340
rect 3976 150220 4028 150272
rect 118424 150220 118476 150272
rect 112904 149336 112956 149388
rect 114008 149336 114060 149388
rect 3424 149064 3476 149116
rect 5080 149064 5132 149116
rect 115296 147636 115348 147688
rect 117688 147636 117740 147688
rect 3240 146684 3292 146736
rect 3424 146684 3476 146736
rect 112628 146208 112680 146260
rect 117320 146208 117372 146260
rect 115388 142536 115440 142588
rect 117320 142536 117372 142588
rect 115480 140768 115532 140820
rect 117320 140768 117372 140820
rect 115572 137980 115624 138032
rect 117688 137980 117740 138032
rect 115112 133832 115164 133884
rect 117872 133832 117924 133884
rect 114284 133764 114336 133816
rect 117320 133764 117372 133816
rect 116492 115948 116544 116000
rect 117504 115948 117556 116000
rect 112720 113976 112772 114028
rect 115848 113976 115900 114028
rect 112628 94324 112680 94376
rect 115112 94324 115164 94376
rect 115756 88272 115808 88324
rect 117688 88272 117740 88324
rect 115848 81812 115900 81864
rect 117872 81812 117924 81864
rect 114192 81336 114244 81388
rect 117320 81336 117372 81388
rect 115112 79296 115164 79348
rect 117780 79296 117832 79348
rect 115664 78616 115716 78668
rect 117688 78616 117740 78668
rect 112536 74536 112588 74588
rect 114560 74536 114612 74588
rect 114100 71680 114152 71732
rect 117320 71680 117372 71732
rect 114560 68960 114612 69012
rect 117320 68960 117372 69012
rect 116400 67532 116452 67584
rect 119436 67532 119488 67584
rect 112444 66172 112496 66224
rect 117320 66172 117372 66224
rect 114008 61616 114060 61668
rect 117320 61616 117372 61668
rect 2780 56856 2832 56908
rect 4804 56856 4856 56908
rect 114008 55564 114060 55616
rect 117320 55564 117372 55616
rect 115664 52436 115716 52488
rect 117320 52436 117372 52488
rect 114100 48220 114152 48272
rect 117320 48288 117372 48340
rect 115756 46112 115808 46164
rect 117228 46112 117280 46164
rect 114192 44072 114244 44124
rect 117872 44140 117924 44192
rect 3792 39992 3844 40044
rect 4896 39992 4948 40044
rect 114284 39992 114336 40044
rect 117320 40060 117372 40112
rect 112536 38632 112588 38684
rect 117320 38632 117372 38684
rect 114560 37000 114612 37052
rect 117228 37000 117280 37052
rect 114652 36184 114704 36236
rect 117320 36184 117372 36236
rect 522580 34416 522632 34468
rect 548524 34416 548576 34468
rect 113732 31764 113784 31816
rect 117320 31764 117372 31816
rect 3700 30268 3752 30320
rect 4988 30268 5040 30320
rect 113640 28976 113692 29028
rect 117320 28976 117372 29028
rect 112628 27616 112680 27668
rect 114468 27616 114520 27668
rect 113732 27480 113784 27532
rect 114468 27480 114520 27532
rect 3608 24828 3660 24880
rect 5080 24828 5132 24880
rect 3884 21360 3936 21412
rect 5172 21360 5224 21412
rect 3332 17892 3384 17944
rect 5264 17892 5316 17944
rect 115848 16872 115900 16924
rect 117504 16872 117556 16924
rect 522672 15104 522724 15156
rect 573364 15104 573416 15156
rect 113640 13812 113692 13864
rect 117320 13812 117372 13864
rect 3240 13540 3292 13592
rect 5448 13540 5500 13592
rect 521660 12928 521712 12980
rect 521844 12928 521896 12980
rect 3976 12860 4028 12912
rect 5356 12860 5408 12912
rect 117688 11704 117740 11756
rect 117964 11704 118016 11756
rect 115112 9664 115164 9716
rect 117320 9664 117372 9716
rect 3332 8916 3384 8968
rect 3608 8916 3660 8968
rect 3608 8780 3660 8832
rect 4068 8780 4120 8832
rect 116032 8304 116084 8356
rect 118976 8304 119028 8356
rect 114560 7148 114612 7200
rect 117320 7148 117372 7200
rect 112444 5924 112496 5976
rect 112720 5924 112772 5976
rect 2964 5856 3016 5908
rect 118516 5856 118568 5908
rect 2872 5788 2924 5840
rect 117872 5788 117924 5840
rect 2780 5720 2832 5772
rect 117136 5720 117188 5772
rect 3792 5652 3844 5704
rect 117780 5652 117832 5704
rect 3148 5584 3200 5636
rect 114468 5584 114520 5636
rect 3056 5516 3108 5568
rect 113732 5516 113784 5568
rect 3976 5448 4028 5500
rect 117228 5448 117280 5500
rect 3424 5380 3476 5432
rect 3700 5312 3752 5364
rect 112444 5380 112496 5432
rect 112628 5380 112680 5432
rect 115296 5380 115348 5432
rect 115664 5312 115716 5364
rect 116584 5312 116636 5364
rect 116952 5312 117004 5364
rect 3240 5244 3292 5296
rect 114560 5244 114612 5296
rect 4068 5176 4120 5228
rect 115112 5176 115164 5228
rect 3516 5108 3568 5160
rect 114376 5108 114428 5160
rect 116676 5108 116728 5160
rect 571984 5108 572036 5160
rect 4988 5040 5040 5092
rect 114008 5040 114060 5092
rect 118884 5040 118936 5092
rect 521752 4972 521804 5024
rect 3332 4904 3384 4956
rect 113640 4904 113692 4956
rect 118700 4904 118752 4956
rect 566556 4904 566608 4956
rect 520832 4836 520884 4888
rect 4896 4768 4948 4820
rect 115848 4768 115900 4820
rect 118792 4768 118844 4820
rect 577228 4768 577280 4820
rect 5080 4700 5132 4752
rect 114100 4700 114152 4752
rect 5172 4632 5224 4684
rect 114192 4632 114244 4684
rect 168840 4675 168892 4684
rect 168840 4641 168849 4675
rect 168849 4641 168883 4675
rect 168883 4641 168892 4675
rect 168840 4632 168892 4641
rect 474464 4675 474516 4684
rect 474464 4641 474473 4675
rect 474473 4641 474507 4675
rect 474507 4641 474516 4675
rect 474464 4632 474516 4641
rect 518624 4675 518676 4684
rect 518624 4641 518633 4675
rect 518633 4641 518667 4675
rect 518667 4641 518676 4675
rect 518624 4632 518676 4641
rect 519636 4632 519688 4684
rect 522396 4632 522448 4684
rect 5356 4564 5408 4616
rect 114284 4564 114336 4616
rect 5264 4496 5316 4548
rect 5448 4428 5500 4480
rect 115756 4496 115808 4548
rect 112720 4428 112772 4480
rect 42616 4360 42668 4412
rect 118332 4360 118384 4412
rect 62672 4292 62724 4344
rect 116768 4292 116820 4344
rect 65984 4267 66036 4276
rect 65984 4233 65993 4267
rect 65993 4233 66027 4267
rect 66027 4233 66036 4267
rect 65984 4224 66036 4233
rect 66168 4224 66220 4276
rect 118056 4224 118108 4276
rect 2964 4156 3016 4208
rect 117320 4156 117372 4208
rect 520096 4156 520148 4208
rect 522120 4156 522172 4208
rect 7840 4088 7892 4140
rect 124680 4088 124732 4140
rect 125140 4088 125192 4140
rect 45100 4020 45152 4072
rect 116860 4020 116912 4072
rect 117044 4020 117096 4072
rect 86868 3995 86920 4004
rect 86868 3961 86877 3995
rect 86877 3961 86911 3995
rect 86911 3961 86920 3995
rect 86868 3952 86920 3961
rect 114284 3952 114336 4004
rect 130292 4088 130344 4140
rect 198740 4088 198792 4140
rect 404268 4088 404320 4140
rect 454316 4088 454368 4140
rect 527824 4088 527876 4140
rect 529296 4088 529348 4140
rect 195244 4020 195296 4072
rect 215392 4020 215444 4072
rect 252560 4020 252612 4072
rect 407672 4020 407724 4072
rect 460112 4020 460164 4072
rect 461492 4020 461544 4072
rect 545304 4020 545356 4072
rect 470876 3952 470928 4004
rect 77024 3884 77076 3936
rect 164976 3884 165028 3936
rect 82360 3816 82412 3868
rect 66444 3748 66496 3800
rect 158260 3748 158312 3800
rect 162216 3748 162268 3800
rect 219118 3884 219170 3936
rect 311164 3884 311216 3936
rect 313234 3884 313286 3936
rect 414066 3884 414118 3936
rect 470784 3884 470836 3936
rect 168288 3816 168340 3868
rect 178132 3816 178184 3868
rect 229100 3816 229152 3868
rect 417792 3816 417844 3868
rect 476120 3816 476172 3868
rect 167460 3748 167512 3800
rect 222200 3748 222252 3800
rect 420736 3748 420788 3800
rect 481456 3748 481508 3800
rect 61108 3680 61160 3732
rect 154948 3680 155000 3732
rect 55772 3612 55824 3664
rect 146944 3612 146996 3664
rect 151544 3612 151596 3664
rect 212080 3680 212132 3732
rect 241980 3680 242032 3732
rect 269212 3680 269264 3732
rect 411076 3680 411128 3732
rect 465448 3680 465500 3732
rect 208676 3612 208728 3664
rect 226064 3612 226116 3664
rect 259460 3612 259512 3664
rect 367008 3612 367060 3664
rect 396264 3612 396316 3664
rect 401600 3612 401652 3664
rect 424508 3612 424560 3664
rect 486700 3612 486752 3664
rect 50436 3544 50488 3596
rect 141608 3544 141660 3596
rect 39764 3476 39816 3528
rect 108856 3476 108908 3528
rect 113916 3476 113968 3528
rect 114652 3476 114704 3528
rect 118240 3476 118292 3528
rect 118976 3476 119028 3528
rect 128360 3476 128412 3528
rect 140872 3476 140924 3528
rect 205640 3544 205692 3596
rect 373908 3544 373960 3596
rect 406936 3544 406988 3596
rect 427728 3544 427780 3596
rect 492036 3544 492088 3596
rect 508044 3544 508096 3596
rect 520280 3544 520332 3596
rect 201960 3476 202012 3528
rect 213828 3476 213880 3528
rect 521844 3476 521896 3528
rect 98368 3408 98420 3460
rect 178500 3408 178552 3460
rect 93032 3340 93084 3392
rect 175280 3340 175332 3392
rect 176660 3340 176712 3392
rect 522212 3408 522264 3460
rect 525064 3408 525116 3460
rect 539968 3408 540020 3460
rect 87696 3272 87748 3324
rect 171784 3272 171836 3324
rect 172796 3272 172848 3324
rect 225512 3340 225564 3392
rect 231308 3340 231360 3392
rect 262496 3340 262548 3392
rect 360660 3340 360712 3392
rect 385684 3340 385736 3392
rect 394240 3340 394292 3392
rect 210056 3272 210108 3324
rect 249064 3272 249116 3324
rect 370688 3272 370740 3324
rect 400956 3272 401008 3324
rect 431224 3272 431276 3324
rect 497372 3340 497424 3392
rect 29184 3204 29236 3256
rect 138112 3204 138164 3256
rect 146208 3204 146260 3256
rect 188804 3204 188856 3256
rect 235632 3204 235684 3256
rect 236644 3204 236696 3256
rect 265900 3204 265952 3256
rect 353944 3204 353996 3256
rect 375012 3204 375064 3256
rect 377404 3204 377456 3256
rect 412272 3204 412324 3256
rect 434628 3204 434680 3256
rect 502708 3272 502760 3324
rect 441252 3204 441304 3256
rect 523960 3204 524012 3256
rect 23848 3136 23900 3188
rect 134800 3136 134852 3188
rect 135536 3136 135588 3188
rect 183468 3136 183520 3188
rect 232228 3136 232280 3188
rect 257988 3136 258040 3188
rect 279332 3136 279384 3188
rect 384120 3136 384172 3188
rect 422852 3136 422904 3188
rect 438860 3136 438912 3188
rect 444288 3136 444340 3188
rect 534632 3136 534684 3188
rect 18512 3068 18564 3120
rect 13176 3000 13228 3052
rect 191932 3068 191984 3120
rect 204720 3068 204772 3120
rect 245660 3068 245712 3120
rect 247316 3068 247368 3120
rect 272616 3068 272668 3120
rect 273904 3068 273956 3120
rect 289360 3068 289412 3120
rect 347228 3068 347280 3120
rect 364340 3068 364392 3120
rect 387524 3068 387576 3120
rect 428188 3068 428240 3120
rect 448060 3068 448112 3120
rect 555884 3068 555936 3120
rect 188528 3000 188580 3052
rect 199384 3000 199436 3052
rect 242348 3000 242400 3052
rect 252652 3000 252704 3052
rect 276020 3000 276072 3052
rect 279240 3000 279292 3052
rect 292764 3000 292816 3052
rect 295156 3000 295208 3052
rect 302884 3000 302936 3052
rect 357256 3000 357308 3052
rect 380348 3000 380400 3052
rect 390928 3000 390980 3052
rect 433524 3000 433576 3052
rect 451188 3000 451240 3052
rect 561220 3000 561272 3052
rect 103612 2932 103664 2984
rect 181812 2932 181864 2984
rect 194140 2932 194192 2984
rect 238944 2932 238996 2984
rect 263232 2932 263284 2984
rect 282920 2932 282972 2984
rect 289912 2932 289964 2984
rect 299480 2932 299532 2984
rect 363972 2932 364024 2984
rect 390836 2932 390888 2984
rect 397276 2932 397328 2984
rect 444196 2932 444248 2984
rect 454776 2932 454828 2984
rect 571892 2932 571944 2984
rect 49332 2864 49384 2916
rect 114560 2864 114612 2916
rect 115480 2864 115532 2916
rect 119620 2864 119672 2916
rect 2596 2796 2648 2848
rect 121460 2796 121512 2848
rect 464160 2864 464212 2916
rect 131396 2796 131448 2848
rect 156880 2796 156932 2848
rect 215484 2796 215536 2848
rect 220728 2796 220780 2848
rect 255780 2796 255832 2848
rect 268568 2796 268620 2848
rect 55956 2728 56008 2780
rect 66168 2728 66220 2780
rect 85948 2728 86000 2780
rect 108948 2728 109000 2780
rect 115388 2728 115440 2780
rect 116860 2728 116912 2780
rect 144920 2728 144972 2780
rect 146944 2728 146996 2780
rect 151820 2728 151872 2780
rect 284576 2796 284628 2848
rect 286048 2728 286100 2780
rect 300492 2796 300544 2848
rect 296076 2728 296128 2780
rect 305828 2796 305880 2848
rect 309600 2796 309652 2848
rect 320180 2796 320232 2848
rect 321836 2796 321888 2848
rect 306380 2728 306432 2780
rect 323676 2728 323728 2780
rect 114560 2660 114612 2712
rect 114652 2660 114704 2712
rect 141516 2660 141568 2712
rect 141608 2660 141660 2712
rect 148232 2660 148284 2712
rect 327080 2796 327132 2848
rect 332416 2796 332468 2848
rect 330392 2728 330444 2780
rect 337752 2796 337804 2848
rect 350448 2796 350500 2848
rect 369676 2796 369728 2848
rect 380808 2796 380860 2848
rect 449532 2796 449584 2848
rect 458180 2796 458232 2848
rect 513380 2796 513432 2848
rect 417608 2728 417660 2780
rect 426348 2728 426400 2780
rect 467840 2728 467892 2780
rect 327080 2660 327132 2712
rect 337108 2660 337160 2712
rect 348424 2660 348476 2712
rect 437940 2660 437992 2712
rect 458180 2660 458232 2712
rect 35808 2592 35860 2644
rect 519636 2592 519688 2644
rect 15936 2524 15988 2576
rect 477684 2524 477736 2576
rect 25964 2456 26016 2508
rect 487712 2456 487764 2508
rect 1308 2388 1360 2440
rect 58624 2388 58676 2440
rect 68928 2388 68980 2440
rect 86868 2388 86920 2440
rect 92388 2388 92440 2440
rect 520372 2388 520424 2440
rect 79324 2320 79376 2372
rect 504548 2320 504600 2372
rect 99288 2252 99340 2304
rect 520464 2252 520516 2304
rect 89352 2184 89404 2236
rect 507860 2184 507912 2236
rect 95976 2116 96028 2168
rect 511264 2116 511316 2168
rect 102692 2048 102744 2100
rect 517980 2048 518032 2100
rect 115204 1980 115256 2032
rect 514760 1980 514812 2032
rect 82636 1912 82688 1964
rect 115572 1912 115624 1964
rect 116492 1912 116544 1964
rect 501144 1912 501196 1964
rect 113824 1844 113876 1896
rect 491300 1844 491352 1896
rect 22652 1776 22704 1828
rect 116584 1776 116636 1828
rect 117688 1776 117740 1828
rect 494428 1776 494480 1828
rect 118148 1708 118200 1760
rect 484400 1708 484452 1760
rect 168840 1640 168892 1692
rect 480996 1640 481048 1692
rect 9312 1572 9364 1624
rect 176660 1572 176712 1624
rect 333704 1572 333756 1624
rect 343088 1572 343140 1624
rect 343456 1572 343508 1624
rect 359004 1572 359056 1624
rect 106004 1504 106056 1556
rect 213828 1504 213880 1556
rect 340420 1504 340472 1556
rect 353760 1504 353812 1556
rect 32588 1436 32640 1488
rect 520740 1436 520792 1488
rect 19248 1368 19300 1420
rect 520096 1368 520148 1420
rect 72608 1300 72660 1352
rect 497832 1300 497884 1352
rect 71596 76 71648 128
rect 161664 76 161716 128
rect 34612 8 34664 60
rect 457444 8 457496 60
<< metal2 >>
rect 478 159200 534 160000
rect 1398 159200 1454 160000
rect 2410 159200 2466 160000
rect 3330 159200 3386 160000
rect 4342 159200 4398 160000
rect 5262 159200 5318 160000
rect 6274 159200 6330 160000
rect 7286 159200 7342 160000
rect 8206 159200 8262 160000
rect 9218 159200 9274 160000
rect 10138 159200 10194 160000
rect 11150 159200 11206 160000
rect 12162 159200 12218 160000
rect 13082 159200 13138 160000
rect 14094 159200 14150 160000
rect 15014 159200 15070 160000
rect 16026 159200 16082 160000
rect 17038 159200 17094 160000
rect 17958 159200 18014 160000
rect 18970 159200 19026 160000
rect 19890 159200 19946 160000
rect 20902 159200 20958 160000
rect 21914 159200 21970 160000
rect 22834 159200 22890 160000
rect 23846 159200 23902 160000
rect 24766 159200 24822 160000
rect 25778 159200 25834 160000
rect 26790 159200 26846 160000
rect 27710 159200 27766 160000
rect 28722 159200 28778 160000
rect 29642 159200 29698 160000
rect 30654 159200 30710 160000
rect 31666 159200 31722 160000
rect 32586 159200 32642 160000
rect 33598 159200 33654 160000
rect 34518 159200 34574 160000
rect 35530 159200 35586 160000
rect 36542 159200 36598 160000
rect 37462 159200 37518 160000
rect 38474 159200 38530 160000
rect 39394 159200 39450 160000
rect 40406 159200 40462 160000
rect 41326 159200 41382 160000
rect 42338 159200 42394 160000
rect 43350 159200 43406 160000
rect 44270 159200 44326 160000
rect 45282 159200 45338 160000
rect 46202 159200 46258 160000
rect 47214 159200 47270 160000
rect 48226 159200 48282 160000
rect 49146 159200 49202 160000
rect 50158 159200 50214 160000
rect 51078 159200 51134 160000
rect 52090 159200 52146 160000
rect 53102 159200 53158 160000
rect 54022 159200 54078 160000
rect 55034 159200 55090 160000
rect 55954 159200 56010 160000
rect 56966 159200 57022 160000
rect 57978 159200 58034 160000
rect 58898 159200 58954 160000
rect 59910 159200 59966 160000
rect 60830 159200 60886 160000
rect 61842 159200 61898 160000
rect 62854 159200 62910 160000
rect 63774 159200 63830 160000
rect 64786 159200 64842 160000
rect 65706 159200 65762 160000
rect 66718 159200 66774 160000
rect 67730 159200 67786 160000
rect 68650 159200 68706 160000
rect 69662 159200 69718 160000
rect 70582 159200 70638 160000
rect 71594 159200 71650 160000
rect 72606 159200 72662 160000
rect 73526 159200 73582 160000
rect 74538 159200 74594 160000
rect 75458 159200 75514 160000
rect 76470 159200 76526 160000
rect 77482 159200 77538 160000
rect 78402 159200 78458 160000
rect 79414 159200 79470 160000
rect 80334 159200 80390 160000
rect 81346 159200 81402 160000
rect 82266 159200 82322 160000
rect 83278 159200 83334 160000
rect 84290 159200 84346 160000
rect 85210 159200 85266 160000
rect 86222 159200 86278 160000
rect 87142 159200 87198 160000
rect 88154 159200 88210 160000
rect 89166 159200 89222 160000
rect 90086 159200 90142 160000
rect 91098 159200 91154 160000
rect 92018 159200 92074 160000
rect 93030 159200 93086 160000
rect 94042 159200 94098 160000
rect 94962 159200 95018 160000
rect 95974 159200 96030 160000
rect 96894 159200 96950 160000
rect 97906 159200 97962 160000
rect 98918 159200 98974 160000
rect 99838 159200 99894 160000
rect 100850 159200 100906 160000
rect 101770 159200 101826 160000
rect 102782 159200 102838 160000
rect 103794 159200 103850 160000
rect 104714 159200 104770 160000
rect 105726 159200 105782 160000
rect 106646 159200 106702 160000
rect 107658 159200 107714 160000
rect 108670 159200 108726 160000
rect 109590 159200 109646 160000
rect 110602 159200 110658 160000
rect 111522 159200 111578 160000
rect 112534 159200 112590 160000
rect 113546 159200 113602 160000
rect 114466 159200 114522 160000
rect 115478 159200 115534 160000
rect 116398 159200 116454 160000
rect 117410 159200 117466 160000
rect 118330 159200 118386 160000
rect 119342 159200 119398 160000
rect 120354 159200 120410 160000
rect 121274 159200 121330 160000
rect 122286 159200 122342 160000
rect 123206 159200 123262 160000
rect 124218 159200 124274 160000
rect 125230 159200 125286 160000
rect 126150 159200 126206 160000
rect 127162 159202 127218 160000
rect 127268 159310 127480 159338
rect 127268 159202 127296 159310
rect 127162 159200 127296 159202
rect 492 155242 520 159200
rect 1412 155281 1440 159200
rect 1398 155272 1454 155281
rect 480 155236 532 155242
rect 480 155178 532 155184
rect 1308 155236 1360 155242
rect 1398 155207 1454 155216
rect 1308 155178 1360 155184
rect 1320 154630 1348 155178
rect 1308 154624 1360 154630
rect 1308 154566 1360 154572
rect 1320 2446 1348 154566
rect 2424 152561 2452 159200
rect 3146 157584 3202 157593
rect 3146 157519 3202 157528
rect 2410 152552 2466 152561
rect 2410 152487 2466 152496
rect 3160 152425 3188 157519
rect 3344 156641 3372 159200
rect 3330 156632 3386 156641
rect 3330 156567 3386 156576
rect 4356 155854 4384 159200
rect 4344 155848 4396 155854
rect 4344 155790 4396 155796
rect 5276 155417 5304 159200
rect 6288 156670 6316 159200
rect 6276 156664 6328 156670
rect 6276 156606 6328 156612
rect 5262 155408 5318 155417
rect 5262 155343 5318 155352
rect 3238 152960 3294 152969
rect 3238 152895 3294 152904
rect 3146 152416 3202 152425
rect 3146 152351 3202 152360
rect 3252 151910 3280 152895
rect 7300 152522 7328 159200
rect 8220 155242 8248 159200
rect 8208 155236 8260 155242
rect 8208 155178 8260 155184
rect 9232 153882 9260 159200
rect 10152 156738 10180 159200
rect 11164 158710 11192 159200
rect 11152 158704 11204 158710
rect 11152 158646 11204 158652
rect 10140 156732 10192 156738
rect 10140 156674 10192 156680
rect 12176 155922 12204 159200
rect 12440 158228 12492 158234
rect 12440 158170 12492 158176
rect 12164 155916 12216 155922
rect 12164 155858 12216 155864
rect 12452 155854 12480 158170
rect 12440 155848 12492 155854
rect 12440 155790 12492 155796
rect 13096 153950 13124 159200
rect 14108 155310 14136 159200
rect 15028 158930 15056 159200
rect 15028 158902 15240 158930
rect 15212 158846 15240 158902
rect 15200 158840 15252 158846
rect 15200 158782 15252 158788
rect 16040 155582 16068 159200
rect 16028 155576 16080 155582
rect 16028 155518 16080 155524
rect 14096 155304 14148 155310
rect 14096 155246 14148 155252
rect 17052 154329 17080 159200
rect 17972 156806 18000 159200
rect 18984 158166 19012 159200
rect 18972 158160 19024 158166
rect 18972 158102 19024 158108
rect 17960 156800 18012 156806
rect 17960 156742 18012 156748
rect 17866 156088 17922 156097
rect 17866 156023 17922 156032
rect 17880 155854 17908 156023
rect 17868 155848 17920 155854
rect 17868 155790 17920 155796
rect 19904 155378 19932 159200
rect 19892 155372 19944 155378
rect 19892 155314 19944 155320
rect 17038 154320 17094 154329
rect 17038 154255 17094 154264
rect 20916 154018 20944 159200
rect 20904 154012 20956 154018
rect 20904 153954 20956 153960
rect 13084 153944 13136 153950
rect 13084 153886 13136 153892
rect 9220 153876 9272 153882
rect 9220 153818 9272 153824
rect 9402 153368 9458 153377
rect 9402 153303 9458 153312
rect 7288 152516 7340 152522
rect 7288 152458 7340 152464
rect 9416 151994 9444 153303
rect 12808 153264 12860 153270
rect 12808 153206 12860 153212
rect 19706 153232 19762 153241
rect 12820 151994 12848 153206
rect 19706 153167 19762 153176
rect 19720 151994 19748 153167
rect 21928 152590 21956 159200
rect 22848 158778 22876 159200
rect 22836 158772 22888 158778
rect 22836 158714 22888 158720
rect 23860 155446 23888 159200
rect 24780 155553 24808 159200
rect 25792 156874 25820 159200
rect 26804 158914 26832 159200
rect 26792 158908 26844 158914
rect 26792 158850 26844 158856
rect 25780 156868 25832 156874
rect 25780 156810 25832 156816
rect 24766 155544 24822 155553
rect 27724 155514 27752 159200
rect 24766 155479 24822 155488
rect 27712 155508 27764 155514
rect 27712 155450 27764 155456
rect 23848 155440 23900 155446
rect 23848 155382 23900 155388
rect 24860 155304 24912 155310
rect 24860 155246 24912 155252
rect 24872 152930 24900 155246
rect 28736 154086 28764 159200
rect 29656 155174 29684 159200
rect 30668 157690 30696 159200
rect 30656 157684 30708 157690
rect 30656 157626 30708 157632
rect 31680 155310 31708 159200
rect 31668 155304 31720 155310
rect 31668 155246 31720 155252
rect 29644 155168 29696 155174
rect 29644 155110 29696 155116
rect 31668 155168 31720 155174
rect 31668 155110 31720 155116
rect 28724 154080 28776 154086
rect 28724 154022 28776 154028
rect 30010 153504 30066 153513
rect 30010 153439 30066 153448
rect 26606 153368 26662 153377
rect 26606 153303 26662 153312
rect 24860 152924 24912 152930
rect 24860 152866 24912 152872
rect 21916 152584 21968 152590
rect 21916 152526 21968 152532
rect 26620 151994 26648 153303
rect 26700 153264 26752 153270
rect 26700 153206 26752 153212
rect 9108 151966 9444 151994
rect 12512 151966 12848 151994
rect 19412 151966 19748 151994
rect 26312 151966 26648 151994
rect 3240 151904 3292 151910
rect 3240 151846 3292 151852
rect 3516 151836 3568 151842
rect 3516 151778 3568 151784
rect 2964 151768 3016 151774
rect 2964 151710 3016 151716
rect 2976 143857 3004 151710
rect 3148 151700 3200 151706
rect 3148 151642 3200 151648
rect 2962 143848 3018 143857
rect 2962 143783 3018 143792
rect 3160 142154 3188 151642
rect 3240 151632 3292 151638
rect 3240 151574 3292 151580
rect 3252 146742 3280 151574
rect 3330 149968 3386 149977
rect 3330 149903 3386 149912
rect 3240 146736 3292 146742
rect 3240 146678 3292 146684
rect 3160 142126 3280 142154
rect 3252 139369 3280 142126
rect 3238 139360 3294 139369
rect 3238 139295 3294 139304
rect 3344 134745 3372 149903
rect 3424 149116 3476 149122
rect 3424 149058 3476 149064
rect 3436 146826 3464 149058
rect 3528 148481 3556 151778
rect 16008 151570 16344 151586
rect 26712 151570 26740 153206
rect 30024 151994 30052 153439
rect 31680 152658 31708 155110
rect 32600 154154 32628 159200
rect 33612 155922 33640 159200
rect 34532 158302 34560 159200
rect 34520 158296 34572 158302
rect 34520 158238 34572 158244
rect 34702 156224 34758 156233
rect 34702 156159 34758 156168
rect 34716 155922 34744 156159
rect 33600 155916 33652 155922
rect 33600 155858 33652 155864
rect 34704 155916 34756 155922
rect 34704 155858 34756 155864
rect 35544 154222 35572 159200
rect 36556 155689 36584 159200
rect 36542 155680 36598 155689
rect 36542 155615 36598 155624
rect 35532 154216 35584 154222
rect 35532 154158 35584 154164
rect 32588 154148 32640 154154
rect 32588 154090 32640 154096
rect 37476 152697 37504 159200
rect 38488 157758 38516 159200
rect 38476 157752 38528 157758
rect 38476 157694 38528 157700
rect 39408 155650 39436 159200
rect 39396 155644 39448 155650
rect 39396 155586 39448 155592
rect 40420 154290 40448 159200
rect 40408 154284 40460 154290
rect 40408 154226 40460 154232
rect 39854 153640 39910 153649
rect 39854 153575 39910 153584
rect 37462 152688 37518 152697
rect 31668 152652 31720 152658
rect 37462 152623 37518 152632
rect 31668 152594 31720 152600
rect 29716 151966 30052 151994
rect 39868 151858 39896 153575
rect 41340 152726 41368 159200
rect 42352 156942 42380 159200
rect 42340 156936 42392 156942
rect 42340 156878 42392 156884
rect 43364 155854 43392 159200
rect 43352 155848 43404 155854
rect 43352 155790 43404 155796
rect 44284 154358 44312 159200
rect 44272 154352 44324 154358
rect 44272 154294 44324 154300
rect 45296 152862 45324 159200
rect 45284 152856 45336 152862
rect 45284 152798 45336 152804
rect 46216 152794 46244 159200
rect 47228 157826 47256 159200
rect 47216 157820 47268 157826
rect 47216 157762 47268 157768
rect 48240 154426 48268 159200
rect 48228 154420 48280 154426
rect 48228 154362 48280 154368
rect 46756 153264 46808 153270
rect 46756 153206 46808 153212
rect 46204 152788 46256 152794
rect 46204 152730 46256 152736
rect 41328 152720 41380 152726
rect 41328 152662 41380 152668
rect 43516 151978 43852 151994
rect 43516 151972 43864 151978
rect 43516 151966 43812 151972
rect 43812 151914 43864 151920
rect 46768 151858 46796 153206
rect 49160 152998 49188 159200
rect 50172 156777 50200 159200
rect 51092 158522 51120 159200
rect 51092 158494 51212 158522
rect 51080 158364 51132 158370
rect 51080 158306 51132 158312
rect 50158 156768 50214 156777
rect 50158 156703 50214 156712
rect 51092 155854 51120 158306
rect 51080 155848 51132 155854
rect 51080 155790 51132 155796
rect 51184 155106 51212 158494
rect 52104 155825 52132 159200
rect 53116 157010 53144 159200
rect 53104 157004 53156 157010
rect 53104 156946 53156 156952
rect 52090 155816 52146 155825
rect 52090 155751 52146 155760
rect 51172 155100 51224 155106
rect 51172 155042 51224 155048
rect 50618 153776 50674 153785
rect 50618 153711 50674 153720
rect 49148 152992 49200 152998
rect 49148 152934 49200 152940
rect 50632 151994 50660 153711
rect 54036 153066 54064 159200
rect 55048 155174 55076 159200
rect 55968 155786 55996 159200
rect 56980 157078 57008 159200
rect 57992 157146 58020 159200
rect 58912 157894 58940 159200
rect 58900 157888 58952 157894
rect 58900 157830 58952 157836
rect 57980 157140 58032 157146
rect 57980 157082 58032 157088
rect 56968 157072 57020 157078
rect 56968 157014 57020 157020
rect 55956 155780 56008 155786
rect 55956 155722 56008 155728
rect 55036 155168 55088 155174
rect 55036 155110 55088 155116
rect 59924 154494 59952 159200
rect 59912 154488 59964 154494
rect 59912 154430 59964 154436
rect 60844 153134 60872 159200
rect 60832 153128 60884 153134
rect 60832 153070 60884 153076
rect 54024 153060 54076 153066
rect 54024 153002 54076 153008
rect 61856 152454 61884 159200
rect 62868 155038 62896 159200
rect 63788 155854 63816 159200
rect 64800 156913 64828 159200
rect 65720 157214 65748 159200
rect 65708 157208 65760 157214
rect 65708 157150 65760 157156
rect 64786 156904 64842 156913
rect 64786 156839 64842 156848
rect 66732 155922 66760 159200
rect 67364 158432 67416 158438
rect 67364 158374 67416 158380
rect 66720 155916 66772 155922
rect 66720 155858 66772 155864
rect 63776 155848 63828 155854
rect 63776 155790 63828 155796
rect 67376 155106 67404 158374
rect 67364 155100 67416 155106
rect 67364 155042 67416 155048
rect 62856 155032 62908 155038
rect 62856 154974 62908 154980
rect 67744 154562 67772 159200
rect 68664 157282 68692 159200
rect 68652 157276 68704 157282
rect 68652 157218 68704 157224
rect 67732 154556 67784 154562
rect 67732 154498 67784 154504
rect 61844 152448 61896 152454
rect 61844 152390 61896 152396
rect 69676 152386 69704 159200
rect 70400 158568 70452 158574
rect 70400 158510 70452 158516
rect 70412 155174 70440 158510
rect 70400 155168 70452 155174
rect 70400 155110 70452 155116
rect 70596 154601 70624 159200
rect 71608 154902 71636 159200
rect 71596 154896 71648 154902
rect 71596 154838 71648 154844
rect 70582 154592 70638 154601
rect 70582 154527 70638 154536
rect 72620 153202 72648 159200
rect 73540 157350 73568 159200
rect 73528 157344 73580 157350
rect 73528 157286 73580 157292
rect 74552 155718 74580 159200
rect 75000 158500 75052 158506
rect 75000 158442 75052 158448
rect 74540 155712 74592 155718
rect 74540 155654 74592 155660
rect 75012 155038 75040 158442
rect 75472 155961 75500 159200
rect 76484 156602 76512 159200
rect 76472 156596 76524 156602
rect 76472 156538 76524 156544
rect 75458 155952 75514 155961
rect 75458 155887 75514 155896
rect 75000 155032 75052 155038
rect 75000 154974 75052 154980
rect 72608 153196 72660 153202
rect 72608 153138 72660 153144
rect 69664 152380 69716 152386
rect 69664 152322 69716 152328
rect 77496 152318 77524 159200
rect 78416 153814 78444 159200
rect 78404 153808 78456 153814
rect 78404 153750 78456 153756
rect 79428 153746 79456 159200
rect 79416 153740 79468 153746
rect 79416 153682 79468 153688
rect 77484 152312 77536 152318
rect 77484 152254 77536 152260
rect 80348 152250 80376 159200
rect 81360 156534 81388 159200
rect 82280 157962 82308 159200
rect 82820 158636 82872 158642
rect 82820 158578 82872 158584
rect 82268 157956 82320 157962
rect 82268 157898 82320 157904
rect 81348 156528 81400 156534
rect 81348 156470 81400 156476
rect 82832 155922 82860 158578
rect 82820 155916 82872 155922
rect 82820 155858 82872 155864
rect 83292 155106 83320 159200
rect 84304 156466 84332 159200
rect 84292 156460 84344 156466
rect 84292 156402 84344 156408
rect 83280 155100 83332 155106
rect 83280 155042 83332 155048
rect 81162 153912 81218 153921
rect 81162 153847 81218 153856
rect 80336 152244 80388 152250
rect 80336 152186 80388 152192
rect 50324 151966 50660 151994
rect 57224 151978 57560 151994
rect 60720 151978 60872 151994
rect 64124 151978 64460 151994
rect 67376 151978 67528 151994
rect 57224 151972 57572 151978
rect 57224 151966 57520 151972
rect 60720 151972 60884 151978
rect 60720 151966 60832 151972
rect 57520 151914 57572 151920
rect 64124 151972 64472 151978
rect 64124 151966 64420 151972
rect 60832 151914 60884 151920
rect 64420 151914 64472 151920
rect 67364 151972 67528 151978
rect 67416 151966 67528 151972
rect 74428 151978 74580 151994
rect 77832 151978 78168 151994
rect 74428 151972 74592 151978
rect 74428 151966 74540 151972
rect 67364 151914 67416 151920
rect 77832 151972 78180 151978
rect 77832 151966 78128 151972
rect 74540 151914 74592 151920
rect 78128 151914 78180 151920
rect 39868 151830 40020 151858
rect 46768 151830 46920 151858
rect 81176 151722 81204 153847
rect 85224 152182 85252 159200
rect 86236 154698 86264 159200
rect 87156 154970 87184 159200
rect 87144 154964 87196 154970
rect 87144 154906 87196 154912
rect 86224 154692 86276 154698
rect 86224 154634 86276 154640
rect 88062 154048 88118 154057
rect 88062 153983 88118 153992
rect 85212 152176 85264 152182
rect 85212 152118 85264 152124
rect 84732 151978 85068 151994
rect 84732 151972 85080 151978
rect 84732 151966 85028 151972
rect 85028 151914 85080 151920
rect 88076 151858 88104 153983
rect 88168 152114 88196 159200
rect 89180 157049 89208 159200
rect 89166 157040 89222 157049
rect 89166 156975 89222 156984
rect 90100 155174 90128 159200
rect 90088 155168 90140 155174
rect 91112 155145 91140 159200
rect 92032 156398 92060 159200
rect 92020 156392 92072 156398
rect 92020 156334 92072 156340
rect 90088 155110 90140 155116
rect 91098 155136 91154 155145
rect 91098 155071 91154 155080
rect 91008 154692 91060 154698
rect 91008 154634 91060 154640
rect 88156 152108 88208 152114
rect 88156 152050 88208 152056
rect 91020 151978 91048 154634
rect 91926 154184 91982 154193
rect 91926 154119 91982 154128
rect 91940 151994 91968 154119
rect 93044 153610 93072 159200
rect 94056 158030 94084 159200
rect 94044 158024 94096 158030
rect 94044 157966 94096 157972
rect 94976 153678 95004 159200
rect 94964 153672 95016 153678
rect 94964 153614 95016 153620
rect 93032 153604 93084 153610
rect 93032 153546 93084 153552
rect 92204 153264 92256 153270
rect 92204 153206 92256 153212
rect 91008 151972 91060 151978
rect 91632 151966 91968 151994
rect 91008 151914 91060 151920
rect 88076 151830 88228 151858
rect 81176 151694 81328 151722
rect 16008 151564 16356 151570
rect 16008 151558 16304 151564
rect 16304 151506 16356 151512
rect 26700 151564 26752 151570
rect 26700 151506 26752 151512
rect 5080 151496 5132 151502
rect 33506 151464 33562 151473
rect 5080 151438 5132 151444
rect 3792 151428 3844 151434
rect 3792 151370 3844 151376
rect 3608 151360 3660 151366
rect 3608 151302 3660 151308
rect 3514 148472 3570 148481
rect 3514 148407 3570 148416
rect 3436 146798 3556 146826
rect 3424 146736 3476 146742
rect 3424 146678 3476 146684
rect 3330 134736 3386 134745
rect 3330 134671 3386 134680
rect 3436 102785 3464 146678
rect 3528 107273 3556 146798
rect 3620 111897 3648 151302
rect 3700 150408 3752 150414
rect 3700 150350 3752 150356
rect 3712 116521 3740 150350
rect 3804 121009 3832 151370
rect 4068 150476 4120 150482
rect 4068 150418 4120 150424
rect 3884 150340 3936 150346
rect 3884 150282 3936 150288
rect 3896 125633 3924 150282
rect 3976 150272 4028 150278
rect 3976 150214 4028 150220
rect 3988 130121 4016 150214
rect 3974 130112 4030 130121
rect 3974 130047 4030 130056
rect 3882 125624 3938 125633
rect 3882 125559 3938 125568
rect 3790 121000 3846 121009
rect 3790 120935 3846 120944
rect 3698 116512 3754 116521
rect 3698 116447 3754 116456
rect 3606 111888 3662 111897
rect 3606 111823 3662 111832
rect 3514 107264 3570 107273
rect 3514 107199 3570 107208
rect 3422 102776 3478 102785
rect 3422 102711 3478 102720
rect 3790 98152 3846 98161
rect 3790 98087 3846 98096
rect 3422 93664 3478 93673
rect 3422 93599 3478 93608
rect 3330 66192 3386 66201
rect 3330 66127 3386 66136
rect 3238 61568 3294 61577
rect 3238 61503 3294 61512
rect 2778 57080 2834 57089
rect 2778 57015 2834 57024
rect 2792 56914 2820 57015
rect 2780 56908 2832 56914
rect 2780 56850 2832 56856
rect 3146 52456 3202 52465
rect 3146 52391 3202 52400
rect 3054 47968 3110 47977
rect 3054 47903 3110 47912
rect 2962 43344 3018 43353
rect 2962 43279 3018 43288
rect 2870 38720 2926 38729
rect 2870 38655 2926 38664
rect 2778 29608 2834 29617
rect 2778 29543 2834 29552
rect 2792 5778 2820 29543
rect 2884 5846 2912 38655
rect 2976 5914 3004 43279
rect 2964 5908 3016 5914
rect 2964 5850 3016 5856
rect 2872 5840 2924 5846
rect 2872 5782 2924 5788
rect 2780 5772 2832 5778
rect 2780 5714 2832 5720
rect 3068 5574 3096 47903
rect 3160 5642 3188 52391
rect 3252 13598 3280 61503
rect 3344 17950 3372 66127
rect 3332 17944 3384 17950
rect 3332 17886 3384 17892
rect 3240 13592 3292 13598
rect 3240 13534 3292 13540
rect 3332 8968 3384 8974
rect 3332 8910 3384 8916
rect 3238 6760 3294 6769
rect 3238 6695 3294 6704
rect 3148 5636 3200 5642
rect 3148 5578 3200 5584
rect 3056 5568 3108 5574
rect 3056 5510 3108 5516
rect 3252 5302 3280 6695
rect 3240 5296 3292 5302
rect 3240 5238 3292 5244
rect 3344 4962 3372 8910
rect 3436 5438 3464 93599
rect 3698 89040 3754 89049
rect 3698 88975 3754 88984
rect 3606 84416 3662 84425
rect 3606 84351 3662 84360
rect 3514 75304 3570 75313
rect 3514 75239 3570 75248
rect 3424 5432 3476 5438
rect 3424 5374 3476 5380
rect 3528 5166 3556 75239
rect 3620 24886 3648 84351
rect 3712 30326 3740 88975
rect 3804 40050 3832 98087
rect 3882 79928 3938 79937
rect 3882 79863 3938 79872
rect 3792 40044 3844 40050
rect 3792 39986 3844 39992
rect 3790 34232 3846 34241
rect 3790 34167 3846 34176
rect 3700 30320 3752 30326
rect 3700 30262 3752 30268
rect 3698 25120 3754 25129
rect 3698 25055 3754 25064
rect 3608 24880 3660 24886
rect 3608 24822 3660 24828
rect 3606 20496 3662 20505
rect 3606 20431 3662 20440
rect 3620 8974 3648 20431
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 3608 8832 3660 8838
rect 3608 8774 3660 8780
rect 3516 5160 3568 5166
rect 3516 5102 3568 5108
rect 3620 5001 3648 8774
rect 3712 5370 3740 25055
rect 3804 5710 3832 34167
rect 3896 21418 3924 79863
rect 3974 70816 4030 70825
rect 3974 70751 4030 70760
rect 3884 21412 3936 21418
rect 3884 21354 3936 21360
rect 3882 15872 3938 15881
rect 3882 15807 3938 15816
rect 3896 6914 3924 15807
rect 3988 12918 4016 70751
rect 3976 12912 4028 12918
rect 3976 12854 4028 12860
rect 3974 11384 4030 11393
rect 3974 11319 4030 11328
rect 3988 8650 4016 11319
rect 4080 8838 4108 150418
rect 5092 149122 5120 151438
rect 33212 151422 33506 151450
rect 33506 151399 33562 151408
rect 92216 151337 92244 153206
rect 95988 152046 96016 159200
rect 96908 154698 96936 159200
rect 97920 154873 97948 159200
rect 97906 154864 97962 154873
rect 97906 154799 97962 154808
rect 98932 154766 98960 159200
rect 99852 156330 99880 159200
rect 99840 156324 99892 156330
rect 99840 156266 99892 156272
rect 98920 154760 98972 154766
rect 98920 154702 98972 154708
rect 96896 154692 96948 154698
rect 96896 154634 96948 154640
rect 100864 153542 100892 159200
rect 101784 155038 101812 159200
rect 101772 155032 101824 155038
rect 101772 154974 101824 154980
rect 100852 153536 100904 153542
rect 100852 153478 100904 153484
rect 102796 153474 102824 159200
rect 102784 153468 102836 153474
rect 102784 153410 102836 153416
rect 103808 152833 103836 159200
rect 104728 157486 104756 159200
rect 104716 157480 104768 157486
rect 104716 157422 104768 157428
rect 105740 155009 105768 159200
rect 105726 155000 105782 155009
rect 105726 154935 105782 154944
rect 106660 154834 106688 159200
rect 107672 156262 107700 159200
rect 107660 156256 107712 156262
rect 107660 156198 107712 156204
rect 106648 154828 106700 154834
rect 106648 154770 106700 154776
rect 106188 154624 106240 154630
rect 106188 154566 106240 154572
rect 106200 154465 106228 154566
rect 106186 154456 106242 154465
rect 106186 154391 106242 154400
rect 108684 152969 108712 159200
rect 109604 153406 109632 159200
rect 110616 154630 110644 159200
rect 111536 156194 111564 159200
rect 112548 158098 112576 159200
rect 112536 158092 112588 158098
rect 112536 158034 112588 158040
rect 113560 157554 113588 159200
rect 113548 157548 113600 157554
rect 113548 157490 113600 157496
rect 111524 156188 111576 156194
rect 111524 156130 111576 156136
rect 110604 154624 110656 154630
rect 110604 154566 110656 154572
rect 114480 153406 114508 159200
rect 109592 153400 109644 153406
rect 109592 153342 109644 153348
rect 114468 153400 114520 153406
rect 114468 153342 114520 153348
rect 112444 153332 112496 153338
rect 112444 153274 112496 153280
rect 108948 153264 109000 153270
rect 108948 153206 109000 153212
rect 108670 152960 108726 152969
rect 108670 152895 108726 152904
rect 103794 152824 103850 152833
rect 103794 152759 103850 152768
rect 95976 152040 96028 152046
rect 95036 151978 95188 151994
rect 108960 151994 108988 153206
rect 112456 151994 112484 153274
rect 112536 153264 112588 153270
rect 112536 153206 112588 153212
rect 95976 151982 96028 151988
rect 105340 151978 105676 151994
rect 95036 151972 95200 151978
rect 95036 151966 95148 151972
rect 105340 151972 105688 151978
rect 105340 151966 105636 151972
rect 95148 151914 95200 151920
rect 108836 151966 108988 151994
rect 112240 151966 112484 151994
rect 105636 151914 105688 151920
rect 102046 151872 102102 151881
rect 101936 151830 102046 151858
rect 102046 151807 102102 151816
rect 112548 151814 112576 153206
rect 115492 151978 115520 159200
rect 116412 156126 116440 159200
rect 116400 156120 116452 156126
rect 116400 156062 116452 156068
rect 117424 154834 117452 159200
rect 118344 155582 118372 159200
rect 119356 156058 119384 159200
rect 119436 157412 119488 157418
rect 119436 157354 119488 157360
rect 119344 156052 119396 156058
rect 119344 155994 119396 156000
rect 117964 155576 118016 155582
rect 117964 155518 118016 155524
rect 118332 155576 118384 155582
rect 118332 155518 118384 155524
rect 117412 154828 117464 154834
rect 117412 154770 117464 154776
rect 117976 153270 118004 155518
rect 117780 153264 117832 153270
rect 117780 153206 117832 153212
rect 117964 153264 118016 153270
rect 117964 153206 118016 153212
rect 115754 152416 115810 152425
rect 115754 152351 115810 152360
rect 115480 151972 115532 151978
rect 115480 151914 115532 151920
rect 115112 151904 115164 151910
rect 115112 151846 115164 151852
rect 112548 151786 112668 151814
rect 98826 151464 98882 151473
rect 98532 151422 98826 151450
rect 98826 151399 98882 151408
rect 112442 151464 112498 151473
rect 112442 151399 112498 151408
rect 112536 151428 112588 151434
rect 23110 151328 23166 151337
rect 5552 151286 5704 151314
rect 22816 151286 23110 151314
rect 5552 150482 5580 151286
rect 36910 151328 36966 151337
rect 36616 151286 36910 151314
rect 23110 151263 23166 151272
rect 53930 151328 53986 151337
rect 53820 151286 53930 151314
rect 36910 151263 36966 151272
rect 71318 151328 71374 151337
rect 71024 151286 71318 151314
rect 53930 151263 53986 151272
rect 71318 151263 71374 151272
rect 92202 151328 92258 151337
rect 92202 151263 92258 151272
rect 112456 150521 112484 151399
rect 112536 151370 112588 151376
rect 112442 150512 112498 150521
rect 5540 150476 5592 150482
rect 112442 150447 112498 150456
rect 5540 150418 5592 150424
rect 112444 150408 112496 150414
rect 112444 150350 112496 150356
rect 5080 149116 5132 149122
rect 5080 149058 5132 149064
rect 112456 66230 112484 150350
rect 112548 74594 112576 151370
rect 112640 146266 112668 151786
rect 114192 151768 114244 151774
rect 114192 151710 114244 151716
rect 112904 151632 112956 151638
rect 112904 151574 112956 151580
rect 112812 151496 112864 151502
rect 112812 151438 112864 151444
rect 112628 146260 112680 146266
rect 112628 146202 112680 146208
rect 112824 146010 112852 151438
rect 112916 149394 112944 151574
rect 112996 151360 113048 151366
rect 112996 151302 113048 151308
rect 112904 149388 112956 149394
rect 112904 149330 112956 149336
rect 112640 145982 112852 146010
rect 112640 94382 112668 145982
rect 113008 142154 113036 151302
rect 113916 151156 113968 151162
rect 113916 151098 113968 151104
rect 113822 150648 113878 150657
rect 113822 150583 113878 150592
rect 112732 142126 113036 142154
rect 112732 114034 112760 142126
rect 112720 114028 112772 114034
rect 112720 113970 112772 113976
rect 112628 94376 112680 94382
rect 112628 94318 112680 94324
rect 112536 74588 112588 74594
rect 112536 74530 112588 74536
rect 112444 66224 112496 66230
rect 112444 66166 112496 66172
rect 4804 56908 4856 56914
rect 4804 56850 4856 56856
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 3988 8622 4108 8650
rect 3896 6886 4016 6914
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 3988 5506 4016 6886
rect 3976 5500 4028 5506
rect 3976 5442 4028 5448
rect 3700 5364 3752 5370
rect 3700 5306 3752 5312
rect 4080 5234 4108 8622
rect 4816 6089 4844 56850
rect 4896 40044 4948 40050
rect 4896 39986 4948 39992
rect 4802 6080 4858 6089
rect 4802 6015 4858 6024
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 3606 4992 3662 5001
rect 3332 4956 3384 4962
rect 3606 4927 3662 4936
rect 3332 4898 3384 4904
rect 4908 4826 4936 39986
rect 112536 38684 112588 38690
rect 112536 38626 112588 38632
rect 4988 30320 5040 30326
rect 4988 30262 5040 30268
rect 5000 5098 5028 30262
rect 5080 24880 5132 24886
rect 5080 24822 5132 24828
rect 4988 5092 5040 5098
rect 4988 5034 5040 5040
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 5092 4758 5120 24822
rect 5172 21412 5224 21418
rect 5172 21354 5224 21360
rect 5080 4752 5132 4758
rect 5080 4694 5132 4700
rect 5184 4690 5212 21354
rect 5264 17944 5316 17950
rect 5264 17886 5316 17892
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5276 4554 5304 17886
rect 5448 13592 5500 13598
rect 5448 13534 5500 13540
rect 5356 12912 5408 12918
rect 5356 12854 5408 12860
rect 5368 4622 5396 12854
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 5264 4548 5316 4554
rect 5264 4490 5316 4496
rect 5460 4486 5488 13534
rect 112444 5976 112496 5982
rect 112444 5918 112496 5924
rect 112456 5438 112484 5918
rect 112548 5522 112576 38626
rect 113732 31816 113784 31822
rect 113732 31758 113784 31764
rect 113640 29028 113692 29034
rect 113640 28970 113692 28976
rect 112628 27668 112680 27674
rect 112628 27610 112680 27616
rect 112640 16574 112668 27610
rect 113652 26234 113680 28970
rect 113744 27538 113772 31758
rect 113732 27532 113784 27538
rect 113732 27474 113784 27480
rect 113652 26206 113772 26234
rect 112640 16546 112760 16574
rect 112732 5982 112760 16546
rect 113640 13864 113692 13870
rect 113640 13806 113692 13812
rect 112720 5976 112772 5982
rect 112720 5918 112772 5924
rect 112548 5494 112760 5522
rect 112444 5432 112496 5438
rect 112444 5374 112496 5380
rect 112628 5432 112680 5438
rect 112628 5374 112680 5380
rect 112640 4706 112668 5374
rect 112332 4678 112668 4706
rect 39302 4584 39358 4593
rect 39008 4542 39302 4570
rect 45926 4584 45982 4593
rect 45632 4542 45926 4570
rect 39302 4519 39358 4528
rect 52458 4584 52514 4593
rect 52348 4542 52458 4570
rect 45926 4519 45982 4528
rect 52458 4519 52514 4528
rect 112732 4486 112760 5494
rect 113652 4962 113680 13806
rect 113744 5574 113772 26206
rect 113732 5568 113784 5574
rect 113732 5510 113784 5516
rect 113640 4956 113692 4962
rect 113640 4898 113692 4904
rect 5448 4480 5500 4486
rect 112720 4480 112772 4486
rect 75826 4448 75882 4457
rect 5448 4422 5500 4428
rect 42320 4418 42656 4434
rect 42320 4412 42668 4418
rect 42320 4406 42616 4412
rect 75716 4406 75826 4434
rect 112720 4422 112772 4428
rect 75826 4383 75882 4392
rect 42616 4354 42668 4360
rect 62672 4344 62724 4350
rect 62376 4292 62672 4298
rect 62376 4286 62724 4292
rect 62376 4270 62712 4286
rect 65688 4282 66024 4298
rect 65688 4276 66036 4282
rect 65688 4270 65984 4276
rect 65984 4218 66036 4224
rect 66168 4276 66220 4282
rect 66168 4218 66220 4224
rect 2964 4208 3016 4214
rect 2964 4150 3016 4156
rect 2596 2848 2648 2854
rect 2596 2790 2648 2796
rect 1308 2440 1360 2446
rect 1308 2382 1360 2388
rect 2608 800 2636 2790
rect 2976 2281 3004 4150
rect 5704 4134 6040 4162
rect 6012 2689 6040 4134
rect 7840 4140 7892 4146
rect 9016 4134 9352 4162
rect 7840 4082 7892 4088
rect 5998 2680 6054 2689
rect 5998 2615 6054 2624
rect 2962 2272 3018 2281
rect 2962 2207 3018 2216
rect 7852 800 7880 4082
rect 9324 1630 9352 4134
rect 12314 3890 12342 4148
rect 15640 4134 15976 4162
rect 18952 4134 19288 4162
rect 22356 4134 22692 4162
rect 25668 4134 26004 4162
rect 12314 3862 12388 3890
rect 12360 2553 12388 3862
rect 13176 3052 13228 3058
rect 13176 2994 13228 3000
rect 12346 2544 12402 2553
rect 12346 2479 12402 2488
rect 9312 1624 9364 1630
rect 9312 1566 9364 1572
rect 13188 800 13216 2994
rect 15948 2582 15976 4134
rect 18512 3120 18564 3126
rect 18512 3062 18564 3068
rect 15936 2576 15988 2582
rect 15936 2518 15988 2524
rect 18524 800 18552 3062
rect 19260 1426 19288 4134
rect 22664 1834 22692 4134
rect 23848 3188 23900 3194
rect 23848 3130 23900 3136
rect 22652 1828 22704 1834
rect 22652 1770 22704 1776
rect 19248 1420 19300 1426
rect 19248 1362 19300 1368
rect 23860 800 23888 3130
rect 25976 2514 26004 4134
rect 28966 3890 28994 4148
rect 32292 4134 32628 4162
rect 35696 4134 35848 4162
rect 49036 4134 49372 4162
rect 55660 4134 55996 4162
rect 28920 3862 28994 3890
rect 25964 2508 26016 2514
rect 25964 2450 26016 2456
rect 28920 2417 28948 3862
rect 29184 3256 29236 3262
rect 29184 3198 29236 3204
rect 28906 2408 28962 2417
rect 28906 2343 28962 2352
rect 29196 800 29224 3198
rect 32600 1494 32628 4134
rect 35820 2650 35848 4134
rect 45100 4072 45152 4078
rect 45100 4014 45152 4020
rect 39764 3528 39816 3534
rect 39764 3470 39816 3476
rect 35808 2644 35860 2650
rect 35808 2586 35860 2592
rect 32588 1488 32640 1494
rect 32588 1430 32640 1436
rect 34532 870 34652 898
rect 34532 800 34560 870
rect 2594 0 2650 800
rect 7838 0 7894 800
rect 13174 0 13230 800
rect 18510 0 18566 800
rect 23846 0 23902 800
rect 29182 0 29238 800
rect 34518 0 34574 800
rect 34624 66 34652 870
rect 39776 800 39804 3470
rect 45112 800 45140 4014
rect 49344 2922 49372 4134
rect 55772 3664 55824 3670
rect 55772 3606 55824 3612
rect 50436 3596 50488 3602
rect 50436 3538 50488 3544
rect 49332 2916 49384 2922
rect 49332 2858 49384 2864
rect 50448 800 50476 3538
rect 55784 800 55812 3606
rect 55968 2786 55996 4134
rect 58636 4134 58972 4162
rect 55956 2780 56008 2786
rect 55956 2722 56008 2728
rect 58636 2446 58664 4134
rect 61108 3732 61160 3738
rect 61108 3674 61160 3680
rect 58624 2440 58676 2446
rect 58624 2382 58676 2388
rect 61120 800 61148 3674
rect 66180 2786 66208 4218
rect 68986 3890 69014 4148
rect 72312 4134 72648 4162
rect 79028 4134 79364 4162
rect 82340 4134 82676 4162
rect 85652 4134 85988 4162
rect 89056 4134 89392 4162
rect 68940 3862 69014 3890
rect 66444 3800 66496 3806
rect 66444 3742 66496 3748
rect 66168 2780 66220 2786
rect 66168 2722 66220 2728
rect 66456 800 66484 3742
rect 68940 2446 68968 3862
rect 68928 2440 68980 2446
rect 68928 2382 68980 2388
rect 72620 1358 72648 4134
rect 77024 3936 77076 3942
rect 77024 3878 77076 3884
rect 72608 1352 72660 1358
rect 72608 1294 72660 1300
rect 71608 870 71728 898
rect 34612 60 34664 66
rect 34612 2 34664 8
rect 39762 0 39818 800
rect 45098 0 45154 800
rect 50434 0 50490 800
rect 55770 0 55826 800
rect 61106 0 61162 800
rect 66442 0 66498 800
rect 71608 134 71636 870
rect 71700 800 71728 870
rect 77036 800 77064 3878
rect 79336 2378 79364 4134
rect 82360 3868 82412 3874
rect 82360 3810 82412 3816
rect 79324 2372 79376 2378
rect 79324 2314 79376 2320
rect 82372 800 82400 3810
rect 82648 1970 82676 4134
rect 85960 2786 85988 4134
rect 86868 4004 86920 4010
rect 86868 3946 86920 3952
rect 85948 2780 86000 2786
rect 85948 2722 86000 2728
rect 86880 2446 86908 3946
rect 87696 3324 87748 3330
rect 87696 3266 87748 3272
rect 86868 2440 86920 2446
rect 86868 2382 86920 2388
rect 82636 1964 82688 1970
rect 82636 1906 82688 1912
rect 87708 800 87736 3266
rect 89364 2242 89392 4134
rect 92354 3890 92382 4148
rect 95680 4134 96016 4162
rect 98992 4134 99328 4162
rect 102396 4134 102732 4162
rect 105708 4134 106044 4162
rect 92354 3862 92428 3890
rect 92400 2446 92428 3862
rect 93032 3392 93084 3398
rect 93032 3334 93084 3340
rect 92388 2440 92440 2446
rect 92388 2382 92440 2388
rect 89352 2236 89404 2242
rect 89352 2178 89404 2184
rect 93044 800 93072 3334
rect 95988 2174 96016 4134
rect 98368 3460 98420 3466
rect 98368 3402 98420 3408
rect 95976 2168 96028 2174
rect 95976 2110 96028 2116
rect 98380 800 98408 3402
rect 99300 2310 99328 4134
rect 99288 2304 99340 2310
rect 99288 2246 99340 2252
rect 102704 2106 102732 4134
rect 103612 2984 103664 2990
rect 103612 2926 103664 2932
rect 102692 2100 102744 2106
rect 102692 2042 102744 2048
rect 103624 800 103652 2926
rect 106016 1562 106044 4134
rect 109006 3890 109034 4148
rect 108960 3862 109034 3890
rect 108856 3528 108908 3534
rect 108856 3470 108908 3476
rect 108868 1850 108896 3470
rect 108960 2786 108988 3862
rect 108948 2780 109000 2786
rect 108948 2722 109000 2728
rect 113836 1902 113864 150583
rect 113928 3534 113956 151098
rect 114100 150340 114152 150346
rect 114100 150282 114152 150288
rect 114008 149388 114060 149394
rect 114008 149330 114060 149336
rect 114020 61674 114048 149330
rect 114112 71738 114140 150282
rect 114204 81394 114232 151710
rect 114284 151088 114336 151094
rect 114284 151030 114336 151036
rect 114296 133822 114324 151030
rect 115124 133890 115152 151846
rect 115664 151700 115716 151706
rect 115664 151642 115716 151648
rect 115202 150512 115258 150521
rect 115202 150447 115258 150456
rect 115112 133884 115164 133890
rect 115112 133826 115164 133832
rect 114284 133816 114336 133822
rect 114284 133758 114336 133764
rect 115112 94376 115164 94382
rect 115112 94318 115164 94324
rect 114192 81388 114244 81394
rect 114192 81330 114244 81336
rect 115124 79354 115152 94318
rect 115112 79348 115164 79354
rect 115112 79290 115164 79296
rect 114560 74588 114612 74594
rect 114560 74530 114612 74536
rect 114100 71732 114152 71738
rect 114100 71674 114152 71680
rect 114572 69018 114600 74530
rect 114560 69012 114612 69018
rect 114560 68954 114612 68960
rect 114008 61668 114060 61674
rect 114008 61610 114060 61616
rect 114008 55616 114060 55622
rect 114008 55558 114060 55564
rect 114020 5098 114048 55558
rect 114100 48272 114152 48278
rect 114100 48214 114152 48220
rect 114008 5092 114060 5098
rect 114008 5034 114060 5040
rect 114112 4758 114140 48214
rect 114192 44124 114244 44130
rect 114192 44066 114244 44072
rect 114100 4752 114152 4758
rect 114100 4694 114152 4700
rect 114204 4690 114232 44066
rect 114284 40044 114336 40050
rect 114284 39986 114336 39992
rect 114192 4684 114244 4690
rect 114192 4626 114244 4632
rect 114296 4622 114324 39986
rect 114560 37052 114612 37058
rect 114560 36994 114612 37000
rect 114572 31770 114600 36994
rect 114652 36236 114704 36242
rect 114652 36178 114704 36184
rect 114388 31742 114600 31770
rect 114388 5166 114416 31742
rect 114664 31634 114692 36178
rect 114480 31606 114692 31634
rect 114480 27674 114508 31606
rect 114468 27668 114520 27674
rect 114468 27610 114520 27616
rect 114468 27532 114520 27538
rect 114468 27474 114520 27480
rect 114480 5642 114508 27474
rect 115112 9716 115164 9722
rect 115112 9658 115164 9664
rect 114560 7200 114612 7206
rect 114560 7142 114612 7148
rect 114468 5636 114520 5642
rect 114468 5578 114520 5584
rect 114572 5302 114600 7142
rect 114560 5296 114612 5302
rect 114560 5238 114612 5244
rect 115124 5234 115152 9658
rect 115112 5228 115164 5234
rect 115112 5170 115164 5176
rect 114376 5160 114428 5166
rect 114376 5102 114428 5108
rect 114284 4616 114336 4622
rect 114284 4558 114336 4564
rect 114284 4004 114336 4010
rect 114284 3946 114336 3952
rect 113916 3528 113968 3534
rect 113916 3470 113968 3476
rect 113824 1896 113876 1902
rect 108868 1822 108988 1850
rect 113824 1838 113876 1844
rect 106004 1556 106056 1562
rect 106004 1498 106056 1504
rect 108960 800 108988 1822
rect 114296 800 114324 3946
rect 114652 3528 114704 3534
rect 114652 3470 114704 3476
rect 114560 2916 114612 2922
rect 114560 2858 114612 2864
rect 114572 2718 114600 2858
rect 114664 2718 114692 3470
rect 114560 2712 114612 2718
rect 114560 2654 114612 2660
rect 114652 2712 114704 2718
rect 114652 2654 114704 2660
rect 115216 2038 115244 150447
rect 115296 147688 115348 147694
rect 115296 147630 115348 147636
rect 115308 5438 115336 147630
rect 115388 142588 115440 142594
rect 115388 142530 115440 142536
rect 115296 5432 115348 5438
rect 115296 5374 115348 5380
rect 115400 2786 115428 142530
rect 115480 140820 115532 140826
rect 115480 140762 115532 140768
rect 115492 2922 115520 140762
rect 115572 138032 115624 138038
rect 115572 137974 115624 137980
rect 115480 2916 115532 2922
rect 115480 2858 115532 2864
rect 115388 2780 115440 2786
rect 115388 2722 115440 2728
rect 115204 2032 115256 2038
rect 115204 1974 115256 1980
rect 115584 1970 115612 137974
rect 115676 78674 115704 151642
rect 115768 88330 115796 152351
rect 117044 151836 117096 151842
rect 117044 151778 117096 151784
rect 116952 151360 117004 151366
rect 116952 151302 117004 151308
rect 116582 151192 116638 151201
rect 116582 151127 116638 151136
rect 116492 116000 116544 116006
rect 116492 115942 116544 115948
rect 115848 114028 115900 114034
rect 115848 113970 115900 113976
rect 115756 88324 115808 88330
rect 115756 88266 115808 88272
rect 115860 81870 115888 113970
rect 116504 89185 116532 115942
rect 116490 89176 116546 89185
rect 116490 89111 116546 89120
rect 115848 81864 115900 81870
rect 115848 81806 115900 81812
rect 115664 78668 115716 78674
rect 115664 78610 115716 78616
rect 116400 67584 116452 67590
rect 116400 67526 116452 67532
rect 116412 66473 116440 67526
rect 116398 66464 116454 66473
rect 116398 66399 116454 66408
rect 115664 52488 115716 52494
rect 115664 52430 115716 52436
rect 115676 5370 115704 52430
rect 115756 46164 115808 46170
rect 115756 46106 115808 46112
rect 115664 5364 115716 5370
rect 115664 5306 115716 5312
rect 115768 4554 115796 46106
rect 115848 16924 115900 16930
rect 115848 16866 115900 16872
rect 115860 4826 115888 16866
rect 116030 9616 116086 9625
rect 116030 9551 116086 9560
rect 116044 8362 116072 9551
rect 116032 8356 116084 8362
rect 116032 8298 116084 8304
rect 116596 6914 116624 151127
rect 116860 150544 116912 150550
rect 116860 150486 116912 150492
rect 116674 134736 116730 134745
rect 116674 134671 116730 134680
rect 116504 6886 116624 6914
rect 115848 4820 115900 4826
rect 115848 4762 115900 4768
rect 115756 4548 115808 4554
rect 115756 4490 115808 4496
rect 116504 1970 116532 6886
rect 116584 5364 116636 5370
rect 116584 5306 116636 5312
rect 115572 1964 115624 1970
rect 115572 1906 115624 1912
rect 116492 1964 116544 1970
rect 116492 1906 116544 1912
rect 116596 1834 116624 5306
rect 116688 5166 116716 134671
rect 116766 131200 116822 131209
rect 116766 131135 116822 131144
rect 116676 5160 116728 5166
rect 116676 5102 116728 5108
rect 116780 4350 116808 131135
rect 116872 121553 116900 150486
rect 116964 123321 116992 151302
rect 116950 123312 117006 123321
rect 116950 123247 117006 123256
rect 116858 121544 116914 121553
rect 116858 121479 116914 121488
rect 116858 112024 116914 112033
rect 116858 111959 116914 111968
rect 116872 5250 116900 111959
rect 116950 111752 117006 111761
rect 116950 111687 117006 111696
rect 116964 5370 116992 111687
rect 117056 82657 117084 151778
rect 117136 151020 117188 151026
rect 117136 150962 117188 150968
rect 117148 128761 117176 150962
rect 117792 150657 117820 153206
rect 118698 152416 118754 152425
rect 118698 152351 118754 152360
rect 118608 151564 118660 151570
rect 118608 151506 118660 151512
rect 118146 151328 118202 151337
rect 118146 151263 118202 151272
rect 118056 151224 118108 151230
rect 118056 151166 118108 151172
rect 117962 150784 118018 150793
rect 117962 150719 118018 150728
rect 117778 150648 117834 150657
rect 117778 150583 117834 150592
rect 117780 150476 117832 150482
rect 117780 150418 117832 150424
rect 117686 148200 117742 148209
rect 117686 148135 117742 148144
rect 117700 147694 117728 148135
rect 117688 147688 117740 147694
rect 117688 147630 117740 147636
rect 117320 146260 117372 146266
rect 117320 146202 117372 146208
rect 117226 146160 117282 146169
rect 117226 146095 117282 146104
rect 117134 128752 117190 128761
rect 117134 128687 117190 128696
rect 117134 106992 117190 107001
rect 117134 106927 117190 106936
rect 117042 82648 117098 82657
rect 117042 82583 117098 82592
rect 117148 43761 117176 106927
rect 117240 92449 117268 146095
rect 117332 145761 117360 146202
rect 117318 145752 117374 145761
rect 117318 145687 117374 145696
rect 117318 143304 117374 143313
rect 117318 143239 117374 143248
rect 117332 142594 117360 143239
rect 117320 142588 117372 142594
rect 117320 142530 117372 142536
rect 117318 140856 117374 140865
rect 117318 140791 117320 140800
rect 117372 140791 117374 140800
rect 117320 140762 117372 140768
rect 117686 138408 117742 138417
rect 117686 138343 117742 138352
rect 117700 138038 117728 138343
rect 117688 138032 117740 138038
rect 117688 137974 117740 137980
rect 117320 133816 117372 133822
rect 117320 133758 117372 133764
rect 117332 133657 117360 133758
rect 117318 133648 117374 133657
rect 117318 133583 117374 133592
rect 117502 116648 117558 116657
rect 117502 116583 117558 116592
rect 117516 116006 117544 116583
rect 117504 116000 117556 116006
rect 117504 115942 117556 115948
rect 117792 109313 117820 150418
rect 117872 133884 117924 133890
rect 117872 133826 117924 133832
rect 117778 109304 117834 109313
rect 117778 109239 117834 109248
rect 117318 102096 117374 102105
rect 117318 102031 117374 102040
rect 117332 100881 117360 102031
rect 117318 100872 117374 100881
rect 117318 100807 117374 100816
rect 117226 92440 117282 92449
rect 117226 92375 117282 92384
rect 117688 88324 117740 88330
rect 117688 88266 117740 88272
rect 117700 87553 117728 88266
rect 117686 87544 117742 87553
rect 117686 87479 117742 87488
rect 117884 85105 117912 133826
rect 117870 85096 117926 85105
rect 117870 85031 117926 85040
rect 117872 81864 117924 81870
rect 117872 81806 117924 81812
rect 117320 81388 117372 81394
rect 117320 81330 117372 81336
rect 117332 80209 117360 81330
rect 117318 80200 117374 80209
rect 117318 80135 117374 80144
rect 117780 79348 117832 79354
rect 117780 79290 117832 79296
rect 117688 78668 117740 78674
rect 117688 78610 117740 78616
rect 117700 77897 117728 78610
rect 117686 77888 117742 77897
rect 117686 77823 117742 77832
rect 117320 71732 117372 71738
rect 117320 71674 117372 71680
rect 117332 70553 117360 71674
rect 117318 70544 117374 70553
rect 117318 70479 117374 70488
rect 117320 69012 117372 69018
rect 117320 68954 117372 68960
rect 117332 68105 117360 68954
rect 117318 68096 117374 68105
rect 117318 68031 117374 68040
rect 117320 66224 117372 66230
rect 117320 66166 117372 66172
rect 117332 65657 117360 66166
rect 117318 65648 117374 65657
rect 117318 65583 117374 65592
rect 117320 61668 117372 61674
rect 117320 61610 117372 61616
rect 117332 58449 117360 61610
rect 117792 60897 117820 79290
rect 117884 63345 117912 81806
rect 117870 63336 117926 63345
rect 117870 63271 117926 63280
rect 117778 60888 117834 60897
rect 117778 60823 117834 60832
rect 117318 58440 117374 58449
rect 117318 58375 117374 58384
rect 117318 55992 117374 56001
rect 117318 55927 117374 55936
rect 117332 55622 117360 55927
rect 117320 55616 117372 55622
rect 117320 55558 117372 55564
rect 117318 53544 117374 53553
rect 117318 53479 117374 53488
rect 117332 52494 117360 53479
rect 117320 52488 117372 52494
rect 117320 52430 117372 52436
rect 117226 51096 117282 51105
rect 117226 51031 117282 51040
rect 117240 46170 117268 51031
rect 117318 48784 117374 48793
rect 117318 48719 117374 48728
rect 117332 48346 117360 48719
rect 117320 48340 117372 48346
rect 117320 48282 117372 48288
rect 117870 46336 117926 46345
rect 117870 46271 117926 46280
rect 117228 46164 117280 46170
rect 117228 46106 117280 46112
rect 117884 44198 117912 46271
rect 117872 44192 117924 44198
rect 117872 44134 117924 44140
rect 117226 43888 117282 43897
rect 117226 43823 117282 43832
rect 117134 43752 117190 43761
rect 117134 43687 117190 43696
rect 117240 37058 117268 43823
rect 117318 41440 117374 41449
rect 117318 41375 117374 41384
rect 117332 40118 117360 41375
rect 117320 40112 117372 40118
rect 117320 40054 117372 40060
rect 117318 38992 117374 39001
rect 117318 38927 117374 38936
rect 117332 38690 117360 38927
rect 117320 38684 117372 38690
rect 117320 38626 117372 38632
rect 117228 37052 117280 37058
rect 117228 36994 117280 37000
rect 117318 36544 117374 36553
rect 117318 36479 117374 36488
rect 117332 36242 117360 36479
rect 117320 36236 117372 36242
rect 117320 36178 117372 36184
rect 117042 32328 117098 32337
rect 117042 32263 117098 32272
rect 116952 5364 117004 5370
rect 116952 5306 117004 5312
rect 116872 5222 116992 5250
rect 116768 4344 116820 4350
rect 116768 4286 116820 4292
rect 116860 4072 116912 4078
rect 116860 4014 116912 4020
rect 116872 2786 116900 4014
rect 116964 3505 116992 5222
rect 117056 4078 117084 32263
rect 117320 31816 117372 31822
rect 117318 31784 117320 31793
rect 117372 31784 117374 31793
rect 117318 31719 117374 31728
rect 117318 29336 117374 29345
rect 117318 29271 117374 29280
rect 117332 29034 117360 29271
rect 117320 29028 117372 29034
rect 117320 28970 117372 28976
rect 117870 24440 117926 24449
rect 117870 24375 117926 24384
rect 117778 21992 117834 22001
rect 117778 21927 117834 21936
rect 117134 19680 117190 19689
rect 117134 19615 117190 19624
rect 117148 5778 117176 19615
rect 117502 17232 117558 17241
rect 117502 17167 117558 17176
rect 117516 16930 117544 17167
rect 117504 16924 117556 16930
rect 117504 16866 117556 16872
rect 117318 14784 117374 14793
rect 117318 14719 117374 14728
rect 117332 13870 117360 14719
rect 117320 13864 117372 13870
rect 117320 13806 117372 13812
rect 117226 12336 117282 12345
rect 117226 12271 117282 12280
rect 117136 5772 117188 5778
rect 117136 5714 117188 5720
rect 117240 5506 117268 12271
rect 117688 11756 117740 11762
rect 117688 11698 117740 11704
rect 117318 9888 117374 9897
rect 117318 9823 117374 9832
rect 117332 9722 117360 9823
rect 117320 9716 117372 9722
rect 117320 9658 117372 9664
rect 117318 7440 117374 7449
rect 117318 7375 117374 7384
rect 117332 7206 117360 7375
rect 117320 7200 117372 7206
rect 117320 7142 117372 7148
rect 117228 5500 117280 5506
rect 117228 5442 117280 5448
rect 117318 5128 117374 5137
rect 117318 5063 117374 5072
rect 117332 4214 117360 5063
rect 117320 4208 117372 4214
rect 117320 4150 117372 4156
rect 117044 4072 117096 4078
rect 117044 4014 117096 4020
rect 116950 3496 117006 3505
rect 116950 3431 117006 3440
rect 116860 2780 116912 2786
rect 116860 2722 116912 2728
rect 117700 1834 117728 11698
rect 117792 5710 117820 21927
rect 117884 5846 117912 24375
rect 117976 11762 118004 150719
rect 118068 136105 118096 151166
rect 118054 136096 118110 136105
rect 118054 136031 118110 136040
rect 118054 126304 118110 126313
rect 118054 126239 118110 126248
rect 117964 11756 118016 11762
rect 117964 11698 118016 11704
rect 117872 5840 117924 5846
rect 117872 5782 117924 5788
rect 117780 5704 117832 5710
rect 117780 5646 117832 5652
rect 118068 4282 118096 126239
rect 118056 4276 118108 4282
rect 118056 4218 118108 4224
rect 116584 1828 116636 1834
rect 116584 1770 116636 1776
rect 117688 1828 117740 1834
rect 117688 1770 117740 1776
rect 118160 1766 118188 151263
rect 118424 150272 118476 150278
rect 118424 150214 118476 150220
rect 118238 123856 118294 123865
rect 118238 123791 118294 123800
rect 118252 3534 118280 123791
rect 118330 119096 118386 119105
rect 118330 119031 118386 119040
rect 118344 4418 118372 119031
rect 118436 73001 118464 150214
rect 118514 149968 118570 149977
rect 118514 149903 118570 149912
rect 118528 75449 118556 149903
rect 118620 104553 118648 151506
rect 118712 114209 118740 152351
rect 119448 151814 119476 157354
rect 120078 154456 120134 154465
rect 120078 154391 120134 154400
rect 119526 152008 119582 152017
rect 120092 151994 120120 154391
rect 120368 152130 120396 159200
rect 120630 155272 120686 155281
rect 120630 155207 120686 155216
rect 120368 152102 120488 152130
rect 120092 151966 120336 151994
rect 119526 151943 119582 151952
rect 119356 151786 119476 151814
rect 118698 114200 118754 114209
rect 118698 114135 118754 114144
rect 118606 104544 118662 104553
rect 118606 104479 118662 104488
rect 118606 99648 118662 99657
rect 118606 99583 118662 99592
rect 118514 75440 118570 75449
rect 118514 75375 118570 75384
rect 118422 72992 118478 73001
rect 118422 72927 118478 72936
rect 118422 34232 118478 34241
rect 118422 34167 118478 34176
rect 118436 6089 118464 34167
rect 118514 26888 118570 26897
rect 118514 26823 118570 26832
rect 118422 6080 118478 6089
rect 118422 6015 118478 6024
rect 118528 5914 118556 26823
rect 118516 5908 118568 5914
rect 118516 5850 118568 5856
rect 118332 4412 118384 4418
rect 118332 4354 118384 4360
rect 118240 3528 118292 3534
rect 118240 3470 118292 3476
rect 118620 3369 118648 99583
rect 118698 97200 118754 97209
rect 118698 97135 118754 97144
rect 118712 4962 118740 97135
rect 118790 94752 118846 94761
rect 118790 94687 118846 94696
rect 118700 4956 118752 4962
rect 118700 4898 118752 4904
rect 118804 4826 118832 94687
rect 118882 89992 118938 90001
rect 118882 89927 118938 89936
rect 118896 5098 118924 89927
rect 118976 8356 119028 8362
rect 118976 8298 119028 8304
rect 118884 5092 118936 5098
rect 118884 5034 118936 5040
rect 118792 4820 118844 4826
rect 118792 4762 118844 4768
rect 118988 3534 119016 8298
rect 118976 3528 119028 3534
rect 118976 3470 119028 3476
rect 118606 3360 118662 3369
rect 118606 3295 118662 3304
rect 119356 2417 119384 151786
rect 119436 151088 119488 151094
rect 119436 151030 119488 151036
rect 119448 67590 119476 151030
rect 119436 67584 119488 67590
rect 119436 67526 119488 67532
rect 119540 2689 119568 151943
rect 120460 151910 120488 152102
rect 120644 151994 120672 155207
rect 121288 154737 121316 159200
rect 121918 156632 121974 156641
rect 121918 156567 121974 156576
rect 121458 155408 121514 155417
rect 121458 155343 121514 155352
rect 121274 154728 121330 154737
rect 121274 154663 121330 154672
rect 121472 154465 121500 155343
rect 121458 154456 121514 154465
rect 121458 154391 121514 154400
rect 121458 152552 121514 152561
rect 121458 152487 121514 152496
rect 121472 151994 121500 152487
rect 121932 151994 121960 156567
rect 122300 155417 122328 159200
rect 122840 158228 122892 158234
rect 122840 158170 122892 158176
rect 122286 155408 122342 155417
rect 122286 155343 122342 155352
rect 122852 151994 122880 158170
rect 123220 156641 123248 159200
rect 124232 156670 124260 159200
rect 123852 156664 123904 156670
rect 123206 156632 123262 156641
rect 123852 156606 123904 156612
rect 124220 156664 124272 156670
rect 124220 156606 124272 156612
rect 123206 156567 123262 156576
rect 123206 154456 123262 154465
rect 123206 154391 123262 154400
rect 123220 151994 123248 154391
rect 123864 151994 123892 156606
rect 125244 155446 125272 159200
rect 125232 155440 125284 155446
rect 125232 155382 125284 155388
rect 126164 155378 126192 159200
rect 127176 159174 127296 159200
rect 127072 158704 127124 158710
rect 127072 158646 127124 158652
rect 126428 156732 126480 156738
rect 126428 156674 126480 156680
rect 126060 155372 126112 155378
rect 126060 155314 126112 155320
rect 126152 155372 126204 155378
rect 126152 155314 126204 155320
rect 125048 155236 125100 155242
rect 125048 155178 125100 155184
rect 124496 152516 124548 152522
rect 124496 152458 124548 152464
rect 124508 151994 124536 152458
rect 125060 151994 125088 155178
rect 126072 153882 126100 155314
rect 125784 153876 125836 153882
rect 125784 153818 125836 153824
rect 126060 153876 126112 153882
rect 126060 153818 126112 153824
rect 125796 151994 125824 153818
rect 126440 151994 126468 156674
rect 127084 151994 127112 158646
rect 127452 152130 127480 159310
rect 128082 159200 128138 160000
rect 129094 159200 129150 160000
rect 130106 159200 130162 160000
rect 131026 159200 131082 160000
rect 132038 159200 132094 160000
rect 132958 159200 133014 160000
rect 133970 159200 134026 160000
rect 134982 159200 135038 160000
rect 135902 159200 135958 160000
rect 136914 159200 136970 160000
rect 137834 159200 137890 160000
rect 138846 159200 138902 160000
rect 139858 159200 139914 160000
rect 140778 159200 140834 160000
rect 141790 159200 141846 160000
rect 142710 159200 142766 160000
rect 143722 159200 143778 160000
rect 144734 159200 144790 160000
rect 145654 159200 145710 160000
rect 146666 159200 146722 160000
rect 147586 159200 147642 160000
rect 148598 159200 148654 160000
rect 149610 159200 149666 160000
rect 150530 159200 150586 160000
rect 151542 159200 151598 160000
rect 152462 159200 152518 160000
rect 153474 159200 153530 160000
rect 154486 159200 154542 160000
rect 155406 159200 155462 160000
rect 156418 159200 156474 160000
rect 157338 159200 157394 160000
rect 158350 159200 158406 160000
rect 159270 159200 159326 160000
rect 160282 159200 160338 160000
rect 161294 159200 161350 160000
rect 162214 159200 162270 160000
rect 163226 159200 163282 160000
rect 164146 159200 164202 160000
rect 165158 159200 165214 160000
rect 166170 159200 166226 160000
rect 167090 159200 167146 160000
rect 168102 159200 168158 160000
rect 169022 159200 169078 160000
rect 170034 159200 170090 160000
rect 171046 159200 171102 160000
rect 171966 159200 172022 160000
rect 172978 159200 173034 160000
rect 173898 159200 173954 160000
rect 174910 159202 174966 160000
rect 175016 159310 175228 159338
rect 175016 159202 175044 159310
rect 174910 159200 175044 159202
rect 127898 156088 127954 156097
rect 127898 156023 127954 156032
rect 127452 152102 127572 152130
rect 120644 151966 120980 151994
rect 121472 151966 121624 151994
rect 121932 151966 122268 151994
rect 122852 151966 122912 151994
rect 123220 151966 123556 151994
rect 123864 151966 124200 151994
rect 124508 151966 124844 151994
rect 125060 151966 125488 151994
rect 125796 151966 126132 151994
rect 126440 151966 126776 151994
rect 127084 151966 127420 151994
rect 120448 151904 120500 151910
rect 120448 151846 120500 151852
rect 127544 151842 127572 152102
rect 127912 151994 127940 156023
rect 128096 152561 128124 159200
rect 129108 157622 129136 159200
rect 129740 158840 129792 158846
rect 129740 158782 129792 158788
rect 129096 157616 129148 157622
rect 129096 157558 129148 157564
rect 128360 153944 128412 153950
rect 128360 153886 128412 153892
rect 128082 152552 128138 152561
rect 128082 152487 128138 152496
rect 128372 151994 128400 153886
rect 129004 152924 129056 152930
rect 129004 152866 129056 152872
rect 129016 151994 129044 152866
rect 129752 151994 129780 158782
rect 130120 153882 130148 159200
rect 131040 157185 131068 159200
rect 131026 157176 131082 157185
rect 131026 157111 131082 157120
rect 131672 156800 131724 156806
rect 131672 156742 131724 156748
rect 131118 154320 131174 154329
rect 131118 154255 131174 154264
rect 130108 153876 130160 153882
rect 130108 153818 130160 153824
rect 130384 153264 130436 153270
rect 130384 153206 130436 153212
rect 130396 151994 130424 153206
rect 131132 151994 131160 154255
rect 131684 151994 131712 156742
rect 132052 156738 132080 159200
rect 132592 158160 132644 158166
rect 132592 158102 132644 158108
rect 132040 156732 132092 156738
rect 132040 156674 132092 156680
rect 132604 151994 132632 158102
rect 132972 155514 133000 159200
rect 132960 155508 133012 155514
rect 132960 155450 133012 155456
rect 133984 155378 134012 159200
rect 134892 158772 134944 158778
rect 134892 158714 134944 158720
rect 133788 155372 133840 155378
rect 133788 155314 133840 155320
rect 133972 155372 134024 155378
rect 133972 155314 134024 155320
rect 133800 153270 133828 155314
rect 133880 154012 133932 154018
rect 133880 153954 133932 153960
rect 132960 153264 133012 153270
rect 132960 153206 133012 153212
rect 133788 153264 133840 153270
rect 133788 153206 133840 153212
rect 132972 151994 133000 153206
rect 133892 151994 133920 153954
rect 134248 152584 134300 152590
rect 134248 152526 134300 152532
rect 134260 151994 134288 152526
rect 134904 151994 134932 158714
rect 134996 156806 135024 159200
rect 134984 156800 135036 156806
rect 134984 156742 135036 156748
rect 135168 155440 135220 155446
rect 135168 155382 135220 155388
rect 135180 154018 135208 155382
rect 135168 154012 135220 154018
rect 135168 153954 135220 153960
rect 135536 153944 135588 153950
rect 135536 153886 135588 153892
rect 135548 151994 135576 153886
rect 135916 152522 135944 159200
rect 136824 156868 136876 156874
rect 136824 156810 136876 156816
rect 136178 155544 136234 155553
rect 136178 155479 136234 155488
rect 135904 152516 135956 152522
rect 135904 152458 135956 152464
rect 136192 151994 136220 155479
rect 136732 155236 136784 155242
rect 136732 155178 136784 155184
rect 136744 153950 136772 155178
rect 136732 153944 136784 153950
rect 136732 153886 136784 153892
rect 136836 151994 136864 156810
rect 136928 155786 136956 159200
rect 137468 158908 137520 158914
rect 137468 158850 137520 158856
rect 136916 155780 136968 155786
rect 136916 155722 136968 155728
rect 137480 151994 137508 158850
rect 137848 155514 137876 159200
rect 137836 155508 137888 155514
rect 137836 155450 137888 155456
rect 138020 155304 138072 155310
rect 138020 155246 138072 155252
rect 138032 154018 138060 155246
rect 138860 154170 138888 159200
rect 139872 156874 139900 159200
rect 140792 157690 140820 159200
rect 140136 157684 140188 157690
rect 140136 157626 140188 157632
rect 140780 157684 140832 157690
rect 140780 157626 140832 157632
rect 139860 156868 139912 156874
rect 139860 156810 139912 156816
rect 138860 154142 138980 154170
rect 138848 154080 138900 154086
rect 138848 154022 138900 154028
rect 138020 154012 138072 154018
rect 138020 153954 138072 153960
rect 138112 153264 138164 153270
rect 138112 153206 138164 153212
rect 138124 151994 138152 153206
rect 138860 151994 138888 154022
rect 138952 152590 138980 154142
rect 139492 152652 139544 152658
rect 139492 152594 139544 152600
rect 138940 152584 138992 152590
rect 138940 152526 138992 152532
rect 139504 151994 139532 152594
rect 140148 151994 140176 157626
rect 140870 155680 140926 155689
rect 140870 155615 140926 155624
rect 140780 155236 140832 155242
rect 140780 155178 140832 155184
rect 140792 154086 140820 155178
rect 140780 154080 140832 154086
rect 140780 154022 140832 154028
rect 140884 153950 140912 155615
rect 141804 155310 141832 159200
rect 142250 156224 142306 156233
rect 142250 156159 142306 156168
rect 141792 155304 141844 155310
rect 141792 155246 141844 155252
rect 141424 154148 141476 154154
rect 141424 154090 141476 154096
rect 140780 153944 140832 153950
rect 140780 153886 140832 153892
rect 140872 153944 140924 153950
rect 140872 153886 140924 153892
rect 140792 151994 140820 153886
rect 141436 151994 141464 154090
rect 142264 151994 142292 156159
rect 142724 152930 142752 159200
rect 142804 158296 142856 158302
rect 142804 158238 142856 158244
rect 142712 152924 142764 152930
rect 142712 152866 142764 152872
rect 142816 151994 142844 158238
rect 143736 155786 143764 159200
rect 144748 155786 144776 159200
rect 145288 157752 145340 157758
rect 145288 157694 145340 157700
rect 143724 155780 143776 155786
rect 143724 155722 143776 155728
rect 144644 155780 144696 155786
rect 144644 155722 144696 155728
rect 144736 155780 144788 155786
rect 144736 155722 144788 155728
rect 144656 155530 144684 155722
rect 144656 155502 144868 155530
rect 144840 155446 144868 155502
rect 144736 155440 144788 155446
rect 144736 155382 144788 155388
rect 144828 155440 144880 155446
rect 144828 155382 144880 155388
rect 144748 154222 144776 155382
rect 144828 154896 144880 154902
rect 144828 154838 144880 154844
rect 143540 154216 143592 154222
rect 143540 154158 143592 154164
rect 144736 154216 144788 154222
rect 144736 154158 144788 154164
rect 143552 151994 143580 154158
rect 144840 154154 144868 154838
rect 144828 154148 144880 154154
rect 144828 154090 144880 154096
rect 144000 153944 144052 153950
rect 144000 153886 144052 153892
rect 144012 151994 144040 153886
rect 144918 152688 144974 152697
rect 144918 152623 144974 152632
rect 144932 151994 144960 152623
rect 145300 151994 145328 157694
rect 145668 153950 145696 159200
rect 146576 154284 146628 154290
rect 146576 154226 146628 154232
rect 145932 154012 145984 154018
rect 145932 153954 145984 153960
rect 145656 153944 145708 153950
rect 145656 153886 145708 153892
rect 145944 151994 145972 153954
rect 146588 151994 146616 154226
rect 146680 152658 146708 159200
rect 147600 155514 147628 159200
rect 148612 157758 148640 159200
rect 148692 158364 148744 158370
rect 148692 158306 148744 158312
rect 148600 157752 148652 157758
rect 148600 157694 148652 157700
rect 147956 156936 148008 156942
rect 147956 156878 148008 156884
rect 147588 155508 147640 155514
rect 147588 155450 147640 155456
rect 146760 155440 146812 155446
rect 146760 155382 146812 155388
rect 146772 155281 146800 155382
rect 146758 155272 146814 155281
rect 146758 155207 146814 155216
rect 147220 152720 147272 152726
rect 147220 152662 147272 152668
rect 146668 152652 146720 152658
rect 146668 152594 146720 152600
rect 147232 151994 147260 152662
rect 147968 151994 147996 156878
rect 148704 151994 148732 158306
rect 149624 155786 149652 159200
rect 150544 156942 150572 159200
rect 151176 157820 151228 157826
rect 151176 157762 151228 157768
rect 150532 156936 150584 156942
rect 150532 156878 150584 156884
rect 149612 155780 149664 155786
rect 149612 155722 149664 155728
rect 149150 155272 149206 155281
rect 149150 155207 149206 155216
rect 149058 154592 149114 154601
rect 149058 154527 149114 154536
rect 149072 154290 149100 154527
rect 149060 154284 149112 154290
rect 149060 154226 149112 154232
rect 149164 152930 149192 155207
rect 149244 154352 149296 154358
rect 149244 154294 149296 154300
rect 149152 152924 149204 152930
rect 149152 152866 149204 152872
rect 149256 151994 149284 154294
rect 149888 152856 149940 152862
rect 149888 152798 149940 152804
rect 149900 151994 149928 152798
rect 150532 152788 150584 152794
rect 150532 152730 150584 152736
rect 150544 151994 150572 152730
rect 151188 151994 151216 157762
rect 151556 152794 151584 159200
rect 152476 157321 152504 159200
rect 152462 157312 152518 157321
rect 152462 157247 152518 157256
rect 153198 156768 153254 156777
rect 153198 156703 153254 156712
rect 153108 155780 153160 155786
rect 153108 155722 153160 155728
rect 152004 154420 152056 154426
rect 152004 154362 152056 154368
rect 151544 152788 151596 152794
rect 151544 152730 151596 152736
rect 152016 151994 152044 154362
rect 153120 154018 153148 155722
rect 153108 154012 153160 154018
rect 153108 153954 153160 153960
rect 152464 152992 152516 152998
rect 152464 152934 152516 152940
rect 152476 151994 152504 152934
rect 153212 151994 153240 156703
rect 153488 155786 153516 159200
rect 153752 158432 153804 158438
rect 153752 158374 153804 158380
rect 153476 155780 153528 155786
rect 153476 155722 153528 155728
rect 153764 151994 153792 158374
rect 154500 152862 154528 159200
rect 155040 157004 155092 157010
rect 155040 156946 155092 156952
rect 154578 155816 154634 155825
rect 154578 155751 154634 155760
rect 154488 152856 154540 152862
rect 154488 152798 154540 152804
rect 154592 151994 154620 155751
rect 155052 151994 155080 156946
rect 155420 155786 155448 159200
rect 156328 158568 156380 158574
rect 156328 158510 156380 158516
rect 155868 155984 155920 155990
rect 155868 155926 155920 155932
rect 155408 155780 155460 155786
rect 155408 155722 155460 155728
rect 155880 155514 155908 155926
rect 155868 155508 155920 155514
rect 155868 155450 155920 155456
rect 155960 153060 156012 153066
rect 155960 153002 156012 153008
rect 155972 151994 156000 153002
rect 156340 151994 156368 158510
rect 156432 153066 156460 159200
rect 157352 154086 157380 159200
rect 157708 157072 157760 157078
rect 157708 157014 157760 157020
rect 156972 154080 157024 154086
rect 156972 154022 157024 154028
rect 157340 154080 157392 154086
rect 157340 154022 157392 154028
rect 156420 153060 156472 153066
rect 156420 153002 156472 153008
rect 156984 151994 157012 154022
rect 157720 151994 157748 157014
rect 158364 157010 158392 159200
rect 158996 157888 159048 157894
rect 158996 157830 159048 157836
rect 158444 157140 158496 157146
rect 158444 157082 158496 157088
rect 158352 157004 158404 157010
rect 158352 156946 158404 156952
rect 158456 151994 158484 157082
rect 158720 155508 158772 155514
rect 158720 155450 158772 155456
rect 158732 154494 158760 155450
rect 158720 154488 158772 154494
rect 158720 154430 158772 154436
rect 159008 151994 159036 157830
rect 159284 155514 159312 159200
rect 160100 157072 160152 157078
rect 160100 157014 160152 157020
rect 160112 155786 160140 157014
rect 160296 155786 160324 159200
rect 160100 155780 160152 155786
rect 160100 155722 160152 155728
rect 160284 155780 160336 155786
rect 160284 155722 160336 155728
rect 159272 155508 159324 155514
rect 159272 155450 159324 155456
rect 161308 155281 161336 159200
rect 161664 158500 161716 158506
rect 161664 158442 161716 158448
rect 161294 155272 161350 155281
rect 161294 155207 161350 155216
rect 159640 154420 159692 154426
rect 159640 154362 159692 154368
rect 159652 151994 159680 154362
rect 160284 153128 160336 153134
rect 160284 153070 160336 153076
rect 160296 151994 160324 153070
rect 160928 152448 160980 152454
rect 160928 152390 160980 152396
rect 160940 151994 160968 152390
rect 161676 151994 161704 158442
rect 162124 155440 162176 155446
rect 162124 155382 162176 155388
rect 162136 154222 162164 155382
rect 162228 155122 162256 159200
rect 163044 157140 163096 157146
rect 163044 157082 163096 157088
rect 162858 156904 162914 156913
rect 162858 156839 162914 156848
rect 162228 155094 162348 155122
rect 161848 154216 161900 154222
rect 161848 154158 161900 154164
rect 162124 154216 162176 154222
rect 162124 154158 162176 154164
rect 161860 152130 161888 154158
rect 162320 153134 162348 155094
rect 162308 153128 162360 153134
rect 162308 153070 162360 153076
rect 161860 152102 162164 152130
rect 162136 151994 162164 152102
rect 162872 151994 162900 156839
rect 163056 155514 163084 157082
rect 163044 155508 163096 155514
rect 163044 155450 163096 155456
rect 163240 155446 163268 159200
rect 163504 157208 163556 157214
rect 163504 157150 163556 157156
rect 163228 155440 163280 155446
rect 163228 155382 163280 155388
rect 163516 151994 163544 157150
rect 164160 155514 164188 159200
rect 164240 158636 164292 158642
rect 164240 158578 164292 158584
rect 164148 155508 164200 155514
rect 164148 155450 164200 155456
rect 164252 151994 164280 158578
rect 165172 154766 165200 159200
rect 165620 157276 165672 157282
rect 165620 157218 165672 157224
rect 165528 155440 165580 155446
rect 165528 155382 165580 155388
rect 164884 154760 164936 154766
rect 164884 154702 164936 154708
rect 165160 154760 165212 154766
rect 165160 154702 165212 154708
rect 164792 154556 164844 154562
rect 164792 154498 164844 154504
rect 164804 151994 164832 154498
rect 164896 154358 164924 154702
rect 164884 154352 164936 154358
rect 164884 154294 164936 154300
rect 165540 152454 165568 155382
rect 165528 152448 165580 152454
rect 165528 152390 165580 152396
rect 165632 151994 165660 157218
rect 166184 157078 166212 159200
rect 167104 157214 167132 159200
rect 167092 157208 167144 157214
rect 167092 157150 167144 157156
rect 166172 157072 166224 157078
rect 166172 157014 166224 157020
rect 167736 155712 167788 155718
rect 167736 155654 167788 155660
rect 167460 154284 167512 154290
rect 167460 154226 167512 154232
rect 167000 154148 167052 154154
rect 167000 154090 167052 154096
rect 166080 152380 166132 152386
rect 166080 152322 166132 152328
rect 166092 151994 166120 152322
rect 167012 151994 167040 154090
rect 167472 151994 167500 154226
rect 167748 153746 167776 155654
rect 167736 153740 167788 153746
rect 167736 153682 167788 153688
rect 168116 153134 168144 159200
rect 168748 157344 168800 157350
rect 168748 157286 168800 157292
rect 168380 155168 168432 155174
rect 168380 155110 168432 155116
rect 168392 154290 168420 155110
rect 168380 154284 168432 154290
rect 168380 154226 168432 154232
rect 168380 153196 168432 153202
rect 168380 153138 168432 153144
rect 168104 153128 168156 153134
rect 168104 153070 168156 153076
rect 168392 151994 168420 153138
rect 168760 151994 168788 157286
rect 169036 155174 169064 159200
rect 169024 155168 169076 155174
rect 169024 155110 169076 155116
rect 169392 153740 169444 153746
rect 169392 153682 169444 153688
rect 169404 151994 169432 153682
rect 170048 153202 170076 159200
rect 170680 157276 170732 157282
rect 170680 157218 170732 157224
rect 170126 155952 170182 155961
rect 170126 155887 170182 155896
rect 170036 153196 170088 153202
rect 170036 153138 170088 153144
rect 170140 151994 170168 155887
rect 170692 151994 170720 157218
rect 171060 155718 171088 159200
rect 171980 155718 172008 159200
rect 172152 155780 172204 155786
rect 172204 155740 172560 155768
rect 172152 155722 172204 155728
rect 171048 155712 171100 155718
rect 171048 155654 171100 155660
rect 171968 155712 172020 155718
rect 171968 155654 172020 155660
rect 172428 155168 172480 155174
rect 172428 155110 172480 155116
rect 171968 154420 172020 154426
rect 171968 154362 172020 154368
rect 171416 152312 171468 152318
rect 171416 152254 171468 152260
rect 171428 151994 171456 152254
rect 171980 151994 172008 154362
rect 172440 154154 172468 155110
rect 172428 154148 172480 154154
rect 172428 154090 172480 154096
rect 172532 152386 172560 155740
rect 172992 155174 173020 159200
rect 173912 157146 173940 159200
rect 174924 159174 175044 159200
rect 174544 157956 174596 157962
rect 174544 157898 174596 157904
rect 173900 157140 173952 157146
rect 173900 157082 173952 157088
rect 173716 156460 173768 156466
rect 173716 156402 173768 156408
rect 173728 156346 173756 156402
rect 173728 156318 173940 156346
rect 172980 155168 173032 155174
rect 172980 155110 173032 155116
rect 172612 153808 172664 153814
rect 172612 153750 172664 153756
rect 172520 152380 172572 152386
rect 172520 152322 172572 152328
rect 172624 151994 172652 153750
rect 173578 152244 173630 152250
rect 173578 152186 173630 152192
rect 127912 151966 128064 151994
rect 128372 151966 128708 151994
rect 129016 151966 129352 151994
rect 129752 151966 130088 151994
rect 130396 151966 130732 151994
rect 131132 151966 131376 151994
rect 131684 151966 132020 151994
rect 132604 151966 132664 151994
rect 132972 151966 133308 151994
rect 133892 151966 133952 151994
rect 134260 151966 134596 151994
rect 134904 151966 135240 151994
rect 135548 151966 135884 151994
rect 136192 151966 136528 151994
rect 136836 151966 137172 151994
rect 137480 151966 137816 151994
rect 138124 151966 138460 151994
rect 138860 151966 139196 151994
rect 139504 151966 139840 151994
rect 140148 151966 140484 151994
rect 140792 151966 141128 151994
rect 141436 151966 141772 151994
rect 142264 151966 142416 151994
rect 142816 151966 143060 151994
rect 143552 151966 143704 151994
rect 144012 151966 144348 151994
rect 144932 151966 144992 151994
rect 145300 151966 145636 151994
rect 145944 151966 146280 151994
rect 146588 151966 146924 151994
rect 147232 151966 147568 151994
rect 147968 151966 148304 151994
rect 148704 151966 148948 151994
rect 149256 151966 149592 151994
rect 149900 151966 150236 151994
rect 150544 151966 150880 151994
rect 151188 151966 151524 151994
rect 152016 151966 152168 151994
rect 152476 151966 152812 151994
rect 153212 151966 153456 151994
rect 153764 151966 154100 151994
rect 154592 151966 154744 151994
rect 155052 151966 155388 151994
rect 155972 151966 156032 151994
rect 156340 151966 156676 151994
rect 156984 151966 157320 151994
rect 157720 151966 158056 151994
rect 158456 151966 158700 151994
rect 159008 151966 159344 151994
rect 159652 151966 159988 151994
rect 160296 151966 160632 151994
rect 160940 151966 161276 151994
rect 161676 151966 161920 151994
rect 162136 151966 162564 151994
rect 162872 151966 163208 151994
rect 163516 151966 163852 151994
rect 164252 151966 164496 151994
rect 164804 151966 165140 151994
rect 165632 151966 165784 151994
rect 166092 151966 166428 151994
rect 167012 151966 167164 151994
rect 167472 151966 167808 151994
rect 168392 151966 168452 151994
rect 168760 151966 169096 151994
rect 169404 151966 169740 151994
rect 170140 151966 170384 151994
rect 170692 151966 171028 151994
rect 171428 151966 171672 151994
rect 171980 151966 172316 151994
rect 172624 151966 172960 151994
rect 173590 151980 173618 152186
rect 173912 151994 173940 156318
rect 174556 151994 174584 157898
rect 175200 154578 175228 159310
rect 175922 159200 175978 160000
rect 176842 159200 176898 160000
rect 177854 159200 177910 160000
rect 178774 159200 178830 160000
rect 179786 159200 179842 160000
rect 180798 159200 180854 160000
rect 181718 159200 181774 160000
rect 182730 159200 182786 160000
rect 183650 159200 183706 160000
rect 184662 159200 184718 160000
rect 185674 159200 185730 160000
rect 186594 159200 186650 160000
rect 187606 159200 187662 160000
rect 188526 159200 188582 160000
rect 189538 159200 189594 160000
rect 190550 159200 190606 160000
rect 191470 159200 191526 160000
rect 192482 159200 192538 160000
rect 193402 159200 193458 160000
rect 194414 159200 194470 160000
rect 195334 159200 195390 160000
rect 196346 159200 196402 160000
rect 197358 159200 197414 160000
rect 198278 159200 198334 160000
rect 199290 159200 199346 160000
rect 200210 159200 200266 160000
rect 201222 159200 201278 160000
rect 202234 159200 202290 160000
rect 203154 159200 203210 160000
rect 204166 159200 204222 160000
rect 205086 159200 205142 160000
rect 206098 159200 206154 160000
rect 207110 159200 207166 160000
rect 208030 159200 208086 160000
rect 209042 159200 209098 160000
rect 209962 159200 210018 160000
rect 210974 159200 211030 160000
rect 211986 159200 212042 160000
rect 212906 159200 212962 160000
rect 213918 159200 213974 160000
rect 214838 159200 214894 160000
rect 215850 159200 215906 160000
rect 216862 159200 216918 160000
rect 217782 159200 217838 160000
rect 218794 159200 218850 160000
rect 219714 159200 219770 160000
rect 220726 159200 220782 160000
rect 221738 159200 221794 160000
rect 222658 159200 222714 160000
rect 223670 159200 223726 160000
rect 224590 159200 224646 160000
rect 225602 159200 225658 160000
rect 226614 159200 226670 160000
rect 227534 159200 227590 160000
rect 228546 159200 228602 160000
rect 229466 159200 229522 160000
rect 230478 159200 230534 160000
rect 231490 159200 231546 160000
rect 232410 159200 232466 160000
rect 233422 159200 233478 160000
rect 234342 159200 234398 160000
rect 235354 159200 235410 160000
rect 236274 159200 236330 160000
rect 237286 159200 237342 160000
rect 238298 159200 238354 160000
rect 239218 159200 239274 160000
rect 240230 159200 240286 160000
rect 241150 159200 241206 160000
rect 242162 159200 242218 160000
rect 243174 159200 243230 160000
rect 244094 159200 244150 160000
rect 245106 159200 245162 160000
rect 246026 159200 246082 160000
rect 247038 159200 247094 160000
rect 248050 159200 248106 160000
rect 248970 159200 249026 160000
rect 249982 159200 250038 160000
rect 250902 159200 250958 160000
rect 251914 159200 251970 160000
rect 252926 159202 252982 160000
rect 253032 159310 253244 159338
rect 253032 159202 253060 159310
rect 252926 159200 253060 159202
rect 175936 157282 175964 159200
rect 175924 157276 175976 157282
rect 175924 157218 175976 157224
rect 176016 157208 176068 157214
rect 176016 157150 176068 157156
rect 175280 154624 175332 154630
rect 175200 154572 175280 154578
rect 175200 154566 175332 154572
rect 175200 154550 175320 154566
rect 175280 154420 175332 154426
rect 175280 154362 175332 154368
rect 175292 151994 175320 154362
rect 176028 151994 176056 157150
rect 176856 155922 176884 159200
rect 177868 157214 177896 159200
rect 177856 157208 177908 157214
rect 177856 157150 177908 157156
rect 178788 156398 178816 159200
rect 179602 157040 179658 157049
rect 179602 156975 179658 156984
rect 178776 156392 178828 156398
rect 178776 156334 178828 156340
rect 176844 155916 176896 155922
rect 176844 155858 176896 155864
rect 179144 155916 179196 155922
rect 179144 155858 179196 155864
rect 179156 154222 179184 155858
rect 179418 154864 179474 154873
rect 179418 154799 179474 154808
rect 179432 154562 179460 154799
rect 179512 154760 179564 154766
rect 179512 154702 179564 154708
rect 179420 154556 179472 154562
rect 179420 154498 179472 154504
rect 178040 154216 178092 154222
rect 178040 154158 178092 154164
rect 179144 154216 179196 154222
rect 179144 154158 179196 154164
rect 176890 152176 176942 152182
rect 176890 152118 176942 152124
rect 173912 151966 174248 151994
rect 174556 151966 174892 151994
rect 175292 151966 175536 151994
rect 176028 151966 176272 151994
rect 176902 151980 176930 152118
rect 178052 151994 178080 154158
rect 179524 153814 179552 154702
rect 179512 153808 179564 153814
rect 179512 153750 179564 153756
rect 178822 152108 178874 152114
rect 178822 152050 178874 152056
rect 178052 151966 178204 151994
rect 178834 151980 178862 152050
rect 179616 151994 179644 156975
rect 179800 154766 179828 159200
rect 180812 155922 180840 159200
rect 181076 157344 181128 157350
rect 181076 157286 181128 157292
rect 180892 156392 180944 156398
rect 180892 156334 180944 156340
rect 180904 156262 180932 156334
rect 180892 156256 180944 156262
rect 180892 156198 180944 156204
rect 180800 155916 180852 155922
rect 180800 155858 180852 155864
rect 180430 155136 180486 155145
rect 180430 155071 180486 155080
rect 179788 154760 179840 154766
rect 179788 154702 179840 154708
rect 179788 154284 179840 154290
rect 179788 154226 179840 154232
rect 179492 151966 179644 151994
rect 179800 151994 179828 154226
rect 180444 151994 180472 155071
rect 181088 151994 181116 157286
rect 181732 153762 181760 159200
rect 182364 158024 182416 158030
rect 182364 157966 182416 157972
rect 182088 155032 182140 155038
rect 182088 154974 182140 154980
rect 181732 153734 181852 153762
rect 181720 153604 181772 153610
rect 181720 153546 181772 153552
rect 181732 151994 181760 153546
rect 181824 152318 181852 153734
rect 182100 153610 182128 154974
rect 182088 153604 182140 153610
rect 182088 153546 182140 153552
rect 181812 152312 181864 152318
rect 181812 152254 181864 152260
rect 182376 151994 182404 157966
rect 182744 155650 182772 159200
rect 183468 156256 183520 156262
rect 183468 156198 183520 156204
rect 183376 155916 183428 155922
rect 183376 155858 183428 155864
rect 182732 155644 182784 155650
rect 182732 155586 182784 155592
rect 183388 154290 183416 155858
rect 183480 154630 183508 156198
rect 183664 154630 183692 159200
rect 184676 154698 184704 159200
rect 185688 155122 185716 159200
rect 186504 156324 186556 156330
rect 186504 156266 186556 156272
rect 186412 155916 186464 155922
rect 186412 155858 186464 155864
rect 186318 155408 186374 155417
rect 186318 155343 186374 155352
rect 185688 155094 185808 155122
rect 185492 155032 185544 155038
rect 185544 154980 185716 154986
rect 185492 154974 185716 154980
rect 185504 154958 185716 154974
rect 185584 154828 185636 154834
rect 185584 154770 185636 154776
rect 184296 154692 184348 154698
rect 184296 154634 184348 154640
rect 184664 154692 184716 154698
rect 184664 154634 184716 154640
rect 183468 154624 183520 154630
rect 183468 154566 183520 154572
rect 183652 154624 183704 154630
rect 183652 154566 183704 154572
rect 184308 154494 184336 154634
rect 184940 154556 184992 154562
rect 184940 154498 184992 154504
rect 184296 154488 184348 154494
rect 184296 154430 184348 154436
rect 183376 154284 183428 154290
rect 183376 154226 183428 154232
rect 183008 153740 183060 153746
rect 183008 153682 183060 153688
rect 183020 151994 183048 153682
rect 184296 153264 184348 153270
rect 184296 153206 184348 153212
rect 183652 152040 183704 152046
rect 179800 151966 180136 151994
rect 180444 151966 180780 151994
rect 181088 151966 181424 151994
rect 181732 151966 182068 151994
rect 182376 151966 182712 151994
rect 183020 151966 183356 151994
rect 184308 151994 184336 153206
rect 184952 151994 184980 154498
rect 185596 153746 185624 154770
rect 185688 154766 185716 154958
rect 185676 154760 185728 154766
rect 185676 154702 185728 154708
rect 185676 154352 185728 154358
rect 185676 154294 185728 154300
rect 185584 153740 185636 153746
rect 185584 153682 185636 153688
rect 185688 151994 185716 154294
rect 185780 152250 185808 155094
rect 186332 154562 186360 155343
rect 186320 154556 186372 154562
rect 186320 154498 186372 154504
rect 186424 154358 186452 155858
rect 186412 154352 186464 154358
rect 186412 154294 186464 154300
rect 185768 152244 185820 152250
rect 185768 152186 185820 152192
rect 186516 151994 186544 156266
rect 186608 155922 186636 159200
rect 186596 155916 186648 155922
rect 186596 155858 186648 155864
rect 186964 153536 187016 153542
rect 186964 153478 187016 153484
rect 186976 151994 187004 153478
rect 187620 152182 187648 159200
rect 187792 155576 187844 155582
rect 187792 155518 187844 155524
rect 187700 155100 187752 155106
rect 187700 155042 187752 155048
rect 187712 153814 187740 155042
rect 187700 153808 187752 153814
rect 187700 153750 187752 153756
rect 187700 153672 187752 153678
rect 187700 153614 187752 153620
rect 187608 152176 187660 152182
rect 187608 152118 187660 152124
rect 187712 151994 187740 153614
rect 187804 152114 187832 155518
rect 188540 155106 188568 159200
rect 189552 157350 189580 159200
rect 189632 157480 189684 157486
rect 189632 157422 189684 157428
rect 189540 157344 189592 157350
rect 189540 157286 189592 157292
rect 188528 155100 188580 155106
rect 188528 155042 188580 155048
rect 189080 154760 189132 154766
rect 189080 154702 189132 154708
rect 188252 153468 188304 153474
rect 188252 153410 188304 153416
rect 187792 152108 187844 152114
rect 187792 152050 187844 152056
rect 188264 151994 188292 153410
rect 189092 153270 189120 154702
rect 189080 153264 189132 153270
rect 189080 153206 189132 153212
rect 189078 152824 189134 152833
rect 189078 152759 189134 152768
rect 189092 151994 189120 152759
rect 189644 151994 189672 157422
rect 190564 155582 190592 159200
rect 191484 155650 191512 159200
rect 191564 156392 191616 156398
rect 191564 156334 191616 156340
rect 191472 155644 191524 155650
rect 191472 155586 191524 155592
rect 190552 155576 190604 155582
rect 190552 155518 190604 155524
rect 190458 155000 190514 155009
rect 190458 154935 190514 154944
rect 190472 151994 190500 154935
rect 190828 153604 190880 153610
rect 190828 153546 190880 153552
rect 190840 151994 190868 153546
rect 191576 151994 191604 156334
rect 191748 156188 191800 156194
rect 191748 156130 191800 156136
rect 191760 154630 191788 156130
rect 191748 154624 191800 154630
rect 191748 154566 191800 154572
rect 192496 154358 192524 159200
rect 193416 156398 193444 159200
rect 193404 156392 193456 156398
rect 193404 156334 193456 156340
rect 194048 156120 194100 156126
rect 194048 156062 194100 156068
rect 193128 155032 193180 155038
rect 193128 154974 193180 154980
rect 192484 154352 192536 154358
rect 192484 154294 192536 154300
rect 193140 153474 193168 154974
rect 193404 154420 193456 154426
rect 193404 154362 193456 154368
rect 193128 153468 193180 153474
rect 193128 153410 193180 153416
rect 192760 153332 192812 153338
rect 192760 153274 192812 153280
rect 192114 152960 192170 152969
rect 192114 152895 192170 152904
rect 192128 151994 192156 152895
rect 192772 151994 192800 153274
rect 193416 151994 193444 154362
rect 194060 151994 194088 156062
rect 194428 154766 194456 159200
rect 194784 158092 194836 158098
rect 194784 158034 194836 158040
rect 194416 154760 194468 154766
rect 194416 154702 194468 154708
rect 194796 151994 194824 158034
rect 195348 155582 195376 159200
rect 195428 157548 195480 157554
rect 195428 157490 195480 157496
rect 195336 155576 195388 155582
rect 195336 155518 195388 155524
rect 195440 151994 195468 157490
rect 195980 154896 196032 154902
rect 195980 154838 196032 154844
rect 195992 153542 196020 154838
rect 196360 154834 196388 159200
rect 197372 156330 197400 159200
rect 197360 156324 197412 156330
rect 197360 156266 197412 156272
rect 197452 156052 197504 156058
rect 197452 155994 197504 156000
rect 197360 154964 197412 154970
rect 197360 154906 197412 154912
rect 196348 154828 196400 154834
rect 196348 154770 196400 154776
rect 196532 154692 196584 154698
rect 196532 154634 196584 154640
rect 195980 153536 196032 153542
rect 195980 153478 196032 153484
rect 196072 153400 196124 153406
rect 196072 153342 196124 153348
rect 196084 151994 196112 153342
rect 183704 151988 184000 151994
rect 183652 151982 184000 151988
rect 183664 151966 184000 151982
rect 184308 151966 184644 151994
rect 184952 151966 185288 151994
rect 185688 151966 186024 151994
rect 186516 151966 186668 151994
rect 186976 151966 187312 151994
rect 187712 151966 187956 151994
rect 188264 151966 188600 151994
rect 189092 151966 189244 151994
rect 189644 151966 189888 151994
rect 190472 151966 190532 151994
rect 190840 151966 191176 151994
rect 191576 151966 191820 151994
rect 192128 151966 192464 151994
rect 192772 151966 193108 151994
rect 193416 151966 193752 151994
rect 194060 151966 194396 151994
rect 194796 151966 195132 151994
rect 195440 151966 195776 151994
rect 196084 151966 196420 151994
rect 196544 151910 196572 154634
rect 197372 153746 197400 154906
rect 197360 153740 197412 153746
rect 197360 153682 197412 153688
rect 197038 152108 197090 152114
rect 197038 152050 197090 152056
rect 197050 151980 197078 152050
rect 197464 151994 197492 155994
rect 198292 154766 198320 159200
rect 198280 154760 198332 154766
rect 198280 154702 198332 154708
rect 198740 154488 198792 154494
rect 198740 154430 198792 154436
rect 198004 153604 198056 153610
rect 198004 153546 198056 153552
rect 198016 151994 198044 153546
rect 198752 151994 198780 154430
rect 199304 154426 199332 159200
rect 199384 156120 199436 156126
rect 199384 156062 199436 156068
rect 199292 154420 199344 154426
rect 199292 154362 199344 154368
rect 199396 151994 199424 156062
rect 200224 155922 200252 159200
rect 200212 155916 200264 155922
rect 200212 155858 200264 155864
rect 200578 154728 200634 154737
rect 200578 154663 200634 154672
rect 200120 152040 200172 152046
rect 197464 151966 197708 151994
rect 198016 151966 198352 151994
rect 198752 151966 198996 151994
rect 199396 151966 199640 151994
rect 200592 151994 200620 154663
rect 201236 152114 201264 159200
rect 201866 156632 201922 156641
rect 201866 156567 201922 156576
rect 201500 154556 201552 154562
rect 201500 154498 201552 154504
rect 201224 152108 201276 152114
rect 201224 152050 201276 152056
rect 201512 151994 201540 154498
rect 201880 151994 201908 156567
rect 202248 154902 202276 159200
rect 202512 156664 202564 156670
rect 202512 156606 202564 156612
rect 202236 154896 202288 154902
rect 202236 154838 202288 154844
rect 202524 151994 202552 156606
rect 202788 155916 202840 155922
rect 202788 155858 202840 155864
rect 202800 154562 202828 155858
rect 202788 154556 202840 154562
rect 202788 154498 202840 154504
rect 203168 154494 203196 159200
rect 204180 155417 204208 159200
rect 204166 155408 204222 155417
rect 204166 155343 204222 155352
rect 203156 154488 203208 154494
rect 203156 154430 203208 154436
rect 203156 153468 203208 153474
rect 203156 153410 203208 153416
rect 203168 151994 203196 153410
rect 203892 153264 203944 153270
rect 203892 153206 203944 153212
rect 203904 151994 203932 153206
rect 205100 152046 205128 159200
rect 205824 157616 205876 157622
rect 205824 157558 205876 157564
rect 205640 156052 205692 156058
rect 205640 155994 205692 156000
rect 205652 154698 205680 155994
rect 205640 154692 205692 154698
rect 205640 154634 205692 154640
rect 205178 152552 205234 152561
rect 205178 152487 205234 152496
rect 205088 152040 205140 152046
rect 200172 151988 200284 151994
rect 200120 151982 200284 151988
rect 200132 151966 200284 151982
rect 200592 151966 200928 151994
rect 201512 151966 201572 151994
rect 201880 151966 202216 151994
rect 202524 151966 202860 151994
rect 203168 151966 203504 151994
rect 203904 151966 204240 151994
rect 205088 151982 205140 151988
rect 205192 151994 205220 152487
rect 205836 151994 205864 157558
rect 206112 155922 206140 159200
rect 206100 155916 206152 155922
rect 206100 155858 206152 155864
rect 207124 154970 207152 159200
rect 207202 157176 207258 157185
rect 207202 157111 207258 157120
rect 207112 154964 207164 154970
rect 207112 154906 207164 154912
rect 206468 153876 206520 153882
rect 206468 153818 206520 153824
rect 206480 151994 206508 153818
rect 207216 151994 207244 157111
rect 207756 156732 207808 156738
rect 207756 156674 207808 156680
rect 207768 151994 207796 156674
rect 208044 153882 208072 159200
rect 209056 156670 209084 159200
rect 209872 156800 209924 156806
rect 209872 156742 209924 156748
rect 209044 156664 209096 156670
rect 209044 156606 209096 156612
rect 209044 155372 209096 155378
rect 209044 155314 209096 155320
rect 208400 155236 208452 155242
rect 208400 155178 208452 155184
rect 208032 153876 208084 153882
rect 208032 153818 208084 153824
rect 208412 151994 208440 155178
rect 209056 151994 209084 155314
rect 209884 151994 209912 156742
rect 209976 155242 210004 159200
rect 210988 155378 211016 159200
rect 210976 155372 211028 155378
rect 210976 155314 211028 155320
rect 209964 155236 210016 155242
rect 209964 155178 210016 155184
rect 212000 154766 212028 159200
rect 212920 156738 212948 159200
rect 213000 156868 213052 156874
rect 213000 156810 213052 156816
rect 212908 156732 212960 156738
rect 212908 156674 212960 156680
rect 211068 154760 211120 154766
rect 211068 154702 211120 154708
rect 211988 154760 212040 154766
rect 211988 154702 212040 154708
rect 210332 152516 210384 152522
rect 210332 152458 210384 152464
rect 210344 151994 210372 152458
rect 205192 151966 205528 151994
rect 205836 151966 206172 151994
rect 206480 151966 206816 151994
rect 207216 151966 207460 151994
rect 207768 151966 208104 151994
rect 208412 151966 208748 151994
rect 209056 151966 209392 151994
rect 209884 151966 210036 151994
rect 210344 151966 210680 151994
rect 196532 151904 196584 151910
rect 196532 151846 196584 151852
rect 204548 151842 204884 151858
rect 211080 151842 211108 154702
rect 211160 153672 211212 153678
rect 211160 153614 211212 153620
rect 211172 151994 211200 153614
rect 211620 153536 211672 153542
rect 211620 153478 211672 153484
rect 211632 151994 211660 153478
rect 212540 152584 212592 152590
rect 212540 152526 212592 152532
rect 212552 151994 212580 152526
rect 213012 151994 213040 156810
rect 213932 155310 213960 159200
rect 214104 157684 214156 157690
rect 214104 157626 214156 157632
rect 213920 155304 213972 155310
rect 213920 155246 213972 155252
rect 211172 151966 211324 151994
rect 211632 151966 211968 151994
rect 212552 151966 212612 151994
rect 213012 151966 213256 151994
rect 214116 151858 214144 157626
rect 214288 154692 214340 154698
rect 214288 154634 214340 154640
rect 214300 151994 214328 154634
rect 214852 152522 214880 159200
rect 215864 155922 215892 159200
rect 215852 155916 215904 155922
rect 215852 155858 215904 155864
rect 216588 155916 216640 155922
rect 216588 155858 216640 155864
rect 216600 153814 216628 155858
rect 216876 154034 216904 159200
rect 217796 155553 217824 159200
rect 218808 156874 218836 159200
rect 218888 157752 218940 157758
rect 218888 157694 218940 157700
rect 218796 156868 218848 156874
rect 218796 156810 218848 156816
rect 218152 156800 218204 156806
rect 218152 156742 218204 156748
rect 217782 155544 217838 155553
rect 217782 155479 217838 155488
rect 216876 154006 216996 154034
rect 216864 153944 216916 153950
rect 216864 153886 216916 153892
rect 216220 153808 216272 153814
rect 216220 153750 216272 153756
rect 216588 153808 216640 153814
rect 216588 153750 216640 153756
rect 215576 152992 215628 152998
rect 215576 152934 215628 152940
rect 214932 152652 214984 152658
rect 214932 152594 214984 152600
rect 214840 152516 214892 152522
rect 214840 152458 214892 152464
rect 214944 151994 214972 152594
rect 215588 151994 215616 152934
rect 216232 151994 216260 153750
rect 216876 151994 216904 153886
rect 216968 152590 216996 154006
rect 217508 152720 217560 152726
rect 217508 152662 217560 152668
rect 216956 152584 217008 152590
rect 216956 152526 217008 152532
rect 217520 151994 217548 152662
rect 218164 151994 218192 156742
rect 218900 151994 218928 157694
rect 219728 155786 219756 159200
rect 220084 156936 220136 156942
rect 220084 156878 220136 156884
rect 219716 155780 219768 155786
rect 219716 155722 219768 155728
rect 219624 154012 219676 154018
rect 219624 153954 219676 153960
rect 219636 151994 219664 153954
rect 220096 151994 220124 156878
rect 220740 152658 220768 159200
rect 221370 157312 221426 157321
rect 221370 157247 221426 157256
rect 220820 152788 220872 152794
rect 220820 152730 220872 152736
rect 220728 152652 220780 152658
rect 220728 152594 220780 152600
rect 220832 151994 220860 152730
rect 221384 151994 221412 157247
rect 221752 156806 221780 159200
rect 221740 156800 221792 156806
rect 221740 156742 221792 156748
rect 222672 155922 222700 159200
rect 223580 156596 223632 156602
rect 223580 156538 223632 156544
rect 222660 155916 222712 155922
rect 222660 155858 222712 155864
rect 222108 155780 222160 155786
rect 222108 155722 222160 155728
rect 222120 153950 222148 155722
rect 222108 153944 222160 153950
rect 222108 153886 222160 153892
rect 222200 153740 222252 153746
rect 222200 153682 222252 153688
rect 222212 151994 222240 153682
rect 222752 152856 222804 152862
rect 222752 152798 222804 152804
rect 222764 151994 222792 152798
rect 223592 151994 223620 156538
rect 223684 154698 223712 159200
rect 223672 154692 223724 154698
rect 223672 154634 223724 154640
rect 224040 152924 224092 152930
rect 224040 152866 224092 152872
rect 224052 151994 224080 152866
rect 224604 152726 224632 159200
rect 225328 157004 225380 157010
rect 225328 156946 225380 156952
rect 225052 155780 225104 155786
rect 225052 155722 225104 155728
rect 224960 154080 225012 154086
rect 224960 154022 225012 154028
rect 224592 152720 224644 152726
rect 224592 152662 224644 152668
rect 224972 151994 225000 154022
rect 225064 153270 225092 155722
rect 225052 153264 225104 153270
rect 225052 153206 225104 153212
rect 225340 151994 225368 156946
rect 225616 155786 225644 159200
rect 225972 156460 226024 156466
rect 225972 156402 226024 156408
rect 225604 155780 225656 155786
rect 225604 155722 225656 155728
rect 225984 151994 226012 156402
rect 226628 155446 226656 159200
rect 226524 155440 226576 155446
rect 226524 155382 226576 155388
rect 226616 155440 226668 155446
rect 226616 155382 226668 155388
rect 226536 151994 226564 155382
rect 227258 155272 227314 155281
rect 227258 155207 227314 155216
rect 227272 151994 227300 155207
rect 227548 154018 227576 159200
rect 228560 156942 228588 159200
rect 228548 156936 228600 156942
rect 228548 156878 228600 156884
rect 229480 155854 229508 159200
rect 229468 155848 229520 155854
rect 229468 155790 229520 155796
rect 230492 155514 230520 159200
rect 230572 157072 230624 157078
rect 230572 157014 230624 157020
rect 229284 155508 229336 155514
rect 229284 155450 229336 155456
rect 230480 155508 230532 155514
rect 230480 155450 230532 155456
rect 229192 155168 229244 155174
rect 229192 155110 229244 155116
rect 227536 154012 227588 154018
rect 227536 153954 227588 153960
rect 229204 153542 229232 155110
rect 229192 153536 229244 153542
rect 229192 153478 229244 153484
rect 227904 153060 227956 153066
rect 227904 153002 227956 153008
rect 227916 151994 227944 153002
rect 228548 152448 228600 152454
rect 228548 152390 228600 152396
rect 228560 151994 228588 152390
rect 229296 151994 229324 155450
rect 229836 153264 229888 153270
rect 229836 153206 229888 153212
rect 229848 151994 229876 153206
rect 230584 151994 230612 157014
rect 231124 156528 231176 156534
rect 231124 156470 231176 156476
rect 231136 151994 231164 156470
rect 231504 155689 231532 159200
rect 231490 155680 231546 155689
rect 231490 155615 231546 155624
rect 231860 153128 231912 153134
rect 231860 153070 231912 153076
rect 231872 151994 231900 153070
rect 232424 152794 232452 159200
rect 233436 155718 233464 159200
rect 233424 155712 233476 155718
rect 233424 155654 233476 155660
rect 233148 155508 233200 155514
rect 233148 155450 233200 155456
rect 232504 154148 232556 154154
rect 232504 154090 232556 154096
rect 232412 152788 232464 152794
rect 232412 152730 232464 152736
rect 232516 151994 232544 154090
rect 233160 154086 233188 155450
rect 233240 155440 233292 155446
rect 233240 155382 233292 155388
rect 233148 154080 233200 154086
rect 233148 154022 233200 154028
rect 233252 153746 233280 155382
rect 234356 155281 234384 159200
rect 234620 155440 234672 155446
rect 234620 155382 234672 155388
rect 234342 155272 234398 155281
rect 234342 155207 234398 155216
rect 233240 153740 233292 153746
rect 233240 153682 233292 153688
rect 233240 153196 233292 153202
rect 233240 153138 233292 153144
rect 233252 151994 233280 153138
rect 233792 152380 233844 152386
rect 233792 152322 233844 152328
rect 233804 151994 233832 152322
rect 234632 151994 234660 155382
rect 235368 154154 235396 159200
rect 236000 157140 236052 157146
rect 236000 157082 236052 157088
rect 235356 154148 235408 154154
rect 235356 154090 235408 154096
rect 235080 153536 235132 153542
rect 235080 153478 235132 153484
rect 235092 151994 235120 153478
rect 236012 151994 236040 157082
rect 236288 157010 236316 159200
rect 237012 157276 237064 157282
rect 237012 157218 237064 157224
rect 236276 157004 236328 157010
rect 236276 156946 236328 156952
rect 236368 156256 236420 156262
rect 236368 156198 236420 156204
rect 236380 151994 236408 156198
rect 237024 151994 237052 157218
rect 237300 155038 237328 159200
rect 238312 155446 238340 159200
rect 238392 157208 238444 157214
rect 238392 157150 238444 157156
rect 238300 155440 238352 155446
rect 238300 155382 238352 155388
rect 237196 155032 237248 155038
rect 237196 154974 237248 154980
rect 237288 155032 237340 155038
rect 237288 154974 237340 154980
rect 237208 154850 237236 154974
rect 237208 154822 237420 154850
rect 237392 153678 237420 154822
rect 237656 154216 237708 154222
rect 237656 154158 237708 154164
rect 237380 153672 237432 153678
rect 237380 153614 237432 153620
rect 237668 151994 237696 154158
rect 238404 151994 238432 157150
rect 239232 155650 239260 159200
rect 239220 155644 239272 155650
rect 239220 155586 239272 155592
rect 239588 155168 239640 155174
rect 239588 155110 239640 155116
rect 239600 151994 239628 155110
rect 240244 154442 240272 159200
rect 241164 155854 241192 159200
rect 241612 156188 241664 156194
rect 241612 156130 241664 156136
rect 241152 155848 241204 155854
rect 241152 155790 241204 155796
rect 241428 155644 241480 155650
rect 241428 155586 241480 155592
rect 240244 154414 240364 154442
rect 240232 154284 240284 154290
rect 240232 154226 240284 154232
rect 240244 151994 240272 154226
rect 240336 152862 240364 154414
rect 241440 154222 241468 155586
rect 241428 154216 241480 154222
rect 241428 154158 241480 154164
rect 240324 152856 240376 152862
rect 240324 152798 240376 152804
rect 240968 152312 241020 152318
rect 240968 152254 241020 152260
rect 240980 151994 241008 152254
rect 241624 151994 241652 156130
rect 242176 155582 242204 159200
rect 243188 155718 243216 159200
rect 244108 157078 244136 159200
rect 244096 157072 244148 157078
rect 244096 157014 244148 157020
rect 244372 156120 244424 156126
rect 244372 156062 244424 156068
rect 243176 155712 243228 155718
rect 243176 155654 243228 155660
rect 242164 155576 242216 155582
rect 242164 155518 242216 155524
rect 242992 155100 243044 155106
rect 242992 155042 243044 155048
rect 242256 154624 242308 154630
rect 242256 154566 242308 154572
rect 242268 151994 242296 154566
rect 242900 153672 242952 153678
rect 242900 153614 242952 153620
rect 242912 151994 242940 153614
rect 243004 153474 243032 155042
rect 242992 153468 243044 153474
rect 242992 153410 243044 153416
rect 243866 152244 243918 152250
rect 243866 152186 243918 152192
rect 214300 151966 214636 151994
rect 214944 151966 215280 151994
rect 215588 151966 215924 151994
rect 216232 151966 216568 151994
rect 216876 151966 217212 151994
rect 217520 151966 217856 151994
rect 218164 151966 218500 151994
rect 218900 151966 219144 151994
rect 219636 151966 219788 151994
rect 220096 151966 220432 151994
rect 220832 151966 221076 151994
rect 221384 151966 221720 151994
rect 222212 151966 222364 151994
rect 222764 151966 223100 151994
rect 223592 151966 223744 151994
rect 224052 151966 224388 151994
rect 224972 151966 225032 151994
rect 225340 151966 225676 151994
rect 225984 151966 226320 151994
rect 226536 151966 226964 151994
rect 227272 151966 227608 151994
rect 227916 151966 228252 151994
rect 228560 151966 228896 151994
rect 229296 151966 229540 151994
rect 229848 151966 230184 151994
rect 230584 151966 230828 151994
rect 231136 151966 231472 151994
rect 231872 151966 232208 151994
rect 232516 151966 232852 151994
rect 233252 151966 233496 151994
rect 233804 151966 234140 151994
rect 234632 151966 234784 151994
rect 235092 151966 235428 151994
rect 236012 151966 236072 151994
rect 236380 151966 236716 151994
rect 237024 151966 237360 151994
rect 237668 151966 238004 151994
rect 238404 151966 238648 151994
rect 238956 151978 239292 151994
rect 238944 151972 239292 151978
rect 238996 151966 239292 151972
rect 239600 151966 239936 151994
rect 240244 151966 240580 151994
rect 240980 151966 241316 151994
rect 241624 151966 241960 151994
rect 242268 151966 242604 151994
rect 242912 151966 243248 151994
rect 243878 151980 243906 152186
rect 244384 151994 244412 156062
rect 245120 155650 245148 159200
rect 245108 155644 245160 155650
rect 245108 155586 245160 155592
rect 245568 154828 245620 154834
rect 245568 154770 245620 154776
rect 245580 153338 245608 154770
rect 246040 154630 246068 159200
rect 246120 157344 246172 157350
rect 246120 157286 246172 157292
rect 246028 154624 246080 154630
rect 246028 154566 246080 154572
rect 245660 153468 245712 153474
rect 245660 153410 245712 153416
rect 245568 153332 245620 153338
rect 245568 153274 245620 153280
rect 245154 152176 245206 152182
rect 245154 152118 245206 152124
rect 244384 151966 244536 151994
rect 245166 151980 245194 152118
rect 245672 151994 245700 153410
rect 246132 151994 246160 157286
rect 247052 154290 247080 159200
rect 248064 157334 248092 159200
rect 248064 157306 248184 157334
rect 247408 154352 247460 154358
rect 247408 154294 247460 154300
rect 247040 154284 247092 154290
rect 247040 154226 247092 154232
rect 247420 151994 247448 154294
rect 248052 153672 248104 153678
rect 248052 153614 248104 153620
rect 248064 151994 248092 153614
rect 248156 152930 248184 157306
rect 248696 156392 248748 156398
rect 248696 156334 248748 156340
rect 248144 152924 248196 152930
rect 248144 152866 248196 152872
rect 248708 151994 248736 156334
rect 248984 154834 249012 159200
rect 249340 155984 249392 155990
rect 249340 155926 249392 155932
rect 248972 154828 249024 154834
rect 248972 154770 249024 154776
rect 249352 151994 249380 155926
rect 249996 155582 250024 159200
rect 250916 155650 250944 159200
rect 251928 157146 251956 159200
rect 252940 159174 253060 159200
rect 251916 157140 251968 157146
rect 251916 157082 251968 157088
rect 251364 156324 251416 156330
rect 251364 156266 251416 156272
rect 250904 155644 250956 155650
rect 250904 155586 250956 155592
rect 249984 155576 250036 155582
rect 249984 155518 250036 155524
rect 251178 155408 251234 155417
rect 251178 155343 251234 155352
rect 249800 154556 249852 154562
rect 249800 154498 249852 154504
rect 249812 153270 249840 154498
rect 249984 154352 250036 154358
rect 249984 154294 250036 154300
rect 249800 153264 249852 153270
rect 249800 153206 249852 153212
rect 249996 151994 250024 154294
rect 251192 153542 251220 155343
rect 251180 153536 251232 153542
rect 251180 153478 251232 153484
rect 250720 153332 250772 153338
rect 250720 153274 250772 153280
rect 250732 151994 250760 153274
rect 251376 151994 251404 156266
rect 253216 155378 253244 159310
rect 253846 159200 253902 160000
rect 254858 159200 254914 160000
rect 255778 159200 255834 160000
rect 256790 159200 256846 160000
rect 257802 159200 257858 160000
rect 258722 159200 258778 160000
rect 259734 159200 259790 160000
rect 260654 159200 260710 160000
rect 261666 159200 261722 160000
rect 262678 159200 262734 160000
rect 263598 159200 263654 160000
rect 264610 159200 264666 160000
rect 265530 159200 265586 160000
rect 266542 159200 266598 160000
rect 267554 159200 267610 160000
rect 268474 159200 268530 160000
rect 269486 159200 269542 160000
rect 270406 159200 270462 160000
rect 271418 159200 271474 160000
rect 272338 159200 272394 160000
rect 273350 159200 273406 160000
rect 274362 159200 274418 160000
rect 275282 159200 275338 160000
rect 276294 159200 276350 160000
rect 277214 159200 277270 160000
rect 278226 159200 278282 160000
rect 279238 159200 279294 160000
rect 280158 159200 280214 160000
rect 281170 159200 281226 160000
rect 282090 159200 282146 160000
rect 283102 159200 283158 160000
rect 284114 159200 284170 160000
rect 285034 159200 285090 160000
rect 286046 159200 286102 160000
rect 286966 159200 287022 160000
rect 287978 159200 288034 160000
rect 288990 159200 289046 160000
rect 289910 159200 289966 160000
rect 290922 159200 290978 160000
rect 291842 159200 291898 160000
rect 292854 159200 292910 160000
rect 293866 159200 293922 160000
rect 294786 159200 294842 160000
rect 295798 159200 295854 160000
rect 296718 159200 296774 160000
rect 297730 159200 297786 160000
rect 298742 159200 298798 160000
rect 299662 159200 299718 160000
rect 300674 159200 300730 160000
rect 301594 159200 301650 160000
rect 302606 159200 302662 160000
rect 303618 159200 303674 160000
rect 304538 159200 304594 160000
rect 305550 159200 305606 160000
rect 306470 159200 306526 160000
rect 307482 159200 307538 160000
rect 308494 159200 308550 160000
rect 309414 159200 309470 160000
rect 310426 159200 310482 160000
rect 311346 159200 311402 160000
rect 312358 159200 312414 160000
rect 313278 159200 313334 160000
rect 314290 159200 314346 160000
rect 315302 159200 315358 160000
rect 316222 159200 316278 160000
rect 317234 159200 317290 160000
rect 318154 159200 318210 160000
rect 319166 159200 319222 160000
rect 320178 159200 320234 160000
rect 321098 159200 321154 160000
rect 322110 159200 322166 160000
rect 323030 159200 323086 160000
rect 324042 159200 324098 160000
rect 325054 159200 325110 160000
rect 325974 159200 326030 160000
rect 326986 159200 327042 160000
rect 327906 159200 327962 160000
rect 328918 159200 328974 160000
rect 329930 159200 329986 160000
rect 330850 159200 330906 160000
rect 331862 159200 331918 160000
rect 332782 159200 332838 160000
rect 333794 159200 333850 160000
rect 334806 159200 334862 160000
rect 335726 159200 335782 160000
rect 336738 159200 336794 160000
rect 337658 159200 337714 160000
rect 338670 159200 338726 160000
rect 339682 159200 339738 160000
rect 340602 159200 340658 160000
rect 341614 159200 341670 160000
rect 342534 159200 342590 160000
rect 343546 159200 343602 160000
rect 344558 159200 344614 160000
rect 345478 159200 345534 160000
rect 346490 159200 346546 160000
rect 347410 159202 347466 160000
rect 347516 159310 347728 159338
rect 347516 159202 347544 159310
rect 347410 159200 347544 159202
rect 253204 155372 253256 155378
rect 253204 155314 253256 155320
rect 253860 154426 253888 159200
rect 252652 154420 252704 154426
rect 252652 154362 252704 154368
rect 253848 154420 253900 154426
rect 253848 154362 253900 154368
rect 252664 151994 252692 154362
rect 254872 154358 254900 159200
rect 255320 154760 255372 154766
rect 255320 154702 255372 154708
rect 255332 154494 255360 154702
rect 255320 154488 255372 154494
rect 255320 154430 255372 154436
rect 254860 154352 254912 154358
rect 254860 154294 254912 154300
rect 255320 153672 255372 153678
rect 255320 153614 255372 153620
rect 253296 153604 253348 153610
rect 253296 153546 253348 153552
rect 253308 151994 253336 153546
rect 254584 153264 254636 153270
rect 254584 153206 254636 153212
rect 254262 152108 254314 152114
rect 254262 152050 254314 152056
rect 245672 151966 245824 151994
rect 246132 151966 246468 151994
rect 247420 151966 247756 151994
rect 248064 151966 248400 151994
rect 248708 151966 249044 151994
rect 249352 151966 249688 151994
rect 249996 151966 250332 151994
rect 250732 151966 251068 151994
rect 251376 151966 251712 151994
rect 252664 151966 253000 151994
rect 253308 151966 253644 151994
rect 254274 151980 254302 152050
rect 254596 151994 254624 153206
rect 255332 151994 255360 153614
rect 255792 152998 255820 159200
rect 256700 154964 256752 154970
rect 256700 154906 256752 154912
rect 255872 153604 255924 153610
rect 255872 153546 255924 153552
rect 255780 152992 255832 152998
rect 255780 152934 255832 152940
rect 255884 151994 255912 153546
rect 256712 153270 256740 154906
rect 256804 154766 256832 159200
rect 257160 156052 257212 156058
rect 257160 155994 257212 156000
rect 256792 154760 256844 154766
rect 256792 154702 256844 154708
rect 256700 153264 256752 153270
rect 256700 153206 256752 153212
rect 256700 152040 256752 152046
rect 254596 151966 254932 151994
rect 255332 151966 255576 151994
rect 255884 151966 256220 151994
rect 257172 151994 257200 155994
rect 257816 154970 257844 159200
rect 258736 155922 258764 159200
rect 259092 156664 259144 156670
rect 259092 156606 259144 156612
rect 258724 155916 258776 155922
rect 258724 155858 258776 155864
rect 257804 154964 257856 154970
rect 257804 154906 257856 154912
rect 258448 153876 258500 153882
rect 258448 153818 258500 153824
rect 258080 153264 258132 153270
rect 258080 153206 258132 153212
rect 258092 151994 258120 153206
rect 258460 151994 258488 153818
rect 259104 151994 259132 156606
rect 259368 154896 259420 154902
rect 259368 154838 259420 154844
rect 259380 153406 259408 154838
rect 259368 153400 259420 153406
rect 259368 153342 259420 153348
rect 259748 153066 259776 159200
rect 260668 155242 260696 159200
rect 261680 155417 261708 159200
rect 261760 156732 261812 156738
rect 261760 156674 261812 156680
rect 261666 155408 261722 155417
rect 261666 155343 261722 155352
rect 259828 155236 259880 155242
rect 259828 155178 259880 155184
rect 260656 155236 260708 155242
rect 260656 155178 260708 155184
rect 259736 153060 259788 153066
rect 259736 153002 259788 153008
rect 259840 151994 259868 155178
rect 261116 154488 261168 154494
rect 261116 154430 261168 154436
rect 260472 153400 260524 153406
rect 260472 153342 260524 153348
rect 260484 151994 260512 153342
rect 261128 151994 261156 154430
rect 261772 151994 261800 156674
rect 262128 155916 262180 155922
rect 262128 155858 262180 155864
rect 262140 153882 262168 155858
rect 262692 155666 262720 159200
rect 262692 155650 262812 155666
rect 262692 155644 262824 155650
rect 262692 155638 262772 155644
rect 262772 155586 262824 155592
rect 262218 155544 262274 155553
rect 262218 155479 262274 155488
rect 262128 153876 262180 153882
rect 262128 153818 262180 153824
rect 262232 153678 262260 155479
rect 262404 155304 262456 155310
rect 262404 155246 262456 155252
rect 262220 153672 262272 153678
rect 262220 153614 262272 153620
rect 262416 151994 262444 155246
rect 263612 155242 263640 159200
rect 264624 155786 264652 159200
rect 263784 155780 263836 155786
rect 263784 155722 263836 155728
rect 264612 155780 264664 155786
rect 264612 155722 264664 155728
rect 263600 155236 263652 155242
rect 263600 155178 263652 155184
rect 263692 153808 263744 153814
rect 263692 153750 263744 153756
rect 263048 152516 263100 152522
rect 263048 152458 263100 152464
rect 263060 151994 263088 152458
rect 263704 151994 263732 153750
rect 263796 153338 263824 155722
rect 265544 155514 265572 159200
rect 265624 156868 265676 156874
rect 265624 156810 265676 156816
rect 265072 155508 265124 155514
rect 265072 155450 265124 155456
rect 265532 155508 265584 155514
rect 265532 155450 265584 155456
rect 264980 153672 265032 153678
rect 264980 153614 265032 153620
rect 263784 153332 263836 153338
rect 263784 153274 263836 153280
rect 264336 152584 264388 152590
rect 264336 152526 264388 152532
rect 264348 151994 264376 152526
rect 264992 151994 265020 153614
rect 265084 153610 265112 155450
rect 265072 153604 265124 153610
rect 265072 153546 265124 153552
rect 265636 151994 265664 156810
rect 266556 155514 266584 159200
rect 267568 155553 267596 159200
rect 267832 156800 267884 156806
rect 267832 156742 267884 156748
rect 267554 155544 267610 155553
rect 266452 155508 266504 155514
rect 266452 155450 266504 155456
rect 266544 155508 266596 155514
rect 267554 155479 267610 155488
rect 266544 155450 266596 155456
rect 266360 155032 266412 155038
rect 266360 154974 266412 154980
rect 266372 154494 266400 154974
rect 266360 154488 266412 154494
rect 266360 154430 266412 154436
rect 266464 153950 266492 155450
rect 266360 153944 266412 153950
rect 266360 153886 266412 153892
rect 266452 153944 266504 153950
rect 266452 153886 266504 153892
rect 266372 151994 266400 153886
rect 266912 152652 266964 152658
rect 266912 152594 266964 152600
rect 266924 151994 266952 152594
rect 267844 151994 267872 156742
rect 268488 155786 268516 159200
rect 268476 155780 268528 155786
rect 268476 155722 268528 155728
rect 269396 155168 269448 155174
rect 269396 155110 269448 155116
rect 269408 154970 269436 155110
rect 269500 155038 269528 159200
rect 270420 155310 270448 159200
rect 270316 155304 270368 155310
rect 270316 155246 270368 155252
rect 270408 155304 270460 155310
rect 270408 155246 270460 155252
rect 269488 155032 269540 155038
rect 269488 154974 269540 154980
rect 269396 154964 269448 154970
rect 269396 154906 269448 154912
rect 269028 154692 269080 154698
rect 269028 154634 269080 154640
rect 268200 153332 268252 153338
rect 268200 153274 268252 153280
rect 268212 151994 268240 153274
rect 269040 153218 269068 154634
rect 270328 153542 270356 155246
rect 270868 153740 270920 153746
rect 270868 153682 270920 153688
rect 270500 153604 270552 153610
rect 270500 153546 270552 153552
rect 270316 153536 270368 153542
rect 270316 153478 270368 153484
rect 269040 153190 269160 153218
rect 269132 151994 269160 153190
rect 269580 152720 269632 152726
rect 269580 152662 269632 152668
rect 269592 151994 269620 152662
rect 270512 151994 270540 153546
rect 270880 151994 270908 153682
rect 271432 152522 271460 159200
rect 272156 156936 272208 156942
rect 272156 156878 272208 156884
rect 271970 155680 272026 155689
rect 271970 155615 272026 155624
rect 271696 154964 271748 154970
rect 271696 154906 271748 154912
rect 271512 154012 271564 154018
rect 271512 153954 271564 153960
rect 271420 152516 271472 152522
rect 271420 152458 271472 152464
rect 271524 151994 271552 153954
rect 271708 153338 271736 154906
rect 271788 154624 271840 154630
rect 271788 154566 271840 154572
rect 271800 153814 271828 154566
rect 271788 153808 271840 153814
rect 271788 153750 271840 153756
rect 271984 153746 272012 155615
rect 271972 153740 272024 153746
rect 271972 153682 272024 153688
rect 271696 153332 271748 153338
rect 271696 153274 271748 153280
rect 272168 151994 272196 156878
rect 272352 154970 272380 159200
rect 273364 155106 273392 159200
rect 274376 155514 274404 159200
rect 274364 155508 274416 155514
rect 274364 155450 274416 155456
rect 275296 155174 275324 159200
rect 275926 155272 275982 155281
rect 275926 155207 275982 155216
rect 274640 155168 274692 155174
rect 274640 155110 274692 155116
rect 275284 155168 275336 155174
rect 275284 155110 275336 155116
rect 273352 155100 273404 155106
rect 273352 155042 273404 155048
rect 272340 154964 272392 154970
rect 272340 154906 272392 154912
rect 273444 154080 273496 154086
rect 273444 154022 273496 154028
rect 272800 153536 272852 153542
rect 272800 153478 272852 153484
rect 272812 151994 272840 153478
rect 273456 151994 273484 154022
rect 274652 154018 274680 155110
rect 275376 154488 275428 154494
rect 275376 154430 275428 154436
rect 274640 154012 274692 154018
rect 274640 153954 274692 153960
rect 274088 153740 274140 153746
rect 274088 153682 274140 153688
rect 274100 151994 274128 153682
rect 274732 152788 274784 152794
rect 274732 152730 274784 152736
rect 274744 151994 274772 152730
rect 275388 151994 275416 154430
rect 275940 153218 275968 155207
rect 276308 154834 276336 159200
rect 277228 154970 277256 159200
rect 277492 157004 277544 157010
rect 277492 156946 277544 156952
rect 277308 155372 277360 155378
rect 277308 155314 277360 155320
rect 277320 155145 277348 155314
rect 277306 155136 277362 155145
rect 277306 155071 277362 155080
rect 277398 155000 277454 155009
rect 276756 154964 276808 154970
rect 276756 154906 276808 154912
rect 277216 154964 277268 154970
rect 277398 154935 277454 154944
rect 277216 154906 277268 154912
rect 276020 154828 276072 154834
rect 276020 154770 276072 154776
rect 276296 154828 276348 154834
rect 276296 154770 276348 154776
rect 276032 154154 276060 154770
rect 276020 154148 276072 154154
rect 276020 154090 276072 154096
rect 276768 154086 276796 154906
rect 276664 154080 276716 154086
rect 276664 154022 276716 154028
rect 276756 154080 276808 154086
rect 276756 154022 276808 154028
rect 275940 153190 276060 153218
rect 276032 151994 276060 153190
rect 276676 151994 276704 154022
rect 277412 153474 277440 154935
rect 277400 153468 277452 153474
rect 277400 153410 277452 153416
rect 277504 151994 277532 156946
rect 278240 155786 278268 159200
rect 278228 155780 278280 155786
rect 278228 155722 278280 155728
rect 279252 155446 279280 159200
rect 280172 155582 280200 159200
rect 280252 155916 280304 155922
rect 280252 155858 280304 155864
rect 280160 155576 280212 155582
rect 280160 155518 280212 155524
rect 279148 155440 279200 155446
rect 279148 155382 279200 155388
rect 279240 155440 279292 155446
rect 279240 155382 279292 155388
rect 279160 153746 279188 155382
rect 279332 154216 279384 154222
rect 279332 154158 279384 154164
rect 279148 153740 279200 153746
rect 279148 153682 279200 153688
rect 278780 153468 278832 153474
rect 278780 153410 278832 153416
rect 277952 153332 278004 153338
rect 277952 153274 278004 153280
rect 277964 151994 277992 153274
rect 278792 151994 278820 153410
rect 279344 151994 279372 154158
rect 280264 153610 280292 155858
rect 281184 154766 281212 159200
rect 281448 155848 281500 155854
rect 281448 155790 281500 155796
rect 281172 154760 281224 154766
rect 281172 154702 281224 154708
rect 280620 153672 280672 153678
rect 280620 153614 280672 153620
rect 280252 153604 280304 153610
rect 280252 153546 280304 153552
rect 280160 152856 280212 152862
rect 280160 152798 280212 152804
rect 280172 151994 280200 152798
rect 280632 151994 280660 153614
rect 281460 153218 281488 155790
rect 282104 155106 282132 159200
rect 282552 157072 282604 157078
rect 282552 157014 282604 157020
rect 282092 155100 282144 155106
rect 282092 155042 282144 155048
rect 281540 154556 281592 154562
rect 281540 154498 281592 154504
rect 281552 153678 281580 154498
rect 281540 153672 281592 153678
rect 281540 153614 281592 153620
rect 281908 153604 281960 153610
rect 281908 153546 281960 153552
rect 281460 153190 281580 153218
rect 281552 151994 281580 153190
rect 281920 151994 281948 153546
rect 282564 151994 282592 157014
rect 283116 155718 283144 159200
rect 284128 155922 284156 159200
rect 284116 155916 284168 155922
rect 284116 155858 284168 155864
rect 284392 155848 284444 155854
rect 284392 155790 284444 155796
rect 282920 155712 282972 155718
rect 282920 155654 282972 155660
rect 283104 155712 283156 155718
rect 283104 155654 283156 155660
rect 282932 154562 282960 155654
rect 283288 154692 283340 154698
rect 283288 154634 283340 154640
rect 282920 154556 282972 154562
rect 282920 154498 282972 154504
rect 283300 153814 283328 154634
rect 284024 154488 284076 154494
rect 284024 154430 284076 154436
rect 283196 153808 283248 153814
rect 283196 153750 283248 153756
rect 283288 153808 283340 153814
rect 283288 153750 283340 153756
rect 283208 151994 283236 153750
rect 284036 151994 284064 154430
rect 284404 153610 284432 155790
rect 285048 154698 285076 159200
rect 286060 154902 286088 159200
rect 286980 155854 287008 159200
rect 287796 157140 287848 157146
rect 287796 157082 287848 157088
rect 286968 155848 287020 155854
rect 286968 155790 287020 155796
rect 285680 154896 285732 154902
rect 285680 154838 285732 154844
rect 286048 154896 286100 154902
rect 286048 154838 286100 154844
rect 285036 154692 285088 154698
rect 285036 154634 285088 154640
rect 285692 154494 285720 154838
rect 285680 154488 285732 154494
rect 285680 154430 285732 154436
rect 284484 154284 284536 154290
rect 284484 154226 284536 154232
rect 284392 153604 284444 153610
rect 284392 153546 284444 153552
rect 284496 151994 284524 154226
rect 285680 154216 285732 154222
rect 285680 154158 285732 154164
rect 285692 153270 285720 154158
rect 285772 154148 285824 154154
rect 285772 154090 285824 154096
rect 285680 153264 285732 153270
rect 285680 153206 285732 153212
rect 285128 152924 285180 152930
rect 285128 152866 285180 152872
rect 285140 151994 285168 152866
rect 285784 151994 285812 154090
rect 286416 153604 286468 153610
rect 286416 153546 286468 153552
rect 286428 151994 286456 153546
rect 287244 153264 287296 153270
rect 287244 153206 287296 153212
rect 287256 151994 287284 153206
rect 287808 151994 287836 157082
rect 287992 155242 288020 159200
rect 287980 155236 288032 155242
rect 287980 155178 288032 155184
rect 289004 154630 289032 159200
rect 289268 154828 289320 154834
rect 289268 154770 289320 154776
rect 288348 154624 288400 154630
rect 288348 154566 288400 154572
rect 288992 154624 289044 154630
rect 288992 154566 289044 154572
rect 288360 153610 288388 154566
rect 289084 154420 289136 154426
rect 289084 154362 289136 154368
rect 288440 154012 288492 154018
rect 288440 153954 288492 153960
rect 288348 153604 288400 153610
rect 288348 153546 288400 153552
rect 288452 151994 288480 153954
rect 289096 151994 289124 154362
rect 289280 154290 289308 154770
rect 289820 154352 289872 154358
rect 289820 154294 289872 154300
rect 289268 154284 289320 154290
rect 289268 154226 289320 154232
rect 289832 151994 289860 154294
rect 289924 154018 289952 159200
rect 290936 155582 290964 159200
rect 291752 155916 291804 155922
rect 291752 155858 291804 155864
rect 290832 155576 290884 155582
rect 290832 155518 290884 155524
rect 290924 155576 290976 155582
rect 290924 155518 290976 155524
rect 290844 154222 290872 155518
rect 290832 154216 290884 154222
rect 290832 154158 290884 154164
rect 291764 154154 291792 155858
rect 291752 154148 291804 154154
rect 291752 154090 291804 154096
rect 291856 154086 291884 159200
rect 292868 155922 292896 159200
rect 292856 155916 292908 155922
rect 292856 155858 292908 155864
rect 292762 155408 292818 155417
rect 292762 155343 292818 155352
rect 292580 155032 292632 155038
rect 292580 154974 292632 154980
rect 292592 154358 292620 154974
rect 292580 154352 292632 154358
rect 292580 154294 292632 154300
rect 291200 154080 291252 154086
rect 291200 154022 291252 154028
rect 291844 154080 291896 154086
rect 291844 154022 291896 154028
rect 289912 154012 289964 154018
rect 289912 153954 289964 153960
rect 290372 152992 290424 152998
rect 290372 152934 290424 152940
rect 290384 151994 290412 152934
rect 291212 151994 291240 154022
rect 292580 153876 292632 153882
rect 292580 153818 292632 153824
rect 291660 153672 291712 153678
rect 291660 153614 291712 153620
rect 291672 151994 291700 153614
rect 292592 151994 292620 153818
rect 292776 153678 292804 155343
rect 293880 154834 293908 159200
rect 294800 155038 294828 159200
rect 295812 155650 295840 159200
rect 295524 155644 295576 155650
rect 295524 155586 295576 155592
rect 295800 155644 295852 155650
rect 295800 155586 295852 155592
rect 294696 155032 294748 155038
rect 294696 154974 294748 154980
rect 294788 155032 294840 155038
rect 294788 154974 294840 154980
rect 293868 154828 293920 154834
rect 293868 154770 293920 154776
rect 293592 153740 293644 153746
rect 293592 153682 293644 153688
rect 292764 153672 292816 153678
rect 292764 153614 292816 153620
rect 292948 153060 293000 153066
rect 292948 153002 293000 153008
rect 292960 151994 292988 153002
rect 293604 151994 293632 153682
rect 294236 153672 294288 153678
rect 294236 153614 294288 153620
rect 294248 151994 294276 153614
rect 294708 152130 294736 154974
rect 295340 154760 295392 154766
rect 295340 154702 295392 154708
rect 295352 153882 295380 154702
rect 295340 153876 295392 153882
rect 295340 153818 295392 153824
rect 294708 152102 294828 152130
rect 294800 151994 294828 152102
rect 295536 151994 295564 155586
rect 296732 155530 296760 159200
rect 296732 155514 296944 155530
rect 296732 155508 296956 155514
rect 296732 155502 296904 155508
rect 296904 155450 296956 155456
rect 296720 155440 296772 155446
rect 296720 155382 296772 155388
rect 296732 155242 296760 155382
rect 296720 155236 296772 155242
rect 296720 155178 296772 155184
rect 297744 154766 297772 159200
rect 298190 155544 298246 155553
rect 298190 155479 298246 155488
rect 298008 155168 298060 155174
rect 298008 155110 298060 155116
rect 297916 154964 297968 154970
rect 297916 154906 297968 154912
rect 297732 154760 297784 154766
rect 297732 154702 297784 154708
rect 296996 153944 297048 153950
rect 296996 153886 297048 153892
rect 296168 153808 296220 153814
rect 296168 153750 296220 153756
rect 296180 151994 296208 153750
rect 297008 151994 297036 153886
rect 297548 153604 297600 153610
rect 297548 153546 297600 153552
rect 297560 151994 297588 153546
rect 297928 153406 297956 154906
rect 298020 153542 298048 155110
rect 298008 153536 298060 153542
rect 298008 153478 298060 153484
rect 297916 153400 297968 153406
rect 297916 153342 297968 153348
rect 298204 151994 298232 155479
rect 298756 155242 298784 159200
rect 298744 155236 298796 155242
rect 298744 155178 298796 155184
rect 299676 154970 299704 159200
rect 300124 155304 300176 155310
rect 300124 155246 300176 155252
rect 299664 154964 299716 154970
rect 299664 154906 299716 154912
rect 298836 154556 298888 154562
rect 298836 154498 298888 154504
rect 298848 151994 298876 154498
rect 299480 154352 299532 154358
rect 299480 154294 299532 154300
rect 299492 151994 299520 154294
rect 300136 151994 300164 155246
rect 300688 155106 300716 159200
rect 301608 155174 301636 159200
rect 302620 155310 302648 159200
rect 302516 155304 302568 155310
rect 302516 155246 302568 155252
rect 302608 155304 302660 155310
rect 302608 155246 302660 155252
rect 301596 155168 301648 155174
rect 301596 155110 301648 155116
rect 300676 155100 300728 155106
rect 300676 155042 300728 155048
rect 300860 154488 300912 154494
rect 300860 154430 300912 154436
rect 300872 153950 300900 154430
rect 301412 154420 301464 154426
rect 301412 154362 301464 154368
rect 300860 153944 300912 153950
rect 300860 153886 300912 153892
rect 300860 152516 300912 152522
rect 300860 152458 300912 152464
rect 300872 151994 300900 152458
rect 301424 151994 301452 154362
rect 302240 153536 302292 153542
rect 302240 153478 302292 153484
rect 302252 151994 302280 153478
rect 302528 152130 302556 155246
rect 303632 154698 303660 159200
rect 303528 154692 303580 154698
rect 303528 154634 303580 154640
rect 303620 154692 303672 154698
rect 303620 154634 303672 154640
rect 303540 154578 303568 154634
rect 304552 154630 304580 159200
rect 305564 155786 305592 159200
rect 305000 155780 305052 155786
rect 305000 155722 305052 155728
rect 305552 155780 305604 155786
rect 305552 155722 305604 155728
rect 303804 154624 303856 154630
rect 303540 154550 303660 154578
rect 303804 154566 303856 154572
rect 304540 154624 304592 154630
rect 304540 154566 304592 154572
rect 302528 152102 302648 152130
rect 302620 151994 302648 152102
rect 303632 151994 303660 154550
rect 303816 153338 303844 154566
rect 305012 154290 305040 155722
rect 305920 155712 305972 155718
rect 305920 155654 305972 155660
rect 303988 154284 304040 154290
rect 303988 154226 304040 154232
rect 305000 154284 305052 154290
rect 305000 154226 305052 154232
rect 303804 153332 303856 153338
rect 303804 153274 303856 153280
rect 304000 151994 304028 154226
rect 305276 153808 305328 153814
rect 305276 153750 305328 153756
rect 304632 153400 304684 153406
rect 304632 153342 304684 153348
rect 304644 151994 304672 153342
rect 305288 151994 305316 153750
rect 305932 151994 305960 155654
rect 306484 155446 306512 159200
rect 306472 155440 306524 155446
rect 306472 155382 306524 155388
rect 307496 155378 307524 159200
rect 308508 155514 308536 159200
rect 308404 155508 308456 155514
rect 308404 155450 308456 155456
rect 308496 155508 308548 155514
rect 308496 155450 308548 155456
rect 307484 155372 307536 155378
rect 307484 155314 307536 155320
rect 307668 154896 307720 154902
rect 307668 154838 307720 154844
rect 306656 154216 306708 154222
rect 306656 154158 306708 154164
rect 306668 151994 306696 154158
rect 307300 153876 307352 153882
rect 307300 153818 307352 153824
rect 307312 151994 307340 153818
rect 307680 153406 307708 154838
rect 308416 154222 308444 155450
rect 309428 155106 309456 159200
rect 309324 155100 309376 155106
rect 309324 155042 309376 155048
rect 309416 155100 309468 155106
rect 309416 155042 309468 155048
rect 308588 154828 308640 154834
rect 308588 154770 308640 154776
rect 308404 154216 308456 154222
rect 308404 154158 308456 154164
rect 307668 153400 307720 153406
rect 307668 153342 307720 153348
rect 307944 153332 307996 153338
rect 307944 153274 307996 153280
rect 307956 151994 307984 153274
rect 308600 151994 308628 154770
rect 309336 154154 309364 155042
rect 310440 154834 310468 159200
rect 311256 155848 311308 155854
rect 311256 155790 311308 155796
rect 310428 154828 310480 154834
rect 310428 154770 310480 154776
rect 311164 154624 311216 154630
rect 311164 154566 311216 154572
rect 309876 154352 309928 154358
rect 309876 154294 309928 154300
rect 309232 154148 309284 154154
rect 309232 154090 309284 154096
rect 309324 154148 309376 154154
rect 309324 154090 309376 154096
rect 309244 151994 309272 154090
rect 309888 151994 309916 154294
rect 311176 153882 311204 154566
rect 311164 153876 311216 153882
rect 311164 153818 311216 153824
rect 310520 153400 310572 153406
rect 310520 153342 310572 153348
rect 310532 151994 310560 153342
rect 311268 151994 311296 155790
rect 311360 154902 311388 159200
rect 311900 155576 311952 155582
rect 311900 155518 311952 155524
rect 311348 154896 311400 154902
rect 311348 154838 311400 154844
rect 311912 151994 311940 155518
rect 312372 154630 312400 159200
rect 313292 155582 313320 159200
rect 313740 155916 313792 155922
rect 313740 155858 313792 155864
rect 313372 155712 313424 155718
rect 313372 155654 313424 155660
rect 313280 155576 313332 155582
rect 313280 155518 313332 155524
rect 312360 154624 312412 154630
rect 312360 154566 312412 154572
rect 313280 154012 313332 154018
rect 313280 153954 313332 153960
rect 312452 153944 312504 153950
rect 312452 153886 312504 153892
rect 312464 151994 312492 153886
rect 313292 151994 313320 153954
rect 313384 153270 313412 155654
rect 313372 153264 313424 153270
rect 313372 153206 313424 153212
rect 313752 151994 313780 155858
rect 314304 155718 314332 159200
rect 315316 155854 315344 159200
rect 316236 155922 316264 159200
rect 316224 155916 316276 155922
rect 316224 155858 316276 155864
rect 315304 155848 315356 155854
rect 315304 155790 315356 155796
rect 314292 155712 314344 155718
rect 314292 155654 314344 155660
rect 317248 155650 317276 159200
rect 317052 155644 317104 155650
rect 317052 155586 317104 155592
rect 317236 155644 317288 155650
rect 317236 155586 317288 155592
rect 316408 155032 316460 155038
rect 316408 154974 316460 154980
rect 314752 154760 314804 154766
rect 314752 154702 314804 154708
rect 314660 154080 314712 154086
rect 314660 154022 314712 154028
rect 314672 151994 314700 154022
rect 314764 153338 314792 154702
rect 315028 154284 315080 154290
rect 315028 154226 315080 154232
rect 314752 153332 314804 153338
rect 314752 153274 314804 153280
rect 315040 151994 315068 154226
rect 316040 153264 316092 153270
rect 316040 153206 316092 153212
rect 316052 151994 316080 153206
rect 316420 151994 316448 154974
rect 317064 151994 317092 155586
rect 318168 155174 318196 159200
rect 318984 155236 319036 155242
rect 318984 155178 319036 155184
rect 317328 155168 317380 155174
rect 317328 155110 317380 155116
rect 318156 155168 318208 155174
rect 318156 155110 318208 155116
rect 317340 153542 317368 155110
rect 318708 154692 318760 154698
rect 318708 154634 318760 154640
rect 317696 154216 317748 154222
rect 317696 154158 317748 154164
rect 317328 153536 317380 153542
rect 317328 153478 317380 153484
rect 317708 151994 317736 154158
rect 318340 153332 318392 153338
rect 318340 153274 318392 153280
rect 318352 151994 318380 153274
rect 318720 153270 318748 154634
rect 318708 153264 318760 153270
rect 318708 153206 318760 153212
rect 318996 151994 319024 155178
rect 319180 154766 319208 159200
rect 319628 154964 319680 154970
rect 319628 154906 319680 154912
rect 319168 154760 319220 154766
rect 319168 154702 319220 154708
rect 319640 151994 319668 154906
rect 320192 154698 320220 159200
rect 321112 155038 321140 159200
rect 321652 155304 321704 155310
rect 321652 155246 321704 155252
rect 321100 155032 321152 155038
rect 321100 154974 321152 154980
rect 321560 154896 321612 154902
rect 321560 154838 321612 154844
rect 320180 154692 320232 154698
rect 320180 154634 320232 154640
rect 320272 154148 320324 154154
rect 320272 154090 320324 154096
rect 320284 151994 320312 154090
rect 321572 153542 321600 154838
rect 320916 153536 320968 153542
rect 320916 153478 320968 153484
rect 321560 153536 321612 153542
rect 321560 153478 321612 153484
rect 320928 151994 320956 153478
rect 321664 151994 321692 155246
rect 322124 154970 322152 159200
rect 323044 155242 323072 159200
rect 323492 155780 323544 155786
rect 323492 155722 323544 155728
rect 323032 155236 323084 155242
rect 323032 155178 323084 155184
rect 323216 155100 323268 155106
rect 323216 155042 323268 155048
rect 322112 154964 322164 154970
rect 322112 154906 322164 154912
rect 323032 154828 323084 154834
rect 323032 154770 323084 154776
rect 322940 154624 322992 154630
rect 322940 154566 322992 154572
rect 322952 153610 322980 154566
rect 322940 153604 322992 153610
rect 322940 153546 322992 153552
rect 323044 153474 323072 154770
rect 323124 153876 323176 153882
rect 323124 153818 323176 153824
rect 323032 153468 323084 153474
rect 323032 153410 323084 153416
rect 322204 153264 322256 153270
rect 322204 153206 322256 153212
rect 322216 151994 322244 153206
rect 323136 151994 323164 153818
rect 323228 153406 323256 155042
rect 323216 153400 323268 153406
rect 323216 153342 323268 153348
rect 323504 151994 323532 155722
rect 324056 154834 324084 159200
rect 324412 155508 324464 155514
rect 324412 155450 324464 155456
rect 324228 155440 324280 155446
rect 324228 155382 324280 155388
rect 324136 155372 324188 155378
rect 324136 155314 324188 155320
rect 324044 154828 324096 154834
rect 324044 154770 324096 154776
rect 324148 153678 324176 155314
rect 324136 153672 324188 153678
rect 324136 153614 324188 153620
rect 324240 153218 324268 155382
rect 324424 153270 324452 155450
rect 325068 155378 325096 159200
rect 325988 155514 326016 159200
rect 325976 155508 326028 155514
rect 325976 155450 326028 155456
rect 325056 155372 325108 155378
rect 325056 155314 325108 155320
rect 327000 155310 327028 159200
rect 327920 155446 327948 159200
rect 328932 155922 328960 159200
rect 328460 155916 328512 155922
rect 328460 155858 328512 155864
rect 328920 155916 328972 155922
rect 328920 155858 328972 155864
rect 327908 155440 327960 155446
rect 327908 155382 327960 155388
rect 326988 155304 327040 155310
rect 326988 155246 327040 155252
rect 328472 153950 328500 155858
rect 329656 155848 329708 155854
rect 329656 155790 329708 155796
rect 329380 155712 329432 155718
rect 329380 155654 329432 155660
rect 328736 155576 328788 155582
rect 328736 155518 328788 155524
rect 328460 153944 328512 153950
rect 328460 153886 328512 153892
rect 324872 153672 324924 153678
rect 324872 153614 324924 153620
rect 324412 153264 324464 153270
rect 324240 153190 324360 153218
rect 324412 153206 324464 153212
rect 324332 151994 324360 153190
rect 324884 151994 324912 153614
rect 328092 153604 328144 153610
rect 328092 153546 328144 153552
rect 327448 153536 327500 153542
rect 327448 153478 327500 153484
rect 327080 153468 327132 153474
rect 327080 153410 327132 153416
rect 326160 153400 326212 153406
rect 326160 153342 326212 153348
rect 325792 153264 325844 153270
rect 325792 153206 325844 153212
rect 325804 151994 325832 153206
rect 326172 151994 326200 153342
rect 327092 151994 327120 153410
rect 327460 151994 327488 153478
rect 328104 151994 328132 153546
rect 328748 151994 328776 155518
rect 329392 151994 329420 155654
rect 329668 153218 329696 155790
rect 329944 155582 329972 159200
rect 330864 155854 330892 159200
rect 330852 155848 330904 155854
rect 330852 155790 330904 155796
rect 331876 155786 331904 159200
rect 331864 155780 331916 155786
rect 331864 155722 331916 155728
rect 331312 155644 331364 155650
rect 331312 155586 331364 155592
rect 329932 155576 329984 155582
rect 329932 155518 329984 155524
rect 329748 155168 329800 155174
rect 329748 155110 329800 155116
rect 329760 153542 329788 155110
rect 330668 153944 330720 153950
rect 330668 153886 330720 153892
rect 329748 153536 329800 153542
rect 329748 153478 329800 153484
rect 329668 153190 329972 153218
rect 329944 151994 329972 153190
rect 330680 151994 330708 153886
rect 331324 151994 331352 155586
rect 332796 155174 332824 159200
rect 333808 155650 333836 159200
rect 334820 155922 334848 159200
rect 334348 155916 334400 155922
rect 334348 155858 334400 155864
rect 334808 155916 334860 155922
rect 334808 155858 334860 155864
rect 333796 155644 333848 155650
rect 333796 155586 333848 155592
rect 334072 155236 334124 155242
rect 334072 155178 334124 155184
rect 332784 155168 332836 155174
rect 332784 155110 332836 155116
rect 332324 155032 332376 155038
rect 332324 154974 332376 154980
rect 331956 153536 332008 153542
rect 331956 153478 332008 153484
rect 331968 151994 331996 153478
rect 332336 153406 332364 154974
rect 333888 154964 333940 154970
rect 333888 154906 333940 154912
rect 332600 154556 332652 154562
rect 332600 154498 332652 154504
rect 332324 153400 332376 153406
rect 332324 153342 332376 153348
rect 332612 151994 332640 154498
rect 333244 154488 333296 154494
rect 333244 154430 333296 154436
rect 333256 151994 333284 154430
rect 333900 153474 333928 154906
rect 333980 154828 334032 154834
rect 333980 154770 334032 154776
rect 333992 153542 334020 154770
rect 333980 153536 334032 153542
rect 333980 153478 334032 153484
rect 333888 153468 333940 153474
rect 333888 153410 333940 153416
rect 333980 153400 334032 153406
rect 333980 153342 334032 153348
rect 333992 151994 334020 153342
rect 334084 153270 334112 155178
rect 334360 153950 334388 155858
rect 335740 155582 335768 159200
rect 336556 155848 336608 155854
rect 336556 155790 336608 155796
rect 335636 155576 335688 155582
rect 335636 155518 335688 155524
rect 335728 155576 335780 155582
rect 335728 155518 335780 155524
rect 334348 153944 334400 153950
rect 334348 153886 334400 153892
rect 335648 153746 335676 155518
rect 335636 153740 335688 153746
rect 335636 153682 335688 153688
rect 335912 153536 335964 153542
rect 335912 153478 335964 153484
rect 334624 153468 334676 153474
rect 334624 153410 334676 153416
rect 334072 153264 334124 153270
rect 334072 153206 334124 153212
rect 334636 151994 334664 153410
rect 335452 153264 335504 153270
rect 335452 153206 335504 153212
rect 335464 151994 335492 153206
rect 335924 151994 335952 153478
rect 336568 153406 336596 155790
rect 336648 155372 336700 155378
rect 336648 155314 336700 155320
rect 336556 153400 336608 153406
rect 336556 153342 336608 153348
rect 336660 153218 336688 155314
rect 336752 154630 336780 159200
rect 337672 155514 337700 159200
rect 337936 155780 337988 155786
rect 337936 155722 337988 155728
rect 337200 155508 337252 155514
rect 337200 155450 337252 155456
rect 337660 155508 337712 155514
rect 337660 155450 337712 155456
rect 336740 154624 336792 154630
rect 336740 154566 336792 154572
rect 336660 153190 336780 153218
rect 336752 151994 336780 153190
rect 337212 151994 337240 155450
rect 337948 153814 337976 155722
rect 338488 155440 338540 155446
rect 338488 155382 338540 155388
rect 338028 155304 338080 155310
rect 338028 155246 338080 155252
rect 337936 153808 337988 153814
rect 337936 153750 337988 153756
rect 338040 153218 338068 155246
rect 338040 153190 338160 153218
rect 338132 151994 338160 153190
rect 338500 151994 338528 155382
rect 338684 155242 338712 159200
rect 338948 155644 339000 155650
rect 338948 155586 339000 155592
rect 338672 155236 338724 155242
rect 338672 155178 338724 155184
rect 338580 155168 338632 155174
rect 338580 155110 338632 155116
rect 338592 153542 338620 155110
rect 338960 153678 338988 155586
rect 339696 154698 339724 159200
rect 340236 155916 340288 155922
rect 340236 155858 340288 155864
rect 339684 154692 339736 154698
rect 339684 154634 339736 154640
rect 340248 153950 340276 155858
rect 340616 154766 340644 159200
rect 340972 155576 341024 155582
rect 340972 155518 341024 155524
rect 340604 154760 340656 154766
rect 340604 154702 340656 154708
rect 340984 154494 341012 155518
rect 341628 154834 341656 159200
rect 342548 155650 342576 159200
rect 342536 155644 342588 155650
rect 342536 155586 342588 155592
rect 342536 155508 342588 155514
rect 342536 155450 342588 155456
rect 341616 154828 341668 154834
rect 341616 154770 341668 154776
rect 340972 154488 341024 154494
rect 340972 154430 341024 154436
rect 339132 153944 339184 153950
rect 339132 153886 339184 153892
rect 340236 153944 340288 153950
rect 340236 153886 340288 153892
rect 338948 153672 339000 153678
rect 338948 153614 339000 153620
rect 338580 153536 338632 153542
rect 338580 153478 338632 153484
rect 339144 151994 339172 153886
rect 341064 153808 341116 153814
rect 341064 153750 341116 153756
rect 339776 153740 339828 153746
rect 339776 153682 339828 153688
rect 339788 151994 339816 153682
rect 340420 153400 340472 153406
rect 340420 153342 340472 153348
rect 340432 151994 340460 153342
rect 341076 151994 341104 153750
rect 342352 153672 342404 153678
rect 342352 153614 342404 153620
rect 341708 153536 341760 153542
rect 341708 153478 341760 153484
rect 341720 151994 341748 153478
rect 342364 151994 342392 153614
rect 342548 153406 342576 155450
rect 343560 155174 343588 159200
rect 344572 155514 344600 159200
rect 345492 155582 345520 159200
rect 345480 155576 345532 155582
rect 345480 155518 345532 155524
rect 344560 155508 344612 155514
rect 344560 155450 344612 155456
rect 343640 155236 343692 155242
rect 343640 155178 343692 155184
rect 343548 155168 343600 155174
rect 343548 155110 343600 155116
rect 342996 153944 343048 153950
rect 342996 153886 343048 153892
rect 342536 153400 342588 153406
rect 342536 153342 342588 153348
rect 343008 151994 343036 153886
rect 343652 153338 343680 155178
rect 346308 154692 346360 154698
rect 346308 154634 346360 154640
rect 344376 154556 344428 154562
rect 344376 154498 344428 154504
rect 343732 154488 343784 154494
rect 343732 154430 343784 154436
rect 343640 153332 343692 153338
rect 343640 153274 343692 153280
rect 343744 151994 343772 154430
rect 344388 151994 344416 154498
rect 345204 153400 345256 153406
rect 345204 153342 345256 153348
rect 345216 151994 345244 153342
rect 345664 153332 345716 153338
rect 345664 153274 345716 153280
rect 345676 151994 345704 153274
rect 346320 153218 346348 154634
rect 346504 154630 346532 159200
rect 347424 159174 347544 159200
rect 347596 155576 347648 155582
rect 347596 155518 347648 155524
rect 347504 154828 347556 154834
rect 347504 154770 347556 154776
rect 346492 154624 346544 154630
rect 346492 154566 346544 154572
rect 347044 154556 347096 154562
rect 347044 154498 347096 154504
rect 346320 153190 346440 153218
rect 346412 151994 346440 153190
rect 347056 151994 347084 154498
rect 347516 153252 347544 154770
rect 347608 154222 347636 155518
rect 347700 154574 347728 159310
rect 348422 159200 348478 160000
rect 349342 159200 349398 160000
rect 350354 159200 350410 160000
rect 351366 159200 351422 160000
rect 352286 159200 352342 160000
rect 353298 159200 353354 160000
rect 354218 159200 354274 160000
rect 355230 159200 355286 160000
rect 356242 159200 356298 160000
rect 357162 159200 357218 160000
rect 358174 159200 358230 160000
rect 359094 159200 359150 160000
rect 360106 159200 360162 160000
rect 361118 159200 361174 160000
rect 362038 159200 362094 160000
rect 363050 159200 363106 160000
rect 363970 159200 364026 160000
rect 364982 159200 365038 160000
rect 365994 159200 366050 160000
rect 366914 159200 366970 160000
rect 367926 159200 367982 160000
rect 368846 159200 368902 160000
rect 369858 159200 369914 160000
rect 370870 159200 370926 160000
rect 371790 159200 371846 160000
rect 372802 159200 372858 160000
rect 373722 159200 373778 160000
rect 374734 159200 374790 160000
rect 375746 159200 375802 160000
rect 376666 159200 376722 160000
rect 377678 159200 377734 160000
rect 378598 159200 378654 160000
rect 379610 159200 379666 160000
rect 380622 159200 380678 160000
rect 381542 159200 381598 160000
rect 382554 159200 382610 160000
rect 383474 159200 383530 160000
rect 384486 159200 384542 160000
rect 385498 159200 385554 160000
rect 386418 159200 386474 160000
rect 387430 159200 387486 160000
rect 388350 159200 388406 160000
rect 389362 159200 389418 160000
rect 390282 159200 390338 160000
rect 391294 159200 391350 160000
rect 392306 159200 392362 160000
rect 393226 159200 393282 160000
rect 394238 159200 394294 160000
rect 395158 159200 395214 160000
rect 396170 159200 396226 160000
rect 397182 159200 397238 160000
rect 398102 159200 398158 160000
rect 398852 159310 399064 159338
rect 348240 155644 348292 155650
rect 348240 155586 348292 155592
rect 347700 154546 347820 154574
rect 347596 154216 347648 154222
rect 347596 154158 347648 154164
rect 347792 153814 347820 154546
rect 347780 153808 347832 153814
rect 347780 153750 347832 153756
rect 347516 153224 347820 153252
rect 347792 151994 347820 153224
rect 348252 151994 348280 155586
rect 348436 154630 348464 159200
rect 349068 155168 349120 155174
rect 349068 155110 349120 155116
rect 348424 154624 348476 154630
rect 348424 154566 348476 154572
rect 349080 153218 349108 155110
rect 349356 154630 349384 159200
rect 349528 155508 349580 155514
rect 349528 155450 349580 155456
rect 349344 154624 349396 154630
rect 349344 154566 349396 154572
rect 349080 153190 349200 153218
rect 349172 151994 349200 153190
rect 349540 151994 349568 155450
rect 350368 154630 350396 159200
rect 351380 154630 351408 159200
rect 352300 154698 352328 159200
rect 353312 155922 353340 159200
rect 353300 155916 353352 155922
rect 353300 155858 353352 155864
rect 354232 155854 354260 159200
rect 354220 155848 354272 155854
rect 354220 155790 354272 155796
rect 355244 155038 355272 159200
rect 355416 155916 355468 155922
rect 355416 155858 355468 155864
rect 355232 155032 355284 155038
rect 355232 154974 355284 154980
rect 352288 154692 352340 154698
rect 352288 154634 352340 154640
rect 353392 154692 353444 154698
rect 353392 154634 353444 154640
rect 350356 154624 350408 154630
rect 350356 154566 350408 154572
rect 351368 154624 351420 154630
rect 351368 154566 351420 154572
rect 352840 154420 352892 154426
rect 352840 154362 352892 154368
rect 352104 154352 352156 154358
rect 352104 154294 352156 154300
rect 350816 154284 350868 154290
rect 350816 154226 350868 154232
rect 350172 154216 350224 154222
rect 350172 154158 350224 154164
rect 350184 151994 350212 154158
rect 350828 151994 350856 154226
rect 351460 153808 351512 153814
rect 351460 153750 351512 153756
rect 351472 151994 351500 153750
rect 352116 151994 352144 154294
rect 352852 151994 352880 154362
rect 353404 153270 353432 154634
rect 354128 154556 354180 154562
rect 354128 154498 354180 154504
rect 353484 154488 353536 154494
rect 353484 154430 353536 154436
rect 353392 153264 353444 153270
rect 353392 153206 353444 153212
rect 353496 151994 353524 154430
rect 354140 151994 354168 154498
rect 354864 153264 354916 153270
rect 354864 153206 354916 153212
rect 354876 151994 354904 153206
rect 355428 151994 355456 155858
rect 355968 155848 356020 155854
rect 355968 155790 356020 155796
rect 355980 153218 356008 155790
rect 356256 155582 356284 159200
rect 356244 155576 356296 155582
rect 356244 155518 356296 155524
rect 356704 155032 356756 155038
rect 356704 154974 356756 154980
rect 355980 153190 356100 153218
rect 356072 151994 356100 153190
rect 356716 151994 356744 154974
rect 357176 154970 357204 159200
rect 358188 155582 358216 159200
rect 357440 155576 357492 155582
rect 357440 155518 357492 155524
rect 358176 155576 358228 155582
rect 358176 155518 358228 155524
rect 358820 155576 358872 155582
rect 358820 155518 358872 155524
rect 357164 154964 357216 154970
rect 357164 154906 357216 154912
rect 357452 151994 357480 155518
rect 357992 154964 358044 154970
rect 357992 154906 358044 154912
rect 358004 151994 358032 154906
rect 358832 151994 358860 155518
rect 359108 151994 359136 159200
rect 360120 154578 360148 159200
rect 360120 154550 360240 154578
rect 360212 151994 360240 154550
rect 361132 151994 361160 159200
rect 362052 154562 362080 159200
rect 363064 154562 363092 159200
rect 361488 154556 361540 154562
rect 361488 154498 361540 154504
rect 362040 154556 362092 154562
rect 362040 154498 362092 154504
rect 362592 154556 362644 154562
rect 362592 154498 362644 154504
rect 363052 154556 363104 154562
rect 363052 154498 363104 154504
rect 256752 151988 256864 151994
rect 256700 151982 256864 151988
rect 256712 151966 256864 151982
rect 257172 151966 257508 151994
rect 258092 151966 258152 151994
rect 258460 151966 258796 151994
rect 259104 151966 259440 151994
rect 259840 151966 260176 151994
rect 260484 151966 260820 151994
rect 261128 151966 261464 151994
rect 261772 151966 262108 151994
rect 262416 151966 262752 151994
rect 263060 151966 263396 151994
rect 263704 151966 264040 151994
rect 264348 151966 264684 151994
rect 264992 151966 265328 151994
rect 265636 151966 265972 151994
rect 266372 151966 266616 151994
rect 266924 151966 267260 151994
rect 267844 151966 267904 151994
rect 268212 151966 268548 151994
rect 269132 151966 269284 151994
rect 269592 151966 269928 151994
rect 270512 151966 270572 151994
rect 270880 151966 271216 151994
rect 271524 151966 271860 151994
rect 272168 151966 272504 151994
rect 272812 151966 273148 151994
rect 273456 151966 273792 151994
rect 274100 151966 274436 151994
rect 274744 151966 275080 151994
rect 275388 151966 275724 151994
rect 276032 151966 276368 151994
rect 276676 151966 277012 151994
rect 277504 151966 277656 151994
rect 277964 151966 278300 151994
rect 278792 151966 279036 151994
rect 279344 151966 279680 151994
rect 280172 151966 280324 151994
rect 280632 151966 280968 151994
rect 281552 151966 281612 151994
rect 281920 151966 282256 151994
rect 282564 151966 282900 151994
rect 283208 151966 283544 151994
rect 284036 151966 284188 151994
rect 284496 151966 284832 151994
rect 285140 151966 285476 151994
rect 285784 151966 286120 151994
rect 286428 151966 286764 151994
rect 287256 151966 287408 151994
rect 287808 151966 288144 151994
rect 288452 151966 288788 151994
rect 289096 151966 289432 151994
rect 289832 151966 290076 151994
rect 290384 151966 290720 151994
rect 291212 151966 291364 151994
rect 291672 151966 292008 151994
rect 292592 151966 292652 151994
rect 292960 151966 293296 151994
rect 293604 151966 293940 151994
rect 294248 151966 294584 151994
rect 294800 151966 295228 151994
rect 295536 151966 295872 151994
rect 296180 151966 296516 151994
rect 297008 151966 297252 151994
rect 297560 151966 297896 151994
rect 298204 151966 298540 151994
rect 298848 151966 299184 151994
rect 299492 151966 299828 151994
rect 300136 151966 300472 151994
rect 300872 151966 301116 151994
rect 301424 151966 301760 151994
rect 302252 151966 302404 151994
rect 302620 151966 303048 151994
rect 303632 151966 303692 151994
rect 304000 151966 304336 151994
rect 304644 151966 304980 151994
rect 305288 151966 305624 151994
rect 305932 151966 306268 151994
rect 306668 151966 307004 151994
rect 307312 151966 307648 151994
rect 307956 151966 308292 151994
rect 308600 151966 308936 151994
rect 309244 151966 309580 151994
rect 309888 151966 310224 151994
rect 310532 151966 310868 151994
rect 311268 151966 311512 151994
rect 311912 151966 312156 151994
rect 312464 151966 312800 151994
rect 313292 151966 313444 151994
rect 313752 151966 314088 151994
rect 314672 151966 314732 151994
rect 315040 151966 315376 151994
rect 316052 151966 316112 151994
rect 316420 151966 316756 151994
rect 317064 151966 317400 151994
rect 317708 151966 318044 151994
rect 318352 151966 318688 151994
rect 318996 151966 319332 151994
rect 319640 151966 319976 151994
rect 320284 151966 320620 151994
rect 320928 151966 321264 151994
rect 321664 151966 321908 151994
rect 322216 151966 322552 151994
rect 323136 151966 323196 151994
rect 323504 151966 323840 151994
rect 324332 151966 324484 151994
rect 324884 151966 325220 151994
rect 325804 151966 325864 151994
rect 326172 151966 326508 151994
rect 327092 151966 327152 151994
rect 327460 151966 327796 151994
rect 328104 151966 328440 151994
rect 328748 151966 329084 151994
rect 329392 151966 329728 151994
rect 329944 151966 330372 151994
rect 330680 151966 331016 151994
rect 331324 151966 331660 151994
rect 331968 151966 332304 151994
rect 332612 151966 332948 151994
rect 333256 151966 333592 151994
rect 333992 151966 334328 151994
rect 334636 151966 334972 151994
rect 335464 151966 335616 151994
rect 335924 151966 336260 151994
rect 336752 151966 336904 151994
rect 337212 151966 337548 151994
rect 338132 151966 338192 151994
rect 338500 151966 338836 151994
rect 339144 151966 339480 151994
rect 339788 151966 340124 151994
rect 340432 151966 340768 151994
rect 341076 151966 341412 151994
rect 341720 151966 342056 151994
rect 342364 151966 342700 151994
rect 343008 151966 343344 151994
rect 343744 151966 344080 151994
rect 344388 151966 344724 151994
rect 345216 151966 345368 151994
rect 345676 151966 346012 151994
rect 346412 151966 346656 151994
rect 347056 151966 347300 151994
rect 347792 151966 347944 151994
rect 348252 151966 348588 151994
rect 349172 151966 349232 151994
rect 349540 151966 349876 151994
rect 350184 151966 350520 151994
rect 350828 151966 351164 151994
rect 351472 151966 351808 151994
rect 352116 151966 352452 151994
rect 352852 151966 353188 151994
rect 353496 151966 353832 151994
rect 354140 151966 354476 151994
rect 354876 151966 355120 151994
rect 355428 151966 355764 151994
rect 356072 151966 356408 151994
rect 356716 151966 357052 151994
rect 357452 151966 357696 151994
rect 358004 151966 358340 151994
rect 358832 151966 358984 151994
rect 359108 151966 359628 151994
rect 360212 151966 360272 151994
rect 360916 151966 361160 151994
rect 361500 151994 361528 154498
rect 362604 151994 362632 154498
rect 363984 154494 364012 159200
rect 362868 154488 362920 154494
rect 362868 154430 362920 154436
rect 363972 154488 364024 154494
rect 363972 154430 364024 154436
rect 361500 151966 361560 151994
rect 362296 151966 362632 151994
rect 362880 151994 362908 154430
rect 364156 153332 364208 153338
rect 364156 153274 364208 153280
rect 363880 153264 363932 153270
rect 363880 153206 363932 153212
rect 363892 151994 363920 153206
rect 362880 151966 362940 151994
rect 363584 151966 363920 151994
rect 238944 151914 238996 151920
rect 127532 151836 127584 151842
rect 127532 151778 127584 151784
rect 204536 151836 204884 151842
rect 204588 151830 204884 151836
rect 211068 151836 211120 151842
rect 204536 151778 204588 151784
rect 213992 151830 214144 151858
rect 246948 151904 247000 151910
rect 364168 151858 364196 153274
rect 364996 153270 365024 159200
rect 366008 154970 366036 159200
rect 365260 154964 365312 154970
rect 365260 154906 365312 154912
rect 365996 154964 366048 154970
rect 365996 154906 366048 154912
rect 365168 153468 365220 153474
rect 365168 153410 365220 153416
rect 364984 153264 365036 153270
rect 364984 153206 365036 153212
rect 365180 151994 365208 153410
rect 365272 153338 365300 154906
rect 365628 154556 365680 154562
rect 365628 154498 365680 154504
rect 366456 154556 366508 154562
rect 366456 154498 366508 154504
rect 365260 153332 365312 153338
rect 365260 153274 365312 153280
rect 365640 151994 365668 154498
rect 366468 151994 366496 154498
rect 366928 153474 366956 159200
rect 367940 154630 367968 159200
rect 368860 154630 368888 159200
rect 367928 154624 367980 154630
rect 367928 154566 367980 154572
rect 368848 154624 368900 154630
rect 368848 154566 368900 154572
rect 369872 154494 369900 159200
rect 370884 154630 370912 159200
rect 370872 154624 370924 154630
rect 370872 154566 370924 154572
rect 367008 154488 367060 154494
rect 367008 154430 367060 154436
rect 369860 154488 369912 154494
rect 369860 154430 369912 154436
rect 366916 153468 366968 153474
rect 366916 153410 366968 153416
rect 367020 151994 367048 154430
rect 367744 154420 367796 154426
rect 367744 154362 367796 154368
rect 367756 151994 367784 154362
rect 371804 154358 371832 159200
rect 368388 154352 368440 154358
rect 368388 154294 368440 154300
rect 371792 154352 371844 154358
rect 371792 154294 371844 154300
rect 368400 151994 368428 154294
rect 369676 154284 369728 154290
rect 369676 154226 369728 154232
rect 369032 154012 369084 154018
rect 369032 153954 369084 153960
rect 369044 151994 369072 153954
rect 369688 151994 369716 154226
rect 372344 154216 372396 154222
rect 372344 154158 372396 154164
rect 370964 153536 371016 153542
rect 370964 153478 371016 153484
rect 370320 153468 370372 153474
rect 370320 153410 370372 153416
rect 370332 151994 370360 153410
rect 370976 151994 371004 153478
rect 371608 153332 371660 153338
rect 371608 153274 371660 153280
rect 371620 151994 371648 153274
rect 372356 151994 372384 154158
rect 372816 154018 372844 159200
rect 372988 154488 373040 154494
rect 372988 154430 373040 154436
rect 372804 154012 372856 154018
rect 372804 153954 372856 153960
rect 373000 151994 373028 154430
rect 373736 154290 373764 159200
rect 373724 154284 373776 154290
rect 373724 154226 373776 154232
rect 373908 154012 373960 154018
rect 373908 153954 373960 153960
rect 373632 153876 373684 153882
rect 373632 153818 373684 153824
rect 373644 151994 373672 153818
rect 364872 151966 365208 151994
rect 365516 151966 365668 151994
rect 366160 151966 366496 151994
rect 366804 151966 367048 151994
rect 367448 151966 367784 151994
rect 368092 151966 368428 151994
rect 368736 151966 369072 151994
rect 369380 151966 369716 151994
rect 370024 151966 370360 151994
rect 370668 151966 371004 151994
rect 371312 151966 371648 151994
rect 372048 151966 372384 151994
rect 372692 151966 373028 151994
rect 373336 151966 373672 151994
rect 373920 151994 373948 153954
rect 374748 153474 374776 159200
rect 374920 154556 374972 154562
rect 374920 154498 374972 154504
rect 374736 153468 374788 153474
rect 374736 153410 374788 153416
rect 374932 151994 374960 154498
rect 375196 154420 375248 154426
rect 375196 154362 375248 154368
rect 373920 151966 373980 151994
rect 374624 151966 374960 151994
rect 375208 151858 375236 154362
rect 375760 153542 375788 159200
rect 376208 154352 376260 154358
rect 376208 154294 376260 154300
rect 375748 153536 375800 153542
rect 375748 153478 375800 153484
rect 376220 151994 376248 154294
rect 376484 153672 376536 153678
rect 376484 153614 376536 153620
rect 375912 151966 376248 151994
rect 376496 151858 376524 153614
rect 376680 153338 376708 159200
rect 377692 154222 377720 159200
rect 378140 155576 378192 155582
rect 378140 155518 378192 155524
rect 377680 154216 377732 154222
rect 377680 154158 377732 154164
rect 378152 154018 378180 155518
rect 378612 154494 378640 159200
rect 379624 154714 379652 159200
rect 379704 155644 379756 155650
rect 379704 155586 379756 155592
rect 379440 154686 379652 154714
rect 378600 154488 378652 154494
rect 378600 154430 378652 154436
rect 378140 154012 378192 154018
rect 378140 153954 378192 153960
rect 377496 153944 377548 153950
rect 377496 153886 377548 153892
rect 376668 153332 376720 153338
rect 376668 153274 376720 153280
rect 377508 151994 377536 153886
rect 379440 153882 379468 154686
rect 379716 154426 379744 155586
rect 380636 155582 380664 159200
rect 380624 155576 380676 155582
rect 380624 155518 380676 155524
rect 380900 155508 380952 155514
rect 380900 155450 380952 155456
rect 379704 154420 379756 154426
rect 379704 154362 379756 154368
rect 379428 153876 379480 153882
rect 379428 153818 379480 153824
rect 380912 153678 380940 155450
rect 381556 154630 381584 159200
rect 382372 155916 382424 155922
rect 382372 155858 382424 155864
rect 382280 155236 382332 155242
rect 382280 155178 382332 155184
rect 381544 154624 381596 154630
rect 381544 154566 381596 154572
rect 382096 154556 382148 154562
rect 382096 154498 382148 154504
rect 381452 154148 381504 154154
rect 381452 154090 381504 154096
rect 380900 153672 380952 153678
rect 380900 153614 380952 153620
rect 380072 153604 380124 153610
rect 380072 153546 380124 153552
rect 378784 153536 378836 153542
rect 378784 153478 378836 153484
rect 378048 153468 378100 153474
rect 378048 153410 378100 153416
rect 378060 151994 378088 153410
rect 378796 151994 378824 153478
rect 379428 153400 379480 153406
rect 379428 153342 379480 153348
rect 379440 151994 379468 153342
rect 380084 151994 380112 153546
rect 380716 153264 380768 153270
rect 380716 153206 380768 153212
rect 380728 151994 380756 153206
rect 381464 151994 381492 154090
rect 382108 151994 382136 154498
rect 382292 153474 382320 155178
rect 382384 153950 382412 155858
rect 382568 155650 382596 159200
rect 382556 155644 382608 155650
rect 382556 155586 382608 155592
rect 383488 154630 383516 159200
rect 384500 155514 384528 159200
rect 385512 155922 385540 159200
rect 385500 155916 385552 155922
rect 385500 155858 385552 155864
rect 385500 155780 385552 155786
rect 385500 155722 385552 155728
rect 384488 155508 384540 155514
rect 384488 155450 384540 155456
rect 384764 155508 384816 155514
rect 384764 155450 384816 155456
rect 384580 154828 384632 154834
rect 384580 154770 384632 154776
rect 383476 154624 383528 154630
rect 383476 154566 383528 154572
rect 384028 154488 384080 154494
rect 384028 154430 384080 154436
rect 382372 153944 382424 153950
rect 382372 153886 382424 153892
rect 383292 153944 383344 153950
rect 383292 153886 383344 153892
rect 382740 153808 382792 153814
rect 382740 153750 382792 153756
rect 382280 153468 382332 153474
rect 382280 153410 382332 153416
rect 382752 151994 382780 153750
rect 383304 151994 383332 153886
rect 384040 151994 384068 154430
rect 384592 153542 384620 154770
rect 384672 154420 384724 154426
rect 384672 154362 384724 154368
rect 384580 153536 384632 153542
rect 384580 153478 384632 153484
rect 384684 151994 384712 154362
rect 384776 153406 384804 155450
rect 384948 154284 385000 154290
rect 384948 154226 385000 154232
rect 384764 153400 384816 153406
rect 384764 153342 384816 153348
rect 377200 151966 377536 151994
rect 377844 151966 378088 151994
rect 378488 151966 378824 151994
rect 379132 151966 379468 151994
rect 379776 151966 380112 151994
rect 380420 151966 380756 151994
rect 381156 151966 381492 151994
rect 381800 151966 382136 151994
rect 382444 151966 382780 151994
rect 383088 151966 383332 151994
rect 383732 151966 384068 151994
rect 384376 151966 384712 151994
rect 384960 151994 384988 154226
rect 385512 153270 385540 155722
rect 386328 155576 386380 155582
rect 386328 155518 386380 155524
rect 385960 154352 386012 154358
rect 385960 154294 386012 154300
rect 385500 153264 385552 153270
rect 385500 153206 385552 153212
rect 385972 151994 386000 154294
rect 386236 154216 386288 154222
rect 386236 154158 386288 154164
rect 384960 151966 385020 151994
rect 385664 151966 386000 151994
rect 386248 151994 386276 154158
rect 386340 153610 386368 155518
rect 386432 155242 386460 159200
rect 387340 155848 387392 155854
rect 387340 155790 387392 155796
rect 386420 155236 386472 155242
rect 386420 155178 386472 155184
rect 387352 154154 387380 155790
rect 387444 154834 387472 159200
rect 388364 155514 388392 159200
rect 388444 155916 388496 155922
rect 388444 155858 388496 155864
rect 388352 155508 388404 155514
rect 388352 155450 388404 155456
rect 387432 154828 387484 154834
rect 387432 154770 387484 154776
rect 387340 154148 387392 154154
rect 387340 154090 387392 154096
rect 387708 154080 387760 154086
rect 387708 154022 387760 154028
rect 386328 153604 386380 153610
rect 386328 153546 386380 153552
rect 387248 153332 387300 153338
rect 387248 153274 387300 153280
rect 387260 151994 387288 153274
rect 387720 151994 387748 154022
rect 388456 153814 388484 155858
rect 389376 155582 389404 159200
rect 390296 155786 390324 159200
rect 391308 155854 391336 159200
rect 391296 155848 391348 155854
rect 391296 155790 391348 155796
rect 390284 155780 390336 155786
rect 390284 155722 390336 155728
rect 389364 155576 389416 155582
rect 389364 155518 389416 155524
rect 392320 154562 392348 159200
rect 393240 155922 393268 159200
rect 393228 155916 393280 155922
rect 393228 155858 393280 155864
rect 392308 154556 392360 154562
rect 392308 154498 392360 154504
rect 390468 154148 390520 154154
rect 390468 154090 390520 154096
rect 388536 154012 388588 154018
rect 388536 153954 388588 153960
rect 388444 153808 388496 153814
rect 388444 153750 388496 153756
rect 388548 151994 388576 153954
rect 389088 153672 389140 153678
rect 389088 153614 389140 153620
rect 389100 151994 389128 153614
rect 389824 153604 389876 153610
rect 389824 153546 389876 153552
rect 389836 151994 389864 153546
rect 390480 151994 390508 154090
rect 394252 153950 394280 159200
rect 395172 154494 395200 159200
rect 395988 154556 396040 154562
rect 395988 154498 396040 154504
rect 395160 154488 395212 154494
rect 395160 154430 395212 154436
rect 395712 154488 395764 154494
rect 395712 154430 395764 154436
rect 394240 153944 394292 153950
rect 394240 153886 394292 153892
rect 394424 153944 394476 153950
rect 394424 153886 394476 153892
rect 391204 153876 391256 153882
rect 391204 153818 391256 153824
rect 391216 151994 391244 153818
rect 393044 153740 393096 153746
rect 393044 153682 393096 153688
rect 392492 153468 392544 153474
rect 392492 153410 392544 153416
rect 391848 153400 391900 153406
rect 391848 153342 391900 153348
rect 391860 151994 391888 153342
rect 392504 151994 392532 153410
rect 393056 151994 393084 153682
rect 393780 153536 393832 153542
rect 393780 153478 393832 153484
rect 393792 151994 393820 153478
rect 394436 151994 394464 153886
rect 395068 153808 395120 153814
rect 395068 153750 395120 153756
rect 395080 151994 395108 153750
rect 395724 151994 395752 154430
rect 386248 151966 386308 151994
rect 386952 151966 387288 151994
rect 387596 151966 387748 151994
rect 388240 151966 388576 151994
rect 388884 151966 389128 151994
rect 389528 151966 389864 151994
rect 390264 151966 390508 151994
rect 390908 151966 391244 151994
rect 391552 151966 391888 151994
rect 392196 151966 392532 151994
rect 392840 151966 393084 151994
rect 393484 151966 393820 151994
rect 394128 151966 394464 151994
rect 394772 151966 395108 151994
rect 395416 151966 395752 151994
rect 396000 151994 396028 154498
rect 396184 154426 396212 159200
rect 396172 154420 396224 154426
rect 396172 154362 396224 154368
rect 397000 154420 397052 154426
rect 397000 154362 397052 154368
rect 397012 151994 397040 154362
rect 397196 154290 397224 159200
rect 398116 154358 398144 159200
rect 398564 155168 398616 155174
rect 398564 155110 398616 155116
rect 398104 154352 398156 154358
rect 398104 154294 398156 154300
rect 398288 154352 398340 154358
rect 398288 154294 398340 154300
rect 397184 154284 397236 154290
rect 397184 154226 397236 154232
rect 397276 154284 397328 154290
rect 397276 154226 397328 154232
rect 396000 151966 396060 151994
rect 396704 151966 397040 151994
rect 397288 151994 397316 154226
rect 398300 151994 398328 154294
rect 397288 151966 397348 151994
rect 397992 151966 398328 151994
rect 398576 151858 398604 155110
rect 398852 154578 398880 159310
rect 399036 159202 399064 159310
rect 399114 159202 399170 160000
rect 399036 159200 399170 159202
rect 400034 159200 400090 160000
rect 401046 159200 401102 160000
rect 402058 159200 402114 160000
rect 402978 159200 403034 160000
rect 403990 159200 404046 160000
rect 404910 159200 404966 160000
rect 405922 159200 405978 160000
rect 406934 159200 406990 160000
rect 407854 159200 407910 160000
rect 408866 159200 408922 160000
rect 409786 159200 409842 160000
rect 410798 159200 410854 160000
rect 411810 159200 411866 160000
rect 412730 159200 412786 160000
rect 413742 159200 413798 160000
rect 414662 159200 414718 160000
rect 415674 159200 415730 160000
rect 416686 159200 416742 160000
rect 417606 159200 417662 160000
rect 418618 159200 418674 160000
rect 419538 159200 419594 160000
rect 420550 159200 420606 160000
rect 421562 159200 421618 160000
rect 422482 159200 422538 160000
rect 423494 159200 423550 160000
rect 424414 159200 424470 160000
rect 425426 159200 425482 160000
rect 426346 159200 426402 160000
rect 427358 159200 427414 160000
rect 428370 159200 428426 160000
rect 429290 159200 429346 160000
rect 430302 159200 430358 160000
rect 431222 159200 431278 160000
rect 432234 159200 432290 160000
rect 433246 159200 433302 160000
rect 434166 159200 434222 160000
rect 435178 159200 435234 160000
rect 436098 159200 436154 160000
rect 437110 159200 437166 160000
rect 438122 159200 438178 160000
rect 439042 159200 439098 160000
rect 440054 159200 440110 160000
rect 440974 159200 441030 160000
rect 441986 159200 442042 160000
rect 442998 159200 443054 160000
rect 443918 159200 443974 160000
rect 444930 159200 444986 160000
rect 445850 159200 445906 160000
rect 446862 159200 446918 160000
rect 447874 159200 447930 160000
rect 448794 159200 448850 160000
rect 449806 159200 449862 160000
rect 450726 159200 450782 160000
rect 451738 159200 451794 160000
rect 452750 159200 452806 160000
rect 453670 159200 453726 160000
rect 454682 159200 454738 160000
rect 455602 159200 455658 160000
rect 456614 159200 456670 160000
rect 457626 159200 457682 160000
rect 458546 159200 458602 160000
rect 459558 159200 459614 160000
rect 460478 159200 460534 160000
rect 461490 159200 461546 160000
rect 462502 159200 462558 160000
rect 463422 159200 463478 160000
rect 464434 159200 464490 160000
rect 465354 159200 465410 160000
rect 466366 159200 466422 160000
rect 467286 159200 467342 160000
rect 468298 159200 468354 160000
rect 469310 159200 469366 160000
rect 470230 159200 470286 160000
rect 471242 159200 471298 160000
rect 472162 159200 472218 160000
rect 473174 159200 473230 160000
rect 474186 159200 474242 160000
rect 475106 159200 475162 160000
rect 476118 159200 476174 160000
rect 477038 159200 477094 160000
rect 478050 159200 478106 160000
rect 479062 159200 479118 160000
rect 479982 159200 480038 160000
rect 480994 159200 481050 160000
rect 481914 159200 481970 160000
rect 482926 159200 482982 160000
rect 483938 159200 483994 160000
rect 484858 159200 484914 160000
rect 485870 159200 485926 160000
rect 486790 159200 486846 160000
rect 487802 159200 487858 160000
rect 488814 159200 488870 160000
rect 489288 159310 489684 159338
rect 399036 159174 399156 159200
rect 398932 155100 398984 155106
rect 398932 155042 398984 155048
rect 398760 154550 398880 154578
rect 398760 154222 398788 154550
rect 398748 154216 398800 154222
rect 398748 154158 398800 154164
rect 398944 154086 398972 155042
rect 399484 154760 399536 154766
rect 399484 154702 399536 154708
rect 398932 154080 398984 154086
rect 398932 154022 398984 154028
rect 399496 151994 399524 154702
rect 400048 153338 400076 159200
rect 401060 155106 401088 159200
rect 401600 155372 401652 155378
rect 401600 155314 401652 155320
rect 401508 155236 401560 155242
rect 401508 155178 401560 155184
rect 401048 155100 401100 155106
rect 401048 155042 401100 155048
rect 400956 155032 401008 155038
rect 400956 154974 401008 154980
rect 400312 154964 400364 154970
rect 400312 154906 400364 154912
rect 400220 154828 400272 154834
rect 400220 154770 400272 154776
rect 400128 154216 400180 154222
rect 400128 154158 400180 154164
rect 400036 153332 400088 153338
rect 400036 153274 400088 153280
rect 400140 151994 400168 154158
rect 400232 154018 400260 154770
rect 400220 154012 400272 154018
rect 400220 153954 400272 153960
rect 400324 153678 400352 154906
rect 400312 153672 400364 153678
rect 400312 153614 400364 153620
rect 400968 151994 400996 154974
rect 401520 151994 401548 155178
rect 401612 154154 401640 155314
rect 401692 155032 401744 155038
rect 401692 154974 401744 154980
rect 401600 154148 401652 154154
rect 401600 154090 401652 154096
rect 401704 153610 401732 154974
rect 402072 154834 402100 159200
rect 402244 155848 402296 155854
rect 402244 155790 402296 155796
rect 402060 154828 402112 154834
rect 402060 154770 402112 154776
rect 401692 153604 401744 153610
rect 401692 153546 401744 153552
rect 402256 151994 402284 155790
rect 402992 154970 403020 159200
rect 404004 155038 404032 159200
rect 404176 155916 404228 155922
rect 404176 155858 404228 155864
rect 404084 155644 404136 155650
rect 404084 155586 404136 155592
rect 403992 155032 404044 155038
rect 403992 154974 404044 154980
rect 402980 154964 403032 154970
rect 402980 154906 403032 154912
rect 403992 154624 404044 154630
rect 403992 154566 404044 154572
rect 403532 154148 403584 154154
rect 403532 154090 403584 154096
rect 402704 154080 402756 154086
rect 402704 154022 402756 154028
rect 402716 151994 402744 154022
rect 403544 151994 403572 154090
rect 404004 153882 404032 154566
rect 403992 153876 404044 153882
rect 403992 153818 404044 153824
rect 404096 151994 404124 155586
rect 404188 153406 404216 155858
rect 404820 155712 404872 155718
rect 404820 155654 404872 155660
rect 404636 155508 404688 155514
rect 404636 155450 404688 155456
rect 404648 153474 404676 155450
rect 404636 153468 404688 153474
rect 404636 153410 404688 153416
rect 404176 153400 404228 153406
rect 404176 153342 404228 153348
rect 404832 151994 404860 155654
rect 404924 155378 404952 159200
rect 405832 155780 405884 155786
rect 405832 155722 405884 155728
rect 404912 155372 404964 155378
rect 404912 155314 404964 155320
rect 405464 154012 405516 154018
rect 405464 153954 405516 153960
rect 405476 151994 405504 153954
rect 405844 153542 405872 155722
rect 405936 154630 405964 159200
rect 406948 155922 406976 159200
rect 406936 155916 406988 155922
rect 406936 155858 406988 155864
rect 406752 155576 406804 155582
rect 406752 155518 406804 155524
rect 406108 154692 406160 154698
rect 406108 154634 406160 154640
rect 405924 154624 405976 154630
rect 405924 154566 405976 154572
rect 405832 153536 405884 153542
rect 405832 153478 405884 153484
rect 406120 151994 406148 154634
rect 406764 151994 406792 155518
rect 407868 155514 407896 159200
rect 407856 155508 407908 155514
rect 407856 155450 407908 155456
rect 408316 155508 408368 155514
rect 408316 155450 408368 155456
rect 407028 154760 407080 154766
rect 407028 154702 407080 154708
rect 399280 151966 399524 151994
rect 400016 151966 400168 151994
rect 400660 151966 400996 151994
rect 401304 151966 401548 151994
rect 401948 151966 402284 151994
rect 402592 151966 402744 151994
rect 403236 151966 403572 151994
rect 403880 151966 404124 151994
rect 404524 151966 404860 151994
rect 405168 151966 405504 151994
rect 405812 151966 406148 151994
rect 406456 151966 406792 151994
rect 407040 151994 407068 154702
rect 408040 153876 408092 153882
rect 408040 153818 408092 153824
rect 408052 151994 408080 153818
rect 407040 151966 407100 151994
rect 407744 151966 408080 151994
rect 408328 151858 408356 155450
rect 408880 153746 408908 159200
rect 409800 155786 409828 159200
rect 409788 155780 409840 155786
rect 409788 155722 409840 155728
rect 409696 155440 409748 155446
rect 409696 155382 409748 155388
rect 409420 154624 409472 154630
rect 409420 154566 409472 154572
rect 408868 153740 408920 153746
rect 408868 153682 408920 153688
rect 409432 151994 409460 154566
rect 409124 151966 409460 151994
rect 409708 151858 409736 155382
rect 410812 153950 410840 159200
rect 411352 155780 411404 155786
rect 411352 155722 411404 155728
rect 411260 155712 411312 155718
rect 411260 155654 411312 155660
rect 411168 155372 411220 155378
rect 411168 155314 411220 155320
rect 410800 153944 410852 153950
rect 410800 153886 410852 153892
rect 410708 153604 410760 153610
rect 410708 153546 410760 153552
rect 410720 151994 410748 153546
rect 411180 151994 411208 155314
rect 411272 154562 411300 155654
rect 411260 154556 411312 154562
rect 411260 154498 411312 154504
rect 411364 154494 411392 155722
rect 411352 154488 411404 154494
rect 411352 154430 411404 154436
rect 411824 153814 411852 159200
rect 412744 155786 412772 159200
rect 412732 155780 412784 155786
rect 412732 155722 412784 155728
rect 413284 155780 413336 155786
rect 413284 155722 413336 155728
rect 411996 154692 412048 154698
rect 411996 154634 412048 154640
rect 411812 153808 411864 153814
rect 411812 153750 411864 153756
rect 412008 151994 412036 154634
rect 413296 154426 413324 155722
rect 413756 155718 413784 159200
rect 414676 155786 414704 159200
rect 414664 155780 414716 155786
rect 414664 155722 414716 155728
rect 413744 155712 413796 155718
rect 413744 155654 413796 155660
rect 414112 155712 414164 155718
rect 414112 155654 414164 155660
rect 413836 154828 413888 154834
rect 413836 154770 413888 154776
rect 413284 154420 413336 154426
rect 413284 154362 413336 154368
rect 413284 153740 413336 153746
rect 413284 153682 413336 153688
rect 412456 153264 412508 153270
rect 412456 153206 412508 153212
rect 412468 151994 412496 153206
rect 413296 151994 413324 153682
rect 413848 153270 413876 154770
rect 414124 154358 414152 155654
rect 414572 155304 414624 155310
rect 414572 155246 414624 155252
rect 414112 154352 414164 154358
rect 414112 154294 414164 154300
rect 413928 153672 413980 153678
rect 413928 153614 413980 153620
rect 413836 153264 413888 153270
rect 413836 153206 413888 153212
rect 413940 151994 413968 153614
rect 414584 151994 414612 155246
rect 415216 154760 415268 154766
rect 415216 154702 415268 154708
rect 415228 151994 415256 154702
rect 415688 154290 415716 159200
rect 416700 155718 416728 159200
rect 416688 155712 416740 155718
rect 416688 155654 416740 155660
rect 417620 155174 417648 159200
rect 417608 155168 417660 155174
rect 417608 155110 417660 155116
rect 418632 155038 418660 159200
rect 419448 155168 419500 155174
rect 419448 155110 419500 155116
rect 418620 155032 418672 155038
rect 418620 154974 418672 154980
rect 417792 154964 417844 154970
rect 417792 154906 417844 154912
rect 415860 154556 415912 154562
rect 415860 154498 415912 154504
rect 415676 154284 415728 154290
rect 415676 154226 415728 154232
rect 415872 151994 415900 154498
rect 416504 154488 416556 154494
rect 416504 154430 416556 154436
rect 416516 151994 416544 154430
rect 417148 153332 417200 153338
rect 417148 153274 417200 153280
rect 417160 151994 417188 153274
rect 417804 151994 417832 154906
rect 417976 154828 418028 154834
rect 417976 154770 418028 154776
rect 417988 153338 418016 154770
rect 419172 154420 419224 154426
rect 419172 154362 419224 154368
rect 418528 153808 418580 153814
rect 418528 153750 418580 153756
rect 417976 153332 418028 153338
rect 417976 153274 418028 153280
rect 418540 151994 418568 153750
rect 419184 151994 419212 154362
rect 410412 151966 410748 151994
rect 411056 151966 411208 151994
rect 411700 151966 412036 151994
rect 412344 151966 412496 151994
rect 412988 151966 413324 151994
rect 413632 151966 413968 151994
rect 414276 151966 414612 151994
rect 414920 151966 415256 151994
rect 415564 151966 415900 151994
rect 416208 151966 416544 151994
rect 416852 151966 417188 151994
rect 417496 151966 417832 151994
rect 418232 151966 418568 151994
rect 418876 151966 419212 151994
rect 419460 151994 419488 155110
rect 419552 154222 419580 159200
rect 420564 155106 420592 159200
rect 420736 156664 420788 156670
rect 420736 156606 420788 156612
rect 420552 155100 420604 155106
rect 420552 155042 420604 155048
rect 420460 155032 420512 155038
rect 420460 154974 420512 154980
rect 419540 154216 419592 154222
rect 419540 154158 419592 154164
rect 420472 151994 420500 154974
rect 419460 151966 419520 151994
rect 420164 151966 420500 151994
rect 420748 151858 420776 156606
rect 421576 155242 421604 159200
rect 422496 155854 422524 159200
rect 422484 155848 422536 155854
rect 422484 155790 422536 155796
rect 421564 155236 421616 155242
rect 421564 155178 421616 155184
rect 422208 155236 422260 155242
rect 422208 155178 422260 155184
rect 421748 154352 421800 154358
rect 421748 154294 421800 154300
rect 421760 151994 421788 154294
rect 421452 151966 421788 151994
rect 422220 151858 422248 155178
rect 423036 155100 423088 155106
rect 423036 155042 423088 155048
rect 423048 151994 423076 155042
rect 423508 154086 423536 159200
rect 424324 154284 424376 154290
rect 424324 154226 424376 154232
rect 423496 154080 423548 154086
rect 423496 154022 423548 154028
rect 423588 152516 423640 152522
rect 423588 152458 423640 152464
rect 423600 151994 423628 152458
rect 424336 151994 424364 154226
rect 424428 154154 424456 159200
rect 424968 155848 425020 155854
rect 424968 155790 425020 155796
rect 424416 154148 424468 154154
rect 424416 154090 424468 154096
rect 424980 151994 425008 155790
rect 425440 155650 425468 159200
rect 426256 157344 426308 157350
rect 426256 157286 426308 157292
rect 425612 155848 425664 155854
rect 425612 155790 425664 155796
rect 425428 155644 425480 155650
rect 425428 155586 425480 155592
rect 425624 151994 425652 155790
rect 426268 151994 426296 157286
rect 426360 155922 426388 159200
rect 426348 155916 426400 155922
rect 426348 155858 426400 155864
rect 426900 154216 426952 154222
rect 426900 154158 426952 154164
rect 426912 151994 426940 154158
rect 427372 154018 427400 159200
rect 428280 155848 428332 155854
rect 428280 155790 428332 155796
rect 427636 155644 427688 155650
rect 427636 155586 427688 155592
rect 427360 154012 427412 154018
rect 427360 153954 427412 153960
rect 427648 151994 427676 155586
rect 428292 151994 428320 155790
rect 428384 155786 428412 159200
rect 428924 157276 428976 157282
rect 428924 157218 428976 157224
rect 428372 155780 428424 155786
rect 428372 155722 428424 155728
rect 428936 151994 428964 157218
rect 429304 155582 429332 159200
rect 430316 155718 430344 159200
rect 430304 155712 430356 155718
rect 430304 155654 430356 155660
rect 430396 155712 430448 155718
rect 430396 155654 430448 155660
rect 429292 155576 429344 155582
rect 429292 155518 429344 155524
rect 429568 154148 429620 154154
rect 429568 154090 429620 154096
rect 429580 151994 429608 154090
rect 430408 151994 430436 155654
rect 430488 155576 430540 155582
rect 430488 155518 430540 155524
rect 422740 151966 423076 151994
rect 423384 151966 423628 151994
rect 424028 151966 424364 151994
rect 424672 151966 425008 151994
rect 425316 151966 425652 151994
rect 425960 151966 426296 151994
rect 426604 151966 426940 151994
rect 427340 151966 427676 151994
rect 427984 151966 428320 151994
rect 428628 151966 428964 151994
rect 429272 151966 429608 151994
rect 429916 151966 430436 151994
rect 430500 151994 430528 155518
rect 431236 153882 431264 159200
rect 432248 155514 432276 159200
rect 432236 155508 432288 155514
rect 432236 155450 432288 155456
rect 433064 155508 433116 155514
rect 433064 155450 433116 155456
rect 431776 154080 431828 154086
rect 431776 154022 431828 154028
rect 431224 153876 431276 153882
rect 431224 153818 431276 153824
rect 431500 153128 431552 153134
rect 431500 153070 431552 153076
rect 431512 151994 431540 153070
rect 430500 151966 430560 151994
rect 431204 151966 431540 151994
rect 431788 151994 431816 154022
rect 432788 154012 432840 154018
rect 432788 153954 432840 153960
rect 432800 151994 432828 153954
rect 431788 151966 431848 151994
rect 432492 151966 432828 151994
rect 247000 151852 247112 151858
rect 246948 151846 247112 151852
rect 246960 151830 247112 151846
rect 252020 151842 252356 151858
rect 252008 151836 252356 151842
rect 211068 151778 211120 151784
rect 252060 151830 252356 151836
rect 364168 151830 364228 151858
rect 375208 151830 375268 151858
rect 376496 151830 376556 151858
rect 398576 151830 398636 151858
rect 408328 151830 408388 151858
rect 409708 151830 409768 151858
rect 420748 151830 420808 151858
rect 422096 151830 422248 151858
rect 433076 151858 433104 155450
rect 433260 154630 433288 159200
rect 434180 155446 434208 159200
rect 434168 155440 434220 155446
rect 434168 155382 434220 155388
rect 433248 154624 433300 154630
rect 433248 154566 433300 154572
rect 434628 153876 434680 153882
rect 434628 153818 434680 153824
rect 434076 153060 434128 153066
rect 434076 153002 434128 153008
rect 434088 151994 434116 153002
rect 434640 151994 434668 153818
rect 435192 153610 435220 159200
rect 436008 155440 436060 155446
rect 436008 155382 436060 155388
rect 435364 153944 435416 153950
rect 435364 153886 435416 153892
rect 435180 153604 435232 153610
rect 435180 153546 435232 153552
rect 435376 151994 435404 153886
rect 436020 151994 436048 155382
rect 436112 155378 436140 159200
rect 436652 157208 436704 157214
rect 436652 157150 436704 157156
rect 436100 155372 436152 155378
rect 436100 155314 436152 155320
rect 436664 151994 436692 157150
rect 437124 154698 437152 159200
rect 438032 157140 438084 157146
rect 438032 157082 438084 157088
rect 437388 157072 437440 157078
rect 437388 157014 437440 157020
rect 437112 154692 437164 154698
rect 437112 154634 437164 154640
rect 437400 151994 437428 157014
rect 438044 151994 438072 157082
rect 438136 154766 438164 159200
rect 438676 155372 438728 155378
rect 438676 155314 438728 155320
rect 438124 154760 438176 154766
rect 438124 154702 438176 154708
rect 438688 151994 438716 155314
rect 439056 153746 439084 159200
rect 439044 153740 439096 153746
rect 439044 153682 439096 153688
rect 440068 153678 440096 159200
rect 440608 156460 440660 156466
rect 440608 156402 440660 156408
rect 440056 153672 440108 153678
rect 440056 153614 440108 153620
rect 439964 152992 440016 152998
rect 439964 152934 440016 152940
rect 439320 152448 439372 152454
rect 439320 152390 439372 152396
rect 439332 151994 439360 152390
rect 439976 151994 440004 152934
rect 440620 151994 440648 156402
rect 440988 155310 441016 159200
rect 440976 155304 441028 155310
rect 440976 155246 441028 155252
rect 441252 155304 441304 155310
rect 441252 155246 441304 155252
rect 441264 151994 441292 155246
rect 442000 154902 442028 159200
rect 442540 157004 442592 157010
rect 442540 156946 442592 156952
rect 441988 154896 442040 154902
rect 441988 154838 442040 154844
rect 441712 152924 441764 152930
rect 441712 152866 441764 152872
rect 433780 151966 434116 151994
rect 434424 151966 434668 151994
rect 435068 151966 435404 151994
rect 435712 151966 436048 151994
rect 436356 151966 436692 151994
rect 437092 151966 437428 151994
rect 437736 151966 438072 151994
rect 438380 151966 438716 151994
rect 439024 151966 439360 151994
rect 439668 151966 440004 151994
rect 440312 151966 440648 151994
rect 440956 151966 441292 151994
rect 441724 151858 441752 152866
rect 442552 151994 442580 156946
rect 442816 156936 442868 156942
rect 442816 156878 442868 156884
rect 442244 151966 442580 151994
rect 433076 151830 433136 151858
rect 441600 151830 441752 151858
rect 442828 151858 442856 156878
rect 443012 154562 443040 159200
rect 443000 154556 443052 154562
rect 443000 154498 443052 154504
rect 443932 154494 443960 159200
rect 444944 154834 444972 159200
rect 445116 156868 445168 156874
rect 445116 156810 445168 156816
rect 444932 154828 444984 154834
rect 444932 154770 444984 154776
rect 443920 154488 443972 154494
rect 443920 154430 443972 154436
rect 444288 152856 444340 152862
rect 444288 152798 444340 152804
rect 443828 152040 443880 152046
rect 443532 151988 443828 151994
rect 444300 151994 444328 152798
rect 445128 151994 445156 156810
rect 445668 156800 445720 156806
rect 445668 156742 445720 156748
rect 445680 151994 445708 156742
rect 445864 154970 445892 159200
rect 446496 156052 446548 156058
rect 446496 155994 446548 156000
rect 445852 154964 445904 154970
rect 445852 154906 445904 154912
rect 446508 151994 446536 155994
rect 446876 153814 446904 159200
rect 447784 155984 447836 155990
rect 447784 155926 447836 155932
rect 446864 153808 446916 153814
rect 446864 153750 446916 153756
rect 447048 152788 447100 152794
rect 447048 152730 447100 152736
rect 447060 151994 447088 152730
rect 447796 151994 447824 155926
rect 447888 154426 447916 159200
rect 448808 155174 448836 159200
rect 449072 156732 449124 156738
rect 449072 156674 449124 156680
rect 448796 155168 448848 155174
rect 448796 155110 448848 155116
rect 447876 154420 447928 154426
rect 447876 154362 447928 154368
rect 448428 152720 448480 152726
rect 448428 152662 448480 152668
rect 448440 151994 448468 152662
rect 449084 151994 449112 156674
rect 449820 155038 449848 159200
rect 450740 156670 450768 159200
rect 450728 156664 450780 156670
rect 450728 156606 450780 156612
rect 450360 156120 450412 156126
rect 450360 156062 450412 156068
rect 449808 155032 449860 155038
rect 449808 154974 449860 154980
rect 449394 152108 449446 152114
rect 449394 152050 449446 152056
rect 443532 151982 443880 151988
rect 443532 151966 443868 151982
rect 444176 151966 444328 151994
rect 444820 151966 445156 151994
rect 445464 151966 445708 151994
rect 446200 151966 446536 151994
rect 446844 151966 447088 151994
rect 447488 151966 447824 151994
rect 448132 151966 448468 151994
rect 448776 151966 449112 151994
rect 449406 151980 449434 152050
rect 450372 151994 450400 156062
rect 451752 154358 451780 159200
rect 452292 156188 452344 156194
rect 452292 156130 452344 156136
rect 451740 154352 451792 154358
rect 451740 154294 451792 154300
rect 451648 152652 451700 152658
rect 451648 152594 451700 152600
rect 450912 152584 450964 152590
rect 450912 152526 450964 152532
rect 450924 151994 450952 152526
rect 451660 151994 451688 152594
rect 452304 151994 452332 156130
rect 452764 155242 452792 159200
rect 453580 156256 453632 156262
rect 453580 156198 453632 156204
rect 452752 155236 452804 155242
rect 452752 155178 452804 155184
rect 452614 152176 452666 152182
rect 452614 152118 452666 152124
rect 450064 151966 450400 151994
rect 450708 151966 450952 151994
rect 451352 151966 451688 151994
rect 451996 151966 452332 151994
rect 452626 151980 452654 152118
rect 453592 151994 453620 156198
rect 453684 155106 453712 159200
rect 453672 155100 453724 155106
rect 453672 155042 453724 155048
rect 454696 152522 454724 159200
rect 454868 155236 454920 155242
rect 454868 155178 454920 155184
rect 454684 152516 454736 152522
rect 454684 152458 454736 152464
rect 453902 152244 453954 152250
rect 453902 152186 453954 152192
rect 453284 151966 453620 151994
rect 453914 151980 453942 152186
rect 454880 151994 454908 155178
rect 455616 154290 455644 159200
rect 456628 155854 456656 159200
rect 456708 156664 456760 156670
rect 456708 156606 456760 156612
rect 456616 155848 456668 155854
rect 456616 155790 456668 155796
rect 455604 154284 455656 154290
rect 455604 154226 455656 154232
rect 455236 153468 455288 153474
rect 455236 153410 455288 153416
rect 454572 151966 454908 151994
rect 455248 151994 455276 153410
rect 456248 153400 456300 153406
rect 456248 153342 456300 153348
rect 456260 151994 456288 153342
rect 456720 151994 456748 156606
rect 457640 155922 457668 159200
rect 458560 157350 458588 159200
rect 458548 157344 458600 157350
rect 458548 157286 458600 157292
rect 457628 155916 457680 155922
rect 457628 155858 457680 155864
rect 459468 154828 459520 154834
rect 459468 154770 459520 154776
rect 457536 154624 457588 154630
rect 457536 154566 457588 154572
rect 457548 151994 457576 154566
rect 458088 153604 458140 153610
rect 458088 153546 458140 153552
rect 458100 151994 458128 153546
rect 458824 152516 458876 152522
rect 458824 152458 458876 152464
rect 458836 151994 458864 152458
rect 459480 151994 459508 154770
rect 459572 154222 459600 159200
rect 460492 155650 460520 159200
rect 460664 156324 460716 156330
rect 460664 156266 460716 156272
rect 460480 155644 460532 155650
rect 460480 155586 460532 155592
rect 460112 154760 460164 154766
rect 460112 154702 460164 154708
rect 459560 154216 459612 154222
rect 459560 154158 459612 154164
rect 460124 151994 460152 154702
rect 460676 151994 460704 156266
rect 461504 155786 461532 159200
rect 462516 157282 462544 159200
rect 462504 157276 462556 157282
rect 462504 157218 462556 157224
rect 461492 155780 461544 155786
rect 461492 155722 461544 155728
rect 462044 155032 462096 155038
rect 462044 154974 462096 154980
rect 461400 154692 461452 154698
rect 461400 154634 461452 154640
rect 461412 151994 461440 154634
rect 462056 151994 462084 154974
rect 463332 154896 463384 154902
rect 463332 154838 463384 154844
rect 462688 152312 462740 152318
rect 462688 152254 462740 152260
rect 462700 151994 462728 152254
rect 463344 151994 463372 154838
rect 463436 154154 463464 159200
rect 464448 155718 464476 159200
rect 464436 155712 464488 155718
rect 464436 155654 464488 155660
rect 465368 155582 465396 159200
rect 466000 156528 466052 156534
rect 466000 156470 466052 156476
rect 465356 155576 465408 155582
rect 465356 155518 465408 155524
rect 463608 155100 463660 155106
rect 463608 155042 463660 155048
rect 463424 154148 463476 154154
rect 463424 154090 463476 154096
rect 455248 151966 455308 151994
rect 455952 151966 456288 151994
rect 456596 151966 456748 151994
rect 457240 151966 457576 151994
rect 457884 151966 458128 151994
rect 458528 151966 458864 151994
rect 459172 151966 459508 151994
rect 459816 151966 460152 151994
rect 460460 151966 460704 151994
rect 461104 151966 461440 151994
rect 461748 151966 462084 151994
rect 462392 151966 462728 151994
rect 463036 151966 463372 151994
rect 463620 151994 463648 155042
rect 464620 154964 464672 154970
rect 464620 154906 464672 154912
rect 464632 151994 464660 154906
rect 464988 153672 465040 153678
rect 464988 153614 465040 153620
rect 463620 151966 463680 151994
rect 464324 151966 464660 151994
rect 465000 151994 465028 153614
rect 466012 151994 466040 156470
rect 466276 155916 466328 155922
rect 466276 155858 466328 155864
rect 465000 151966 465060 151994
rect 465704 151966 466040 151994
rect 466288 151994 466316 155858
rect 466380 153134 466408 159200
rect 467196 155168 467248 155174
rect 467196 155110 467248 155116
rect 466368 153128 466420 153134
rect 466368 153070 466420 153076
rect 467208 151994 467236 155110
rect 467300 154086 467328 159200
rect 467288 154080 467340 154086
rect 467288 154022 467340 154028
rect 468312 154018 468340 159200
rect 469128 155848 469180 155854
rect 469128 155790 469180 155796
rect 468300 154012 468352 154018
rect 468300 153954 468352 153960
rect 467748 153740 467800 153746
rect 467748 153682 467800 153688
rect 467760 151994 467788 153682
rect 468576 153196 468628 153202
rect 468576 153138 468628 153144
rect 468588 151994 468616 153138
rect 469140 151994 469168 155790
rect 469324 155514 469352 159200
rect 469864 156596 469916 156602
rect 469864 156538 469916 156544
rect 469312 155508 469364 155514
rect 469312 155450 469364 155456
rect 469876 151994 469904 156538
rect 470244 153066 470272 159200
rect 471152 155780 471204 155786
rect 471152 155722 471204 155728
rect 470324 153808 470376 153814
rect 470324 153750 470376 153756
rect 470232 153060 470284 153066
rect 470232 153002 470284 153008
rect 470336 151994 470364 153750
rect 471164 151994 471192 155722
rect 471256 153882 471284 159200
rect 471796 154556 471848 154562
rect 471796 154498 471848 154504
rect 471244 153876 471296 153882
rect 471244 153818 471296 153824
rect 471808 151994 471836 154498
rect 472176 153950 472204 159200
rect 473188 155446 473216 159200
rect 473728 157276 473780 157282
rect 473728 157218 473780 157224
rect 473176 155440 473228 155446
rect 473176 155382 473228 155388
rect 472164 153944 472216 153950
rect 472164 153886 472216 153892
rect 473084 153264 473136 153270
rect 473084 153206 473136 153212
rect 472440 153128 472492 153134
rect 472440 153070 472492 153076
rect 472452 151994 472480 153070
rect 473096 151994 473124 153206
rect 473740 151994 473768 157218
rect 474200 157214 474228 159200
rect 475016 157344 475068 157350
rect 475016 157286 475068 157292
rect 474188 157208 474240 157214
rect 474188 157150 474240 157156
rect 474464 154148 474516 154154
rect 474464 154090 474516 154096
rect 474476 151994 474504 154090
rect 475028 151994 475056 157286
rect 475120 157078 475148 159200
rect 476132 157146 476160 159200
rect 476120 157140 476172 157146
rect 476120 157082 476172 157088
rect 475108 157072 475160 157078
rect 475108 157014 475160 157020
rect 475752 155712 475804 155718
rect 475752 155654 475804 155660
rect 475764 151994 475792 155654
rect 477052 155378 477080 159200
rect 477316 157276 477368 157282
rect 477316 157218 477368 157224
rect 477040 155372 477092 155378
rect 477040 155314 477092 155320
rect 477040 153536 477092 153542
rect 477040 153478 477092 153484
rect 476120 153264 476172 153270
rect 476120 153206 476172 153212
rect 476028 153060 476080 153066
rect 476028 153002 476080 153008
rect 466288 151966 466348 151994
rect 466992 151966 467236 151994
rect 467636 151966 467788 151994
rect 468280 151966 468616 151994
rect 468924 151966 469168 151994
rect 469568 151966 469904 151994
rect 470212 151966 470364 151994
rect 470856 151966 471192 151994
rect 471500 151966 471836 151994
rect 472144 151966 472480 151994
rect 472788 151966 473124 151994
rect 473432 151966 473768 151994
rect 474168 151966 474504 151994
rect 474812 151966 475056 151994
rect 475456 151966 475792 151994
rect 476040 151994 476068 153002
rect 476132 152386 476160 153206
rect 476120 152380 476172 152386
rect 476120 152322 476172 152328
rect 477052 151994 477080 153478
rect 476040 151966 476100 151994
rect 476744 151966 477080 151994
rect 477328 151858 477356 157218
rect 478064 152454 478092 159200
rect 478788 157140 478840 157146
rect 478788 157082 478840 157088
rect 478328 155644 478380 155650
rect 478328 155586 478380 155592
rect 478052 152448 478104 152454
rect 478052 152390 478104 152396
rect 478340 151994 478368 155586
rect 478800 151994 478828 157082
rect 479076 152998 479104 159200
rect 479996 156466 480024 159200
rect 479984 156460 480036 156466
rect 479984 156402 480036 156408
rect 480076 156460 480128 156466
rect 480076 156402 480128 156408
rect 480088 154154 480116 156402
rect 480904 155576 480956 155582
rect 480904 155518 480956 155524
rect 480076 154148 480128 154154
rect 480076 154090 480128 154096
rect 479616 153876 479668 153882
rect 479616 153818 479668 153824
rect 479064 152992 479116 152998
rect 479064 152934 479116 152940
rect 479628 151994 479656 153818
rect 480076 152992 480128 152998
rect 480076 152934 480128 152940
rect 480088 151994 480116 152934
rect 480916 151994 480944 155518
rect 481008 155310 481036 159200
rect 481548 156392 481600 156398
rect 481548 156334 481600 156340
rect 480996 155304 481048 155310
rect 480996 155246 481048 155252
rect 481560 151994 481588 156334
rect 481928 152930 481956 159200
rect 482940 157010 482968 159200
rect 482928 157004 482980 157010
rect 482928 156946 482980 156952
rect 483020 157004 483072 157010
rect 483020 156946 483072 156952
rect 483032 156890 483060 156946
rect 483952 156942 483980 159200
rect 482940 156862 483060 156890
rect 483940 156936 483992 156942
rect 483940 156878 483992 156884
rect 482192 154420 482244 154426
rect 482192 154362 482244 154368
rect 481916 152924 481968 152930
rect 481916 152866 481968 152872
rect 482204 151994 482232 154362
rect 482744 153536 482796 153542
rect 482744 153478 482796 153484
rect 482756 152454 482784 153478
rect 482744 152448 482796 152454
rect 482744 152390 482796 152396
rect 482940 151994 482968 156862
rect 484872 155666 484900 159200
rect 485504 156936 485556 156942
rect 485504 156878 485556 156884
rect 484872 155638 484992 155666
rect 484860 155508 484912 155514
rect 484860 155450 484912 155456
rect 483572 155440 483624 155446
rect 483572 155382 483624 155388
rect 483584 151994 483612 155382
rect 484216 152924 484268 152930
rect 484216 152866 484268 152872
rect 484228 151994 484256 152866
rect 484872 151994 484900 155450
rect 484964 152046 484992 155638
rect 478032 151966 478368 151994
rect 478676 151966 478828 151994
rect 479320 151966 479656 151994
rect 479964 151966 480116 151994
rect 480608 151966 480944 151994
rect 481252 151966 481588 151994
rect 481896 151966 482232 151994
rect 482540 151966 482968 151994
rect 483276 151966 483612 151994
rect 483920 151966 484256 151994
rect 484564 151966 484900 151994
rect 484952 152040 485004 152046
rect 485516 151994 485544 156878
rect 485884 152862 485912 159200
rect 486804 156874 486832 159200
rect 486792 156868 486844 156874
rect 486792 156810 486844 156816
rect 486884 156868 486936 156874
rect 486884 156810 486936 156816
rect 486148 154352 486200 154358
rect 486148 154294 486200 154300
rect 485872 152856 485924 152862
rect 485872 152798 485924 152804
rect 486160 151994 486188 154294
rect 486896 151994 486924 156810
rect 487816 156806 487844 159200
rect 487804 156800 487856 156806
rect 487804 156742 487856 156748
rect 487160 156392 487212 156398
rect 487160 156334 487212 156340
rect 487068 154284 487120 154290
rect 487068 154226 487120 154232
rect 484952 151982 485004 151988
rect 485208 151966 485544 151994
rect 485852 151966 486188 151994
rect 486496 151966 486924 151994
rect 487080 151994 487108 154226
rect 487172 153882 487200 156334
rect 488828 156058 488856 159200
rect 488816 156052 488868 156058
rect 488816 155994 488868 156000
rect 488356 155304 488408 155310
rect 488356 155246 488408 155252
rect 487160 153876 487212 153882
rect 487160 153818 487212 153824
rect 488080 152856 488132 152862
rect 488080 152798 488132 152804
rect 488092 151994 488120 152798
rect 487080 151966 487140 151994
rect 487784 151966 488120 151994
rect 488368 151994 488396 155246
rect 489288 152794 489316 159310
rect 489656 159202 489684 159310
rect 489734 159202 489790 160000
rect 489656 159200 489790 159202
rect 490746 159200 490802 160000
rect 491666 159200 491722 160000
rect 492678 159200 492734 160000
rect 493690 159200 493746 160000
rect 494610 159200 494666 160000
rect 495622 159200 495678 160000
rect 496542 159200 496598 160000
rect 497554 159200 497610 160000
rect 498566 159200 498622 160000
rect 499486 159200 499542 160000
rect 500498 159200 500554 160000
rect 501418 159200 501474 160000
rect 502430 159200 502486 160000
rect 503350 159200 503406 160000
rect 504362 159200 504418 160000
rect 505374 159200 505430 160000
rect 506294 159200 506350 160000
rect 507306 159200 507362 160000
rect 508226 159200 508282 160000
rect 509238 159200 509294 160000
rect 510250 159200 510306 160000
rect 511170 159200 511226 160000
rect 512182 159200 512238 160000
rect 513102 159200 513158 160000
rect 514114 159200 514170 160000
rect 515126 159200 515182 160000
rect 516046 159200 516102 160000
rect 517058 159200 517114 160000
rect 517978 159200 518034 160000
rect 518990 159200 519046 160000
rect 520002 159200 520058 160000
rect 520922 159200 520978 160000
rect 521934 159200 521990 160000
rect 522854 159200 522910 160000
rect 523866 159200 523922 160000
rect 524878 159200 524934 160000
rect 525798 159200 525854 160000
rect 526810 159200 526866 160000
rect 527730 159200 527786 160000
rect 528742 159200 528798 160000
rect 529754 159200 529810 160000
rect 530674 159200 530730 160000
rect 531686 159200 531742 160000
rect 532606 159200 532662 160000
rect 533618 159200 533674 160000
rect 534630 159200 534686 160000
rect 535550 159200 535606 160000
rect 536562 159200 536618 160000
rect 537482 159200 537538 160000
rect 538494 159200 538550 160000
rect 539506 159200 539562 160000
rect 540426 159200 540482 160000
rect 541438 159200 541494 160000
rect 542358 159200 542414 160000
rect 543370 159200 543426 160000
rect 544290 159200 544346 160000
rect 545302 159200 545358 160000
rect 546314 159200 546370 160000
rect 547234 159200 547290 160000
rect 548246 159200 548302 160000
rect 549166 159200 549222 160000
rect 550178 159200 550234 160000
rect 551190 159200 551246 160000
rect 552110 159200 552166 160000
rect 553122 159200 553178 160000
rect 554042 159200 554098 160000
rect 555054 159200 555110 160000
rect 556066 159200 556122 160000
rect 556986 159200 557042 160000
rect 557998 159200 558054 160000
rect 558918 159200 558974 160000
rect 559930 159200 559986 160000
rect 560942 159200 560998 160000
rect 561862 159200 561918 160000
rect 562874 159200 562930 160000
rect 563794 159200 563850 160000
rect 564806 159200 564862 160000
rect 565818 159200 565874 160000
rect 566738 159200 566794 160000
rect 567750 159200 567806 160000
rect 568670 159200 568726 160000
rect 569682 159200 569738 160000
rect 570694 159200 570750 160000
rect 571352 159310 571564 159338
rect 489656 159174 489776 159200
rect 490656 156800 490708 156806
rect 490656 156742 490708 156748
rect 489644 154216 489696 154222
rect 489644 154158 489696 154164
rect 489276 152788 489328 152794
rect 489276 152730 489328 152736
rect 489368 152788 489420 152794
rect 489368 152730 489420 152736
rect 489380 151994 489408 152730
rect 488368 151966 488428 151994
rect 489072 151966 489408 151994
rect 489656 151994 489684 154158
rect 490668 151994 490696 156742
rect 490760 155990 490788 159200
rect 490748 155984 490800 155990
rect 490748 155926 490800 155932
rect 491208 155372 491260 155378
rect 491208 155314 491260 155320
rect 491220 151994 491248 155314
rect 491680 152726 491708 159200
rect 492692 156738 492720 159200
rect 492680 156732 492732 156738
rect 492680 156674 492732 156680
rect 493324 156732 493376 156738
rect 493324 156674 493376 156680
rect 492588 154148 492640 154154
rect 492588 154090 492640 154096
rect 491668 152720 491720 152726
rect 491668 152662 491720 152668
rect 491944 152720 491996 152726
rect 491944 152662 491996 152668
rect 491956 151994 491984 152662
rect 492600 151994 492628 154090
rect 493336 151994 493364 156674
rect 493704 152114 493732 159200
rect 494624 156126 494652 159200
rect 494612 156120 494664 156126
rect 494612 156062 494664 156068
rect 494610 155952 494666 155961
rect 494610 155887 494666 155896
rect 493966 155816 494022 155825
rect 493966 155751 494022 155760
rect 493692 152108 493744 152114
rect 493692 152050 493744 152056
rect 493980 151994 494008 155751
rect 494624 151994 494652 155887
rect 495256 154080 495308 154086
rect 495256 154022 495308 154028
rect 495268 151994 495296 154022
rect 495636 152590 495664 159200
rect 496556 155938 496584 159200
rect 497568 156194 497596 159200
rect 497556 156188 497608 156194
rect 497556 156130 497608 156136
rect 496464 155910 496584 155938
rect 495900 152652 495952 152658
rect 495900 152594 495952 152600
rect 495624 152584 495676 152590
rect 495624 152526 495676 152532
rect 495912 151994 495940 152594
rect 496464 152590 496492 155910
rect 497186 155680 497242 155689
rect 497186 155615 497242 155624
rect 496542 155544 496598 155553
rect 496542 155479 496598 155488
rect 496452 152584 496504 152590
rect 496452 152526 496504 152532
rect 496556 151994 496584 155479
rect 497200 151994 497228 155615
rect 497832 154012 497884 154018
rect 497832 153954 497884 153960
rect 497844 151994 497872 153954
rect 498108 152584 498160 152590
rect 498108 152526 498160 152532
rect 489656 151966 489716 151994
rect 490360 151966 490696 151994
rect 491004 151966 491248 151994
rect 491648 151966 491984 151994
rect 492292 151966 492628 151994
rect 493028 151966 493364 151994
rect 493672 151966 494008 151994
rect 494316 151966 494652 151994
rect 494960 151966 495296 151994
rect 495604 151966 495940 151994
rect 496248 151966 496584 151994
rect 496892 151966 497228 151994
rect 497536 151966 497872 151994
rect 498120 151994 498148 152526
rect 498580 152182 498608 159200
rect 499500 156262 499528 159200
rect 499488 156256 499540 156262
rect 499488 156198 499540 156204
rect 499394 155408 499450 155417
rect 499394 155343 499450 155352
rect 499120 153944 499172 153950
rect 499120 153886 499172 153892
rect 498568 152176 498620 152182
rect 498568 152118 498620 152124
rect 499132 151994 499160 153886
rect 498120 151966 498180 151994
rect 498824 151966 499160 151994
rect 499408 151994 499436 155343
rect 500408 154488 500460 154494
rect 500408 154430 500460 154436
rect 500420 151994 500448 154430
rect 500512 152250 500540 159200
rect 500866 155272 500922 155281
rect 501432 155242 501460 159200
rect 502444 155938 502472 159200
rect 502168 155910 502472 155938
rect 500866 155207 500922 155216
rect 501420 155236 501472 155242
rect 500500 152244 500552 152250
rect 500500 152186 500552 152192
rect 500880 151994 500908 155207
rect 501420 155178 501472 155184
rect 501696 153876 501748 153882
rect 501696 153818 501748 153824
rect 501708 151994 501736 153818
rect 502168 153474 502196 155910
rect 503076 155236 503128 155242
rect 503076 155178 503128 155184
rect 502248 153536 502300 153542
rect 502248 153478 502300 153484
rect 502156 153468 502208 153474
rect 502156 153410 502208 153416
rect 502260 151994 502288 153478
rect 503088 151994 503116 155178
rect 503364 153406 503392 159200
rect 504376 156670 504404 159200
rect 504364 156664 504416 156670
rect 504364 156606 504416 156612
rect 505388 154630 505416 159200
rect 505376 154624 505428 154630
rect 505376 154566 505428 154572
rect 506308 153610 506336 159200
rect 506296 153604 506348 153610
rect 506296 153546 506348 153552
rect 503352 153400 503404 153406
rect 503352 153342 503404 153348
rect 506478 153232 506534 153241
rect 506478 153167 506534 153176
rect 499408 151966 499468 151994
rect 500112 151966 500448 151994
rect 500756 151966 500908 151994
rect 501400 151966 501736 151994
rect 502136 151966 502288 151994
rect 502780 151966 503116 151994
rect 505650 152008 505706 152017
rect 506492 151994 506520 153167
rect 507320 152522 507348 159200
rect 508240 154834 508268 159200
rect 508780 156664 508832 156670
rect 508780 156606 508832 156612
rect 508228 154828 508280 154834
rect 508228 154770 508280 154776
rect 507308 152516 507360 152522
rect 507308 152458 507360 152464
rect 508792 151994 508820 156606
rect 509252 154766 509280 159200
rect 510264 156330 510292 159200
rect 510252 156324 510304 156330
rect 510252 156266 510304 156272
rect 509240 154760 509292 154766
rect 509240 154702 509292 154708
rect 511184 154698 511212 159200
rect 511540 157412 511592 157418
rect 511540 157354 511592 157360
rect 511172 154692 511224 154698
rect 511172 154634 511224 154640
rect 510894 153368 510950 153377
rect 510894 153303 510950 153312
rect 508870 153232 508926 153241
rect 508870 153167 508926 153176
rect 505706 151966 506000 151994
rect 506492 151966 506644 151994
rect 508576 151966 508820 151994
rect 508884 151994 508912 153167
rect 510160 152516 510212 152522
rect 510160 152458 510212 152464
rect 510172 151994 510200 152458
rect 508884 151966 509220 151994
rect 509864 151966 510200 151994
rect 510908 151994 510936 153303
rect 511552 151994 511580 157354
rect 512196 155038 512224 159200
rect 512184 155032 512236 155038
rect 512184 154974 512236 154980
rect 512182 153504 512238 153513
rect 512182 153439 512238 153448
rect 512196 151994 512224 153439
rect 513116 152318 513144 159200
rect 514128 154902 514156 159200
rect 515140 155106 515168 159200
rect 515128 155100 515180 155106
rect 515128 155042 515180 155048
rect 516060 154970 516088 159200
rect 516048 154964 516100 154970
rect 516048 154906 516100 154912
rect 514116 154896 514168 154902
rect 514116 154838 514168 154844
rect 516690 154048 516746 154057
rect 516690 153983 516746 153992
rect 516138 153912 516194 153921
rect 516138 153847 516194 153856
rect 514758 153776 514814 153785
rect 514758 153711 514814 153720
rect 513470 153640 513526 153649
rect 513470 153575 513526 153584
rect 513104 152312 513156 152318
rect 513104 152254 513156 152260
rect 513484 151994 513512 153575
rect 514668 153332 514720 153338
rect 514668 153274 514720 153280
rect 514680 151994 514708 153274
rect 510908 151966 511244 151994
rect 511552 151966 511888 151994
rect 512196 151966 512532 151994
rect 513484 151966 513820 151994
rect 514464 151966 514708 151994
rect 514772 151994 514800 153711
rect 516048 153264 516100 153270
rect 516048 153206 516100 153212
rect 516060 151994 516088 153206
rect 514772 151966 515108 151994
rect 515752 151966 516088 151994
rect 516152 151994 516180 153847
rect 516704 151994 516732 153983
rect 517072 153678 517100 159200
rect 517992 156534 518020 159200
rect 517980 156528 518032 156534
rect 517980 156470 518032 156476
rect 519004 155922 519032 159200
rect 518992 155916 519044 155922
rect 518992 155858 519044 155864
rect 520016 155174 520044 159200
rect 520004 155168 520056 155174
rect 520004 155110 520056 155116
rect 517978 154184 518034 154193
rect 517978 154119 518034 154128
rect 517060 153672 517112 153678
rect 517060 153614 517112 153620
rect 517992 151994 518020 154119
rect 520936 153746 520964 159200
rect 520924 153740 520976 153746
rect 520924 153682 520976 153688
rect 520556 153332 520608 153338
rect 520556 153274 520608 153280
rect 516152 151966 516396 151994
rect 516704 151966 517040 151994
rect 517992 151966 518328 151994
rect 505650 151943 505706 151952
rect 503628 151904 503680 151910
rect 442828 151830 442888 151858
rect 477328 151830 477388 151858
rect 503424 151852 503628 151858
rect 520280 151904 520332 151910
rect 519266 151872 519322 151881
rect 503424 151846 503680 151852
rect 503424 151830 503668 151846
rect 504712 151842 505048 151858
rect 504712 151836 505060 151842
rect 504712 151830 505008 151836
rect 252008 151778 252060 151784
rect 519322 151830 519616 151858
rect 520280 151846 520332 151852
rect 519266 151807 519322 151816
rect 505008 151778 505060 151784
rect 507780 151570 507932 151586
rect 507768 151564 507932 151570
rect 507820 151558 507932 151564
rect 507768 151506 507820 151512
rect 505652 151496 505704 151502
rect 177224 151434 177560 151450
rect 177212 151428 177560 151434
rect 177264 151422 177560 151428
rect 505356 151444 505652 151450
rect 513288 151496 513340 151502
rect 505356 151438 505704 151444
rect 505356 151422 505692 151438
rect 506952 151434 507288 151450
rect 506940 151428 507288 151434
rect 177212 151370 177264 151376
rect 506992 151422 507288 151428
rect 513176 151444 513288 151450
rect 513176 151438 513340 151444
rect 513176 151422 513328 151438
rect 517684 151434 518020 151450
rect 517684 151428 518032 151434
rect 517684 151422 517980 151428
rect 506940 151370 506992 151376
rect 517980 151370 518032 151376
rect 503720 151360 503772 151366
rect 510160 151360 510212 151366
rect 503772 151308 504068 151314
rect 503720 151302 504068 151308
rect 519268 151360 519320 151366
rect 510212 151308 510508 151314
rect 510160 151302 510508 151308
rect 503732 151286 504068 151302
rect 510172 151286 510508 151302
rect 518972 151308 519268 151314
rect 518972 151302 519320 151308
rect 518972 151286 519308 151302
rect 119712 151224 119764 151230
rect 119712 151166 119764 151172
rect 119620 2916 119672 2922
rect 119620 2858 119672 2864
rect 119526 2680 119582 2689
rect 119526 2615 119582 2624
rect 119342 2408 119398 2417
rect 119342 2343 119398 2352
rect 118148 1760 118200 1766
rect 118148 1702 118200 1708
rect 119632 800 119660 2858
rect 119724 2553 119752 151166
rect 519728 150952 519780 150958
rect 519728 150894 519780 150900
rect 519740 149025 519768 150894
rect 519726 149016 519782 149025
rect 519726 148951 519782 148960
rect 474476 4690 474628 4706
rect 168840 4684 168892 4690
rect 168840 4626 168892 4632
rect 474464 4684 474628 4690
rect 474516 4678 474628 4684
rect 518624 4684 518676 4690
rect 474464 4626 474516 4632
rect 518624 4626 518676 4632
rect 519636 4684 519688 4690
rect 519636 4626 519688 4632
rect 121472 4134 121716 4162
rect 124692 4146 125028 4162
rect 124680 4140 125028 4146
rect 121472 2854 121500 4134
rect 124732 4134 125028 4140
rect 125140 4140 125192 4146
rect 124680 4082 124732 4088
rect 125140 4082 125192 4088
rect 128372 4134 128432 4162
rect 130292 4140 130344 4146
rect 121460 2848 121512 2854
rect 121460 2790 121512 2796
rect 119710 2544 119766 2553
rect 119710 2479 119766 2488
rect 125152 2122 125180 4082
rect 128372 3534 128400 4134
rect 130292 4082 130344 4088
rect 131408 4134 131744 4162
rect 134812 4134 135148 4162
rect 138124 4134 138460 4162
rect 141528 4134 141864 4162
rect 144932 4134 145176 4162
rect 148244 4134 148580 4162
rect 151832 4134 151892 4162
rect 154960 4134 155296 4162
rect 158272 4134 158608 4162
rect 161676 4134 162012 4162
rect 164988 4134 165324 4162
rect 168392 4134 168728 4162
rect 128360 3528 128412 3534
rect 128360 3470 128412 3476
rect 124968 2094 125180 2122
rect 124968 800 124996 2094
rect 130304 800 130332 4082
rect 131408 2854 131436 4134
rect 134812 3194 134840 4134
rect 138124 3262 138152 4134
rect 140872 3528 140924 3534
rect 140872 3470 140924 3476
rect 138112 3256 138164 3262
rect 138112 3198 138164 3204
rect 134800 3188 134852 3194
rect 134800 3130 134852 3136
rect 135536 3188 135588 3194
rect 135536 3130 135588 3136
rect 131396 2848 131448 2854
rect 131396 2790 131448 2796
rect 135548 800 135576 3130
rect 140884 800 140912 3470
rect 141528 2718 141556 4134
rect 141608 3596 141660 3602
rect 141608 3538 141660 3544
rect 141620 2718 141648 3538
rect 144932 2786 144960 4134
rect 146944 3664 146996 3670
rect 146944 3606 146996 3612
rect 146208 3256 146260 3262
rect 146208 3198 146260 3204
rect 144920 2780 144972 2786
rect 144920 2722 144972 2728
rect 141516 2712 141568 2718
rect 141516 2654 141568 2660
rect 141608 2712 141660 2718
rect 141608 2654 141660 2660
rect 146220 800 146248 3198
rect 146956 2786 146984 3606
rect 146944 2780 146996 2786
rect 146944 2722 146996 2728
rect 148244 2718 148272 4134
rect 151544 3664 151596 3670
rect 151544 3606 151596 3612
rect 148232 2712 148284 2718
rect 148232 2654 148284 2660
rect 151556 800 151584 3606
rect 151832 2786 151860 4134
rect 154960 3738 154988 4134
rect 158272 3806 158300 4134
rect 158260 3800 158312 3806
rect 158260 3742 158312 3748
rect 154948 3732 155000 3738
rect 154948 3674 155000 3680
rect 156880 2848 156932 2854
rect 156880 2790 156932 2796
rect 151820 2780 151872 2786
rect 151820 2722 151872 2728
rect 156892 800 156920 2790
rect 71596 128 71648 134
rect 71596 70 71648 76
rect 71686 0 71742 800
rect 77022 0 77078 800
rect 82358 0 82414 800
rect 87694 0 87750 800
rect 93030 0 93086 800
rect 98366 0 98422 800
rect 103610 0 103666 800
rect 108946 0 109002 800
rect 114282 0 114338 800
rect 119618 0 119674 800
rect 124954 0 125010 800
rect 130290 0 130346 800
rect 135534 0 135590 800
rect 140870 0 140926 800
rect 146206 0 146262 800
rect 151542 0 151598 800
rect 156878 0 156934 800
rect 161676 134 161704 4134
rect 164988 3942 165016 4134
rect 164976 3936 165028 3942
rect 168392 3890 168420 4134
rect 164976 3878 165028 3884
rect 168300 3874 168420 3890
rect 168288 3868 168420 3874
rect 168340 3862 168420 3868
rect 168288 3810 168340 3816
rect 162216 3800 162268 3806
rect 162216 3742 162268 3748
rect 167460 3800 167512 3806
rect 167460 3742 167512 3748
rect 162228 800 162256 3742
rect 167472 800 167500 3742
rect 168852 1698 168880 4626
rect 171796 4134 172132 4162
rect 175292 4134 175444 4162
rect 178512 4134 178848 4162
rect 181824 4134 182160 4162
rect 188540 4134 188876 4162
rect 191944 4134 192280 4162
rect 195256 4134 195592 4162
rect 198752 4146 198996 4162
rect 198740 4140 198996 4146
rect 171796 3330 171824 4134
rect 175292 3398 175320 4134
rect 178132 3868 178184 3874
rect 178132 3810 178184 3816
rect 175280 3392 175332 3398
rect 175280 3334 175332 3340
rect 176660 3392 176712 3398
rect 176660 3334 176712 3340
rect 171784 3324 171836 3330
rect 171784 3266 171836 3272
rect 172796 3324 172848 3330
rect 172796 3266 172848 3272
rect 168840 1692 168892 1698
rect 168840 1634 168892 1640
rect 172808 800 172836 3266
rect 176672 1630 176700 3334
rect 176660 1624 176712 1630
rect 176660 1566 176712 1572
rect 178144 800 178172 3810
rect 178512 3466 178540 4134
rect 178500 3460 178552 3466
rect 178500 3402 178552 3408
rect 181824 2990 181852 4134
rect 183468 3188 183520 3194
rect 183468 3130 183520 3136
rect 181812 2984 181864 2990
rect 181812 2926 181864 2932
rect 183480 800 183508 3130
rect 188540 3058 188568 4134
rect 188804 3256 188856 3262
rect 188804 3198 188856 3204
rect 188528 3052 188580 3058
rect 188528 2994 188580 3000
rect 188816 800 188844 3198
rect 191944 3126 191972 4134
rect 195256 4078 195284 4134
rect 198792 4134 198996 4140
rect 201972 4134 202308 4162
rect 205652 4134 205712 4162
rect 208688 4134 209024 4162
rect 212092 4134 212428 4162
rect 215496 4134 215832 4162
rect 198740 4082 198792 4088
rect 195244 4072 195296 4078
rect 195244 4014 195296 4020
rect 201972 3534 202000 4134
rect 205652 3602 205680 4134
rect 208688 3670 208716 4134
rect 212092 3738 212120 4134
rect 215392 4072 215444 4078
rect 215392 4014 215444 4020
rect 212080 3732 212132 3738
rect 212080 3674 212132 3680
rect 208676 3664 208728 3670
rect 208676 3606 208728 3612
rect 205640 3596 205692 3602
rect 205640 3538 205692 3544
rect 201960 3528 202012 3534
rect 201960 3470 202012 3476
rect 213828 3528 213880 3534
rect 213828 3470 213880 3476
rect 210056 3324 210108 3330
rect 210056 3266 210108 3272
rect 191932 3120 191984 3126
rect 191932 3062 191984 3068
rect 204720 3120 204772 3126
rect 204720 3062 204772 3068
rect 199384 3052 199436 3058
rect 199384 2994 199436 3000
rect 194140 2984 194192 2990
rect 194140 2926 194192 2932
rect 194152 800 194180 2926
rect 199396 800 199424 2994
rect 204732 800 204760 3062
rect 210068 800 210096 3266
rect 213840 1562 213868 3470
rect 213828 1556 213880 1562
rect 213828 1498 213880 1504
rect 215404 800 215432 4014
rect 215496 2854 215524 4134
rect 219130 3942 219158 4148
rect 222212 4134 222548 4162
rect 225524 4134 225860 4162
rect 229112 4134 229264 4162
rect 232240 4134 232576 4162
rect 235644 4134 235980 4162
rect 238956 4134 239292 4162
rect 242360 4134 242696 4162
rect 245672 4134 246008 4162
rect 249076 4134 249412 4162
rect 252572 4134 252724 4162
rect 255792 4134 256128 4162
rect 259472 4134 259532 4162
rect 262508 4134 262844 4162
rect 265912 4134 266248 4162
rect 269224 4134 269560 4162
rect 272628 4134 272964 4162
rect 276032 4134 276276 4162
rect 279344 4134 279680 4162
rect 282932 4134 282992 4162
rect 286060 4134 286396 4162
rect 289372 4134 289708 4162
rect 292776 4134 293112 4162
rect 296088 4134 296424 4162
rect 299492 4134 299828 4162
rect 302896 4134 303232 4162
rect 306392 4134 306544 4162
rect 309612 4134 309948 4162
rect 219118 3936 219170 3942
rect 219118 3878 219170 3884
rect 222212 3806 222240 4134
rect 222200 3800 222252 3806
rect 222200 3742 222252 3748
rect 225524 3398 225552 4134
rect 229112 3874 229140 4134
rect 229100 3868 229152 3874
rect 229100 3810 229152 3816
rect 226064 3664 226116 3670
rect 226064 3606 226116 3612
rect 225512 3392 225564 3398
rect 225512 3334 225564 3340
rect 215484 2848 215536 2854
rect 215484 2790 215536 2796
rect 220728 2848 220780 2854
rect 220728 2790 220780 2796
rect 220740 800 220768 2790
rect 226076 800 226104 3606
rect 231308 3392 231360 3398
rect 231308 3334 231360 3340
rect 231320 800 231348 3334
rect 232240 3194 232268 4134
rect 235644 3262 235672 4134
rect 235632 3256 235684 3262
rect 235632 3198 235684 3204
rect 236644 3256 236696 3262
rect 236644 3198 236696 3204
rect 232228 3188 232280 3194
rect 232228 3130 232280 3136
rect 236656 800 236684 3198
rect 238956 2990 238984 4134
rect 241980 3732 242032 3738
rect 241980 3674 242032 3680
rect 238944 2984 238996 2990
rect 238944 2926 238996 2932
rect 241992 800 242020 3674
rect 242360 3058 242388 4134
rect 245672 3126 245700 4134
rect 249076 3330 249104 4134
rect 252572 4078 252600 4134
rect 252560 4072 252612 4078
rect 252560 4014 252612 4020
rect 249064 3324 249116 3330
rect 249064 3266 249116 3272
rect 245660 3120 245712 3126
rect 245660 3062 245712 3068
rect 247316 3120 247368 3126
rect 247316 3062 247368 3068
rect 242348 3052 242400 3058
rect 242348 2994 242400 3000
rect 247328 800 247356 3062
rect 252652 3052 252704 3058
rect 252652 2994 252704 3000
rect 252664 800 252692 2994
rect 255792 2854 255820 4134
rect 259472 3670 259500 4134
rect 259460 3664 259512 3670
rect 259460 3606 259512 3612
rect 262508 3398 262536 4134
rect 262496 3392 262548 3398
rect 262496 3334 262548 3340
rect 265912 3262 265940 4134
rect 269224 3738 269252 4134
rect 269212 3732 269264 3738
rect 269212 3674 269264 3680
rect 265900 3256 265952 3262
rect 265900 3198 265952 3204
rect 257988 3188 258040 3194
rect 257988 3130 258040 3136
rect 255780 2848 255832 2854
rect 255780 2790 255832 2796
rect 258000 800 258028 3130
rect 272628 3126 272656 4134
rect 272616 3120 272668 3126
rect 272616 3062 272668 3068
rect 273904 3120 273956 3126
rect 273904 3062 273956 3068
rect 263232 2984 263284 2990
rect 263232 2926 263284 2932
rect 263244 800 263272 2926
rect 268568 2848 268620 2854
rect 268568 2790 268620 2796
rect 268580 800 268608 2790
rect 273916 800 273944 3062
rect 276032 3058 276060 4134
rect 279344 3194 279372 4134
rect 279332 3188 279384 3194
rect 279332 3130 279384 3136
rect 276020 3052 276072 3058
rect 276020 2994 276072 3000
rect 279240 3052 279292 3058
rect 279240 2994 279292 3000
rect 279252 800 279280 2994
rect 282932 2990 282960 4134
rect 282920 2984 282972 2990
rect 282920 2926 282972 2932
rect 284576 2848 284628 2854
rect 284576 2790 284628 2796
rect 284588 800 284616 2790
rect 286060 2786 286088 4134
rect 289372 3126 289400 4134
rect 289360 3120 289412 3126
rect 289360 3062 289412 3068
rect 292776 3058 292804 4134
rect 292764 3052 292816 3058
rect 292764 2994 292816 3000
rect 295156 3052 295208 3058
rect 295156 2994 295208 3000
rect 289912 2984 289964 2990
rect 289912 2926 289964 2932
rect 286048 2780 286100 2786
rect 286048 2722 286100 2728
rect 289924 800 289952 2926
rect 295168 800 295196 2994
rect 296088 2786 296116 4134
rect 299492 2990 299520 4134
rect 302896 3058 302924 4134
rect 302884 3052 302936 3058
rect 302884 2994 302936 3000
rect 299480 2984 299532 2990
rect 299480 2926 299532 2932
rect 300492 2848 300544 2854
rect 300492 2790 300544 2796
rect 305828 2848 305880 2854
rect 305828 2790 305880 2796
rect 296076 2780 296128 2786
rect 296076 2722 296128 2728
rect 300504 800 300532 2790
rect 305840 800 305868 2790
rect 306392 2786 306420 4134
rect 309612 2854 309640 4134
rect 313246 3942 313274 4148
rect 316512 4134 316664 4162
rect 319976 4134 320220 4162
rect 323380 4134 323716 4162
rect 326692 4134 327028 4162
rect 330096 4134 330432 4162
rect 333408 4134 333744 4162
rect 336812 4134 337148 4162
rect 340124 4134 340460 4162
rect 311164 3936 311216 3942
rect 311164 3878 311216 3884
rect 313234 3936 313286 3942
rect 313234 3878 313286 3884
rect 309600 2848 309652 2854
rect 309600 2790 309652 2796
rect 306380 2780 306432 2786
rect 306380 2722 306432 2728
rect 311176 800 311204 3878
rect 316512 800 316540 4134
rect 320192 2854 320220 4134
rect 320180 2848 320232 2854
rect 320180 2790 320232 2796
rect 321836 2848 321888 2854
rect 321836 2790 321888 2796
rect 321848 800 321876 2790
rect 323688 2786 323716 4134
rect 327000 2938 327028 4134
rect 327000 2910 327120 2938
rect 327092 2854 327120 2910
rect 327080 2848 327132 2854
rect 327080 2790 327132 2796
rect 330404 2786 330432 4134
rect 332416 2848 332468 2854
rect 332416 2790 332468 2796
rect 323676 2780 323728 2786
rect 323676 2722 323728 2728
rect 330392 2780 330444 2786
rect 330392 2722 330444 2728
rect 327080 2712 327132 2718
rect 327080 2654 327132 2660
rect 327092 800 327120 2654
rect 332428 800 332456 2790
rect 333716 1630 333744 4134
rect 337120 2718 337148 4134
rect 337752 2848 337804 2854
rect 337752 2790 337804 2796
rect 337108 2712 337160 2718
rect 337108 2654 337160 2660
rect 333704 1624 333756 1630
rect 333704 1566 333756 1572
rect 337764 800 337792 2790
rect 340432 1562 340460 4134
rect 343468 4134 343528 4162
rect 346932 4134 347268 4162
rect 350244 4134 350488 4162
rect 353648 4134 353984 4162
rect 356960 4134 357296 4162
rect 360364 4134 360700 4162
rect 363676 4134 364012 4162
rect 343468 1630 343496 4134
rect 347240 3126 347268 4134
rect 347228 3120 347280 3126
rect 347228 3062 347280 3068
rect 350460 2854 350488 4134
rect 353956 3262 353984 4134
rect 353944 3256 353996 3262
rect 353944 3198 353996 3204
rect 357268 3058 357296 4134
rect 360672 3398 360700 4134
rect 360660 3392 360712 3398
rect 360660 3334 360712 3340
rect 357256 3052 357308 3058
rect 357256 2994 357308 3000
rect 363984 2990 364012 4134
rect 367020 4134 367080 4162
rect 370392 4134 370728 4162
rect 373796 4134 373948 4162
rect 377108 4134 377444 4162
rect 380512 4134 380848 4162
rect 383824 4134 384160 4162
rect 387228 4134 387564 4162
rect 390632 4134 390968 4162
rect 393944 4134 394280 4162
rect 367020 3670 367048 4134
rect 367008 3664 367060 3670
rect 367008 3606 367060 3612
rect 370700 3330 370728 4134
rect 373920 3602 373948 4134
rect 373908 3596 373960 3602
rect 373908 3538 373960 3544
rect 370688 3324 370740 3330
rect 370688 3266 370740 3272
rect 377416 3262 377444 4134
rect 375012 3256 375064 3262
rect 375012 3198 375064 3204
rect 377404 3256 377456 3262
rect 377404 3198 377456 3204
rect 364340 3120 364392 3126
rect 364340 3062 364392 3068
rect 363972 2984 364024 2990
rect 363972 2926 364024 2932
rect 350448 2848 350500 2854
rect 350448 2790 350500 2796
rect 348424 2712 348476 2718
rect 348424 2654 348476 2660
rect 343088 1624 343140 1630
rect 343088 1566 343140 1572
rect 343456 1624 343508 1630
rect 343456 1566 343508 1572
rect 340420 1556 340472 1562
rect 340420 1498 340472 1504
rect 343100 800 343128 1566
rect 348436 800 348464 2654
rect 359004 1624 359056 1630
rect 359004 1566 359056 1572
rect 353760 1556 353812 1562
rect 353760 1498 353812 1504
rect 353772 800 353800 1498
rect 359016 800 359044 1566
rect 364352 800 364380 3062
rect 369676 2848 369728 2854
rect 369676 2790 369728 2796
rect 369688 800 369716 2790
rect 375024 800 375052 3198
rect 380348 3052 380400 3058
rect 380348 2994 380400 3000
rect 380360 800 380388 2994
rect 380820 2854 380848 4134
rect 384132 3194 384160 4134
rect 385684 3392 385736 3398
rect 385684 3334 385736 3340
rect 384120 3188 384172 3194
rect 384120 3130 384172 3136
rect 380808 2848 380860 2854
rect 380808 2790 380860 2796
rect 385696 800 385724 3334
rect 387536 3126 387564 4134
rect 387524 3120 387576 3126
rect 387524 3062 387576 3068
rect 390940 3058 390968 4134
rect 394252 3398 394280 4134
rect 397288 4134 397348 4162
rect 400660 4134 400996 4162
rect 404064 4146 404308 4162
rect 404064 4140 404320 4146
rect 404064 4134 404268 4140
rect 396264 3664 396316 3670
rect 396264 3606 396316 3612
rect 394240 3392 394292 3398
rect 394240 3334 394292 3340
rect 390928 3052 390980 3058
rect 390928 2994 390980 3000
rect 390836 2984 390888 2990
rect 390836 2926 390888 2932
rect 390848 1578 390876 2926
rect 390848 1550 390968 1578
rect 390940 800 390968 1550
rect 396276 800 396304 3606
rect 397288 2990 397316 4134
rect 400968 3330 400996 4134
rect 407376 4134 407712 4162
rect 410780 4134 411116 4162
rect 404268 4082 404320 4088
rect 407684 4078 407712 4134
rect 407672 4072 407724 4078
rect 407672 4014 407724 4020
rect 411088 3738 411116 4134
rect 414078 3942 414106 4148
rect 417496 4134 417832 4162
rect 414066 3936 414118 3942
rect 414066 3878 414118 3884
rect 417804 3874 417832 4134
rect 420748 4134 420808 4162
rect 424212 4134 424548 4162
rect 427524 4134 427768 4162
rect 430928 4134 431264 4162
rect 434332 4134 434668 4162
rect 437644 4134 437980 4162
rect 441048 4134 441292 4162
rect 417792 3868 417844 3874
rect 417792 3810 417844 3816
rect 420748 3806 420776 4134
rect 420736 3800 420788 3806
rect 420736 3742 420788 3748
rect 411076 3732 411128 3738
rect 411076 3674 411128 3680
rect 424520 3670 424548 4134
rect 401600 3664 401652 3670
rect 401600 3606 401652 3612
rect 424508 3664 424560 3670
rect 424508 3606 424560 3612
rect 400956 3324 401008 3330
rect 400956 3266 401008 3272
rect 397276 2984 397328 2990
rect 397276 2926 397328 2932
rect 401612 800 401640 3606
rect 427740 3602 427768 4134
rect 406936 3596 406988 3602
rect 406936 3538 406988 3544
rect 427728 3596 427780 3602
rect 427728 3538 427780 3544
rect 406948 800 406976 3538
rect 426346 3496 426402 3505
rect 426346 3431 426402 3440
rect 412272 3256 412324 3262
rect 412272 3198 412324 3204
rect 412284 800 412312 3198
rect 422852 3188 422904 3194
rect 422852 3130 422904 3136
rect 417608 2780 417660 2786
rect 417608 2722 417660 2728
rect 417620 800 417648 2722
rect 422864 800 422892 3130
rect 426360 2786 426388 3431
rect 431236 3330 431264 4134
rect 431224 3324 431276 3330
rect 431224 3266 431276 3272
rect 434640 3262 434668 4134
rect 434628 3256 434680 3262
rect 434628 3198 434680 3204
rect 428188 3120 428240 3126
rect 428188 3062 428240 3068
rect 426348 2780 426400 2786
rect 426348 2722 426400 2728
rect 428200 800 428228 3062
rect 433524 3052 433576 3058
rect 433524 2994 433576 3000
rect 433536 800 433564 2994
rect 437952 2718 437980 4134
rect 441264 3262 441292 4134
rect 444300 4134 444360 4162
rect 447764 4134 448100 4162
rect 451076 4134 451228 4162
rect 441252 3256 441304 3262
rect 441252 3198 441304 3204
rect 444300 3194 444328 4134
rect 438860 3188 438912 3194
rect 438860 3130 438912 3136
rect 444288 3188 444340 3194
rect 444288 3130 444340 3136
rect 437940 2712 437992 2718
rect 437940 2654 437992 2660
rect 438872 800 438900 3130
rect 448072 3126 448100 4134
rect 448060 3120 448112 3126
rect 448060 3062 448112 3068
rect 451200 3058 451228 4134
rect 454316 4140 454368 4146
rect 454480 4134 454816 4162
rect 454316 4082 454368 4088
rect 451188 3052 451240 3058
rect 451188 2994 451240 3000
rect 444196 2984 444248 2990
rect 444196 2926 444248 2932
rect 444208 800 444236 2926
rect 449532 2848 449584 2854
rect 449532 2790 449584 2796
rect 449544 800 449572 2790
rect 454328 898 454356 4082
rect 454788 2990 454816 4134
rect 457456 4134 457792 4162
rect 461196 4134 461532 4162
rect 454776 2984 454828 2990
rect 454776 2926 454828 2932
rect 454328 870 454448 898
rect 161664 128 161716 134
rect 161664 70 161716 76
rect 162214 0 162270 800
rect 167458 0 167514 800
rect 172794 0 172850 800
rect 178130 0 178186 800
rect 183466 0 183522 800
rect 188802 0 188858 800
rect 194138 0 194194 800
rect 199382 0 199438 800
rect 204718 0 204774 800
rect 210054 0 210110 800
rect 215390 0 215446 800
rect 220726 0 220782 800
rect 226062 0 226118 800
rect 231306 0 231362 800
rect 236642 0 236698 800
rect 241978 0 242034 800
rect 247314 0 247370 800
rect 252650 0 252706 800
rect 257986 0 258042 800
rect 263230 0 263286 800
rect 268566 0 268622 800
rect 273902 0 273958 800
rect 279238 0 279294 800
rect 284574 0 284630 800
rect 289910 0 289966 800
rect 295154 0 295210 800
rect 300490 0 300546 800
rect 305826 0 305882 800
rect 311162 0 311218 800
rect 316498 0 316554 800
rect 321834 0 321890 800
rect 327078 0 327134 800
rect 332414 0 332470 800
rect 337750 0 337806 800
rect 343086 0 343142 800
rect 348422 0 348478 800
rect 353758 0 353814 800
rect 359002 0 359058 800
rect 364338 0 364394 800
rect 369674 0 369730 800
rect 375010 0 375066 800
rect 380346 0 380402 800
rect 385682 0 385738 800
rect 390926 0 390982 800
rect 396262 0 396318 800
rect 401598 0 401654 800
rect 406934 0 406990 800
rect 412270 0 412326 800
rect 417606 0 417662 800
rect 422850 0 422906 800
rect 428186 0 428242 800
rect 433522 0 433578 800
rect 438858 0 438914 800
rect 444194 0 444250 800
rect 449530 0 449586 800
rect 454420 762 454448 870
rect 454696 870 454816 898
rect 454696 762 454724 870
rect 454788 800 454816 870
rect 454420 734 454724 762
rect 454774 0 454830 800
rect 457456 66 457484 4134
rect 461504 4078 461532 4134
rect 464172 4134 464508 4162
rect 467852 4134 467912 4162
rect 470888 4134 471224 4162
rect 477696 4134 478032 4162
rect 481008 4134 481344 4162
rect 484412 4134 484748 4162
rect 487724 4134 488060 4162
rect 491312 4134 491464 4162
rect 494440 4134 494776 4162
rect 497844 4134 498180 4162
rect 501156 4134 501492 4162
rect 504560 4134 504896 4162
rect 507872 4134 508208 4162
rect 511276 4134 511612 4162
rect 514772 4134 514924 4162
rect 517992 4134 518328 4162
rect 460112 4072 460164 4078
rect 460112 4014 460164 4020
rect 461492 4072 461544 4078
rect 461492 4014 461544 4020
rect 458180 2848 458232 2854
rect 458180 2790 458232 2796
rect 458192 2718 458220 2790
rect 458180 2712 458232 2718
rect 458180 2654 458232 2660
rect 460124 800 460152 4014
rect 464172 2922 464200 4134
rect 465448 3732 465500 3738
rect 465448 3674 465500 3680
rect 464160 2916 464212 2922
rect 464160 2858 464212 2864
rect 465460 800 465488 3674
rect 467852 2786 467880 4134
rect 470888 4010 470916 4134
rect 470876 4004 470928 4010
rect 470876 3946 470928 3952
rect 470784 3936 470836 3942
rect 470784 3878 470836 3884
rect 467840 2780 467892 2786
rect 467840 2722 467892 2728
rect 470796 800 470824 3878
rect 476120 3868 476172 3874
rect 476120 3810 476172 3816
rect 476132 800 476160 3810
rect 477696 2582 477724 4134
rect 477684 2576 477736 2582
rect 477684 2518 477736 2524
rect 481008 1698 481036 4134
rect 481456 3800 481508 3806
rect 481456 3742 481508 3748
rect 480996 1692 481048 1698
rect 480996 1634 481048 1640
rect 481468 800 481496 3742
rect 484412 1766 484440 4134
rect 486700 3664 486752 3670
rect 486700 3606 486752 3612
rect 484400 1760 484452 1766
rect 484400 1702 484452 1708
rect 486712 800 486740 3606
rect 487724 2514 487752 4134
rect 487712 2508 487764 2514
rect 487712 2450 487764 2456
rect 491312 1902 491340 4134
rect 492036 3596 492088 3602
rect 492036 3538 492088 3544
rect 491300 1896 491352 1902
rect 491300 1838 491352 1844
rect 492048 800 492076 3538
rect 494440 1834 494468 4134
rect 497372 3392 497424 3398
rect 497372 3334 497424 3340
rect 494428 1828 494480 1834
rect 494428 1770 494480 1776
rect 497384 800 497412 3334
rect 497844 1358 497872 4134
rect 501156 1970 501184 4134
rect 502708 3324 502760 3330
rect 502708 3266 502760 3272
rect 501144 1964 501196 1970
rect 501144 1906 501196 1912
rect 497832 1352 497884 1358
rect 497832 1294 497884 1300
rect 502720 800 502748 3266
rect 504560 2378 504588 4134
rect 504548 2372 504600 2378
rect 504548 2314 504600 2320
rect 507872 2242 507900 4134
rect 508044 3596 508096 3602
rect 508044 3538 508096 3544
rect 507860 2236 507912 2242
rect 507860 2178 507912 2184
rect 508056 800 508084 3538
rect 511276 2174 511304 4134
rect 513380 2848 513432 2854
rect 513380 2790 513432 2796
rect 511264 2168 511316 2174
rect 511264 2110 511316 2116
rect 513392 800 513420 2790
rect 514772 2038 514800 4134
rect 517992 2106 518020 4134
rect 517980 2100 518032 2106
rect 517980 2042 518032 2048
rect 514760 2032 514812 2038
rect 514760 1974 514812 1980
rect 518636 800 518664 4626
rect 519648 2650 519676 4626
rect 520096 4208 520148 4214
rect 520096 4150 520148 4156
rect 519636 2644 519688 2650
rect 519636 2586 519688 2592
rect 520108 1426 520136 4150
rect 520292 3602 520320 151846
rect 520372 151428 520424 151434
rect 520372 151370 520424 151376
rect 520280 3596 520332 3602
rect 520280 3538 520332 3544
rect 520384 2446 520412 151370
rect 520464 151360 520516 151366
rect 520464 151302 520516 151308
rect 520372 2440 520424 2446
rect 520372 2382 520424 2388
rect 520476 2310 520504 151302
rect 520568 4729 520596 153274
rect 520648 153264 520700 153270
rect 520648 153206 520700 153212
rect 520554 4720 520610 4729
rect 520554 4655 520610 4664
rect 520660 4457 520688 153206
rect 521948 153202 521976 159200
rect 522868 155854 522896 159200
rect 523880 156602 523908 159200
rect 523868 156596 523920 156602
rect 523868 156538 523920 156544
rect 522856 155848 522908 155854
rect 522856 155790 522908 155796
rect 524892 153814 524920 159200
rect 525812 155786 525840 159200
rect 525800 155780 525852 155786
rect 525800 155722 525852 155728
rect 526824 154562 526852 159200
rect 526812 154556 526864 154562
rect 526812 154498 526864 154504
rect 524880 153808 524932 153814
rect 524880 153750 524932 153756
rect 521936 153196 521988 153202
rect 521936 153138 521988 153144
rect 527744 153134 527772 159200
rect 527732 153128 527784 153134
rect 527732 153070 527784 153076
rect 528756 152386 528784 159200
rect 529768 157350 529796 159200
rect 529756 157344 529808 157350
rect 529756 157286 529808 157292
rect 530688 156466 530716 159200
rect 531700 157282 531728 159200
rect 531688 157276 531740 157282
rect 531688 157218 531740 157224
rect 530676 156460 530728 156466
rect 530676 156402 530728 156408
rect 532620 155718 532648 159200
rect 532608 155712 532660 155718
rect 532608 155654 532660 155660
rect 533632 153066 533660 159200
rect 533620 153060 533672 153066
rect 533620 153002 533672 153008
rect 534644 152454 534672 159200
rect 535564 157214 535592 159200
rect 535552 157208 535604 157214
rect 535552 157150 535604 157156
rect 536576 155650 536604 159200
rect 537496 157146 537524 159200
rect 537484 157140 537536 157146
rect 537484 157082 537536 157088
rect 538508 156398 538536 159200
rect 538496 156392 538548 156398
rect 538496 156334 538548 156340
rect 536564 155644 536616 155650
rect 536564 155586 536616 155592
rect 539520 152998 539548 159200
rect 540440 155582 540468 159200
rect 541452 157078 541480 159200
rect 541440 157072 541492 157078
rect 541440 157014 541492 157020
rect 540428 155576 540480 155582
rect 540428 155518 540480 155524
rect 542372 154578 542400 159200
rect 543384 157010 543412 159200
rect 543372 157004 543424 157010
rect 543372 156946 543424 156952
rect 544304 155446 544332 159200
rect 544292 155440 544344 155446
rect 544292 155382 544344 155388
rect 542280 154550 542400 154578
rect 542280 154426 542308 154550
rect 542268 154420 542320 154426
rect 542268 154362 542320 154368
rect 539508 152992 539560 152998
rect 539508 152934 539560 152940
rect 545316 152930 545344 159200
rect 546328 155514 546356 159200
rect 547248 156942 547276 159200
rect 547236 156936 547288 156942
rect 547236 156878 547288 156884
rect 548260 155922 548288 159200
rect 549180 156874 549208 159200
rect 549168 156868 549220 156874
rect 549168 156810 549220 156816
rect 546500 155916 546552 155922
rect 546500 155858 546552 155864
rect 548248 155916 548300 155922
rect 548248 155858 548300 155864
rect 546316 155508 546368 155514
rect 546316 155450 546368 155456
rect 546512 154358 546540 155858
rect 549168 155440 549220 155446
rect 549168 155382 549220 155388
rect 546500 154352 546552 154358
rect 546500 154294 546552 154300
rect 548524 154352 548576 154358
rect 548524 154294 548576 154300
rect 545304 152924 545356 152930
rect 545304 152866 545356 152872
rect 534632 152448 534684 152454
rect 534632 152390 534684 152396
rect 528744 152380 528796 152386
rect 528744 152322 528796 152328
rect 525064 151836 525116 151842
rect 525064 151778 525116 151784
rect 520740 151496 520792 151502
rect 520740 151438 520792 151444
rect 520646 4448 520702 4457
rect 520646 4383 520702 4392
rect 520464 2304 520516 2310
rect 520464 2246 520516 2252
rect 520752 1494 520780 151438
rect 522026 151056 522082 151065
rect 522026 150991 522082 151000
rect 521842 150920 521898 150929
rect 521842 150855 521898 150864
rect 520832 150748 520884 150754
rect 520832 150690 520884 150696
rect 520844 121553 520872 150690
rect 521752 150612 521804 150618
rect 521752 150554 521804 150560
rect 521658 141808 521714 141817
rect 521658 141743 521714 141752
rect 520830 121544 520886 121553
rect 520830 121479 520886 121488
rect 520830 94616 520886 94625
rect 520830 94551 520886 94560
rect 520844 4894 520872 94551
rect 521672 12986 521700 141743
rect 521764 108089 521792 150554
rect 521750 108080 521806 108089
rect 521750 108015 521806 108024
rect 521750 101416 521806 101425
rect 521750 101351 521806 101360
rect 521660 12980 521712 12986
rect 521660 12922 521712 12928
rect 521658 7304 521714 7313
rect 521658 7239 521714 7248
rect 521672 5001 521700 7239
rect 521764 5030 521792 101351
rect 521856 61033 521884 150855
rect 521936 150680 521988 150686
rect 521936 150622 521988 150628
rect 521948 114889 521976 150622
rect 521934 114880 521990 114889
rect 521934 114815 521990 114824
rect 521934 87952 521990 87961
rect 521934 87887 521990 87896
rect 521842 61024 521898 61033
rect 521842 60959 521898 60968
rect 521844 12980 521896 12986
rect 521844 12922 521896 12928
rect 521752 5024 521804 5030
rect 521658 4992 521714 5001
rect 521752 4966 521804 4972
rect 521658 4927 521714 4936
rect 520832 4888 520884 4894
rect 520832 4830 520884 4836
rect 521856 3534 521884 12922
rect 521948 4593 521976 87887
rect 522040 81297 522068 150991
rect 522120 150884 522172 150890
rect 522120 150826 522172 150832
rect 522132 135017 522160 150826
rect 522212 150816 522264 150822
rect 522212 150758 522264 150764
rect 522118 135008 522174 135017
rect 522118 134943 522174 134952
rect 522224 128353 522252 150758
rect 522210 128344 522266 128353
rect 522210 128279 522266 128288
rect 522026 81288 522082 81297
rect 522026 81223 522082 81232
rect 522026 74488 522082 74497
rect 522026 74423 522082 74432
rect 522040 4865 522068 74423
rect 522394 67824 522450 67833
rect 522394 67759 522450 67768
rect 522118 47560 522174 47569
rect 522118 47495 522174 47504
rect 522026 4856 522082 4865
rect 522026 4791 522082 4800
rect 521934 4584 521990 4593
rect 521934 4519 521990 4528
rect 522132 4214 522160 47495
rect 522210 27432 522266 27441
rect 522210 27367 522266 27376
rect 522120 4208 522172 4214
rect 522120 4150 522172 4156
rect 521844 3528 521896 3534
rect 521844 3470 521896 3476
rect 522224 3466 522252 27367
rect 522408 4690 522436 67759
rect 522580 34468 522632 34474
rect 522580 34410 522632 34416
rect 522592 34105 522620 34410
rect 522578 34096 522634 34105
rect 522578 34031 522634 34040
rect 522672 15156 522724 15162
rect 522672 15098 522724 15104
rect 522684 13977 522712 15098
rect 522670 13968 522726 13977
rect 522670 13903 522726 13912
rect 522396 4684 522448 4690
rect 522396 4626 522448 4632
rect 525076 3466 525104 151778
rect 527824 151156 527876 151162
rect 527824 151098 527876 151104
rect 527836 4146 527864 151098
rect 548536 34474 548564 154294
rect 549180 153542 549208 155382
rect 550192 154290 550220 159200
rect 550180 154284 550232 154290
rect 550180 154226 550232 154232
rect 549168 153536 549220 153542
rect 549168 153478 549220 153484
rect 551204 152862 551232 159200
rect 552124 155310 552152 159200
rect 552112 155304 552164 155310
rect 552112 155246 552164 155252
rect 551192 152856 551244 152862
rect 551192 152798 551244 152804
rect 553136 152794 553164 159200
rect 554056 154222 554084 159200
rect 555068 156806 555096 159200
rect 555056 156800 555108 156806
rect 555056 156742 555108 156748
rect 556080 155378 556108 159200
rect 556068 155372 556120 155378
rect 556068 155314 556120 155320
rect 554780 155304 554832 155310
rect 554780 155246 554832 155252
rect 554792 154494 554820 155246
rect 554780 154488 554832 154494
rect 554780 154430 554832 154436
rect 554044 154216 554096 154222
rect 554044 154158 554096 154164
rect 553124 152788 553176 152794
rect 553124 152730 553176 152736
rect 557000 152726 557028 159200
rect 558012 154154 558040 159200
rect 558932 156738 558960 159200
rect 558920 156732 558972 156738
rect 558920 156674 558972 156680
rect 559944 155825 559972 159200
rect 560956 155961 560984 159200
rect 560942 155952 560998 155961
rect 560942 155887 560998 155896
rect 559930 155816 559986 155825
rect 559930 155751 559986 155760
rect 561876 154714 561904 159200
rect 561600 154686 561904 154714
rect 558000 154148 558052 154154
rect 558000 154090 558052 154096
rect 561600 154086 561628 154686
rect 561588 154080 561640 154086
rect 561588 154022 561640 154028
rect 556988 152720 557040 152726
rect 556988 152662 557040 152668
rect 562888 152658 562916 159200
rect 563808 155553 563836 159200
rect 564820 155689 564848 159200
rect 564806 155680 564862 155689
rect 564806 155615 564862 155624
rect 563794 155544 563850 155553
rect 563794 155479 563850 155488
rect 565832 154578 565860 159200
rect 565740 154550 565860 154578
rect 565740 154018 565768 154550
rect 565728 154012 565780 154018
rect 565728 153954 565780 153960
rect 562876 152652 562928 152658
rect 562876 152594 562928 152600
rect 566752 152590 566780 159200
rect 567764 153950 567792 159200
rect 568684 155417 568712 159200
rect 568670 155408 568726 155417
rect 568670 155343 568726 155352
rect 569696 155310 569724 159200
rect 569684 155304 569736 155310
rect 570708 155281 570736 159200
rect 569684 155246 569736 155252
rect 570694 155272 570750 155281
rect 570694 155207 570750 155216
rect 571352 154578 571380 159310
rect 571536 159202 571564 159310
rect 571614 159202 571670 160000
rect 571536 159200 571670 159202
rect 572626 159200 572682 160000
rect 573546 159200 573602 160000
rect 574558 159200 574614 160000
rect 575570 159200 575626 160000
rect 576490 159200 576546 160000
rect 577502 159200 577558 160000
rect 578422 159200 578478 160000
rect 579434 159200 579490 160000
rect 571536 159174 571656 159200
rect 571984 155644 572036 155650
rect 571984 155586 572036 155592
rect 571260 154550 571380 154578
rect 567752 153944 567804 153950
rect 567752 153886 567804 153892
rect 571260 153882 571288 154550
rect 571248 153876 571300 153882
rect 571248 153818 571300 153824
rect 566740 152584 566792 152590
rect 566740 152526 566792 152532
rect 548524 34468 548576 34474
rect 548524 34410 548576 34416
rect 571996 5166 572024 155586
rect 572640 155446 572668 159200
rect 573364 155576 573416 155582
rect 573364 155518 573416 155524
rect 572628 155440 572680 155446
rect 572628 155382 572680 155388
rect 573376 15162 573404 155518
rect 573560 155242 573588 159200
rect 574572 155582 574600 159200
rect 574560 155576 574612 155582
rect 574560 155518 574612 155524
rect 573548 155236 573600 155242
rect 573548 155178 573600 155184
rect 575584 154358 575612 159200
rect 576504 155650 576532 159200
rect 577516 156670 577544 159200
rect 577504 156664 577556 156670
rect 577504 156606 577556 156612
rect 576492 155644 576544 155650
rect 576492 155586 576544 155592
rect 578436 154630 578464 159200
rect 578424 154624 578476 154630
rect 578424 154566 578476 154572
rect 575572 154352 575624 154358
rect 575572 154294 575624 154300
rect 579448 152425 579476 159200
rect 579434 152416 579490 152425
rect 579434 152351 579490 152360
rect 573364 15156 573416 15162
rect 573364 15098 573416 15104
rect 571984 5160 572036 5166
rect 571984 5102 572036 5108
rect 566556 4956 566608 4962
rect 566556 4898 566608 4904
rect 527824 4140 527876 4146
rect 527824 4082 527876 4088
rect 529296 4140 529348 4146
rect 529296 4082 529348 4088
rect 522212 3460 522264 3466
rect 522212 3402 522264 3408
rect 525064 3460 525116 3466
rect 525064 3402 525116 3408
rect 523960 3256 524012 3262
rect 523960 3198 524012 3204
rect 520740 1488 520792 1494
rect 520740 1430 520792 1436
rect 520096 1420 520148 1426
rect 520096 1362 520148 1368
rect 523972 800 524000 3198
rect 529308 800 529336 4082
rect 545304 4072 545356 4078
rect 545304 4014 545356 4020
rect 539968 3460 540020 3466
rect 539968 3402 540020 3408
rect 534632 3188 534684 3194
rect 534632 3130 534684 3136
rect 534644 800 534672 3130
rect 539980 800 540008 3402
rect 545316 800 545344 4014
rect 550546 3360 550602 3369
rect 550546 3295 550602 3304
rect 550560 800 550588 3295
rect 555884 3120 555936 3126
rect 555884 3062 555936 3068
rect 555896 800 555924 3062
rect 561220 3052 561272 3058
rect 561220 2994 561272 3000
rect 561232 800 561260 2994
rect 566568 800 566596 4898
rect 577228 4820 577280 4826
rect 577228 4762 577280 4768
rect 571892 2984 571944 2990
rect 571892 2926 571944 2932
rect 571904 800 571932 2926
rect 577240 800 577268 4762
rect 457444 60 457496 66
rect 457444 2 457496 8
rect 460110 0 460166 800
rect 465446 0 465502 800
rect 470782 0 470838 800
rect 476118 0 476174 800
rect 481454 0 481510 800
rect 486698 0 486754 800
rect 492034 0 492090 800
rect 497370 0 497426 800
rect 502706 0 502762 800
rect 508042 0 508098 800
rect 513378 0 513434 800
rect 518622 0 518678 800
rect 523958 0 524014 800
rect 529294 0 529350 800
rect 534630 0 534686 800
rect 539966 0 540022 800
rect 545302 0 545358 800
rect 550546 0 550602 800
rect 555882 0 555938 800
rect 561218 0 561274 800
rect 566554 0 566610 800
rect 571890 0 571946 800
rect 577226 0 577282 800
<< via2 >>
rect 1398 155216 1454 155272
rect 3146 157528 3202 157584
rect 2410 152496 2466 152552
rect 3330 156576 3386 156632
rect 5262 155352 5318 155408
rect 3238 152904 3294 152960
rect 3146 152360 3202 152416
rect 17866 156032 17922 156088
rect 17038 154264 17094 154320
rect 9402 153312 9458 153368
rect 19706 153176 19762 153232
rect 24766 155488 24822 155544
rect 30010 153448 30066 153504
rect 26606 153312 26662 153368
rect 2962 143792 3018 143848
rect 3330 149912 3386 149968
rect 3238 139304 3294 139360
rect 34702 156168 34758 156224
rect 36542 155624 36598 155680
rect 39854 153584 39910 153640
rect 37462 152632 37518 152688
rect 50158 156712 50214 156768
rect 52090 155760 52146 155816
rect 50618 153720 50674 153776
rect 64786 156848 64842 156904
rect 70582 154536 70638 154592
rect 75458 155896 75514 155952
rect 81162 153856 81218 153912
rect 88062 153992 88118 154048
rect 89166 156984 89222 157040
rect 91098 155080 91154 155136
rect 91926 154128 91982 154184
rect 3514 148416 3570 148472
rect 3330 134680 3386 134736
rect 3974 130056 4030 130112
rect 3882 125568 3938 125624
rect 3790 120944 3846 121000
rect 3698 116456 3754 116512
rect 3606 111832 3662 111888
rect 3514 107208 3570 107264
rect 3422 102720 3478 102776
rect 3790 98096 3846 98152
rect 3422 93608 3478 93664
rect 3330 66136 3386 66192
rect 3238 61512 3294 61568
rect 2778 57024 2834 57080
rect 3146 52400 3202 52456
rect 3054 47912 3110 47968
rect 2962 43288 3018 43344
rect 2870 38664 2926 38720
rect 2778 29552 2834 29608
rect 3238 6704 3294 6760
rect 3698 88984 3754 89040
rect 3606 84360 3662 84416
rect 3514 75248 3570 75304
rect 3882 79872 3938 79928
rect 3790 34176 3846 34232
rect 3698 25064 3754 25120
rect 3606 20440 3662 20496
rect 3974 70760 4030 70816
rect 3882 15816 3938 15872
rect 3974 11328 4030 11384
rect 33506 151408 33562 151464
rect 97906 154808 97962 154864
rect 105726 154944 105782 155000
rect 106186 154400 106242 154456
rect 108670 152904 108726 152960
rect 103794 152768 103850 152824
rect 102046 151816 102102 151872
rect 115754 152360 115810 152416
rect 98826 151408 98882 151464
rect 112442 151408 112498 151464
rect 23110 151272 23166 151328
rect 36910 151272 36966 151328
rect 53930 151272 53986 151328
rect 71318 151272 71374 151328
rect 92202 151272 92258 151328
rect 112442 150456 112498 150512
rect 113822 150592 113878 150648
rect 4802 6024 4858 6080
rect 3606 4936 3662 4992
rect 39302 4528 39358 4584
rect 45926 4528 45982 4584
rect 52458 4528 52514 4584
rect 75826 4392 75882 4448
rect 5998 2624 6054 2680
rect 2962 2216 3018 2272
rect 12346 2488 12402 2544
rect 28906 2352 28962 2408
rect 115202 150456 115258 150512
rect 116582 151136 116638 151192
rect 116490 89120 116546 89176
rect 116398 66408 116454 66464
rect 116030 9560 116086 9616
rect 116674 134680 116730 134736
rect 116766 131144 116822 131200
rect 116950 123256 117006 123312
rect 116858 121488 116914 121544
rect 116858 111968 116914 112024
rect 116950 111696 117006 111752
rect 118698 152360 118754 152416
rect 118146 151272 118202 151328
rect 117962 150728 118018 150784
rect 117778 150592 117834 150648
rect 117686 148144 117742 148200
rect 117226 146104 117282 146160
rect 117134 128696 117190 128752
rect 117134 106936 117190 106992
rect 117042 82592 117098 82648
rect 117318 145696 117374 145752
rect 117318 143248 117374 143304
rect 117318 140820 117374 140856
rect 117318 140800 117320 140820
rect 117320 140800 117372 140820
rect 117372 140800 117374 140820
rect 117686 138352 117742 138408
rect 117318 133592 117374 133648
rect 117502 116592 117558 116648
rect 117778 109248 117834 109304
rect 117318 102040 117374 102096
rect 117318 100816 117374 100872
rect 117226 92384 117282 92440
rect 117686 87488 117742 87544
rect 117870 85040 117926 85096
rect 117318 80144 117374 80200
rect 117686 77832 117742 77888
rect 117318 70488 117374 70544
rect 117318 68040 117374 68096
rect 117318 65592 117374 65648
rect 117870 63280 117926 63336
rect 117778 60832 117834 60888
rect 117318 58384 117374 58440
rect 117318 55936 117374 55992
rect 117318 53488 117374 53544
rect 117226 51040 117282 51096
rect 117318 48728 117374 48784
rect 117870 46280 117926 46336
rect 117226 43832 117282 43888
rect 117134 43696 117190 43752
rect 117318 41384 117374 41440
rect 117318 38936 117374 38992
rect 117318 36488 117374 36544
rect 117042 32272 117098 32328
rect 117318 31764 117320 31784
rect 117320 31764 117372 31784
rect 117372 31764 117374 31784
rect 117318 31728 117374 31764
rect 117318 29280 117374 29336
rect 117870 24384 117926 24440
rect 117778 21936 117834 21992
rect 117134 19624 117190 19680
rect 117502 17176 117558 17232
rect 117318 14728 117374 14784
rect 117226 12280 117282 12336
rect 117318 9832 117374 9888
rect 117318 7384 117374 7440
rect 117318 5072 117374 5128
rect 116950 3440 117006 3496
rect 118054 136040 118110 136096
rect 118054 126248 118110 126304
rect 118238 123800 118294 123856
rect 118330 119040 118386 119096
rect 118514 149912 118570 149968
rect 120078 154400 120134 154456
rect 119526 151952 119582 152008
rect 120630 155216 120686 155272
rect 118698 114144 118754 114200
rect 118606 104488 118662 104544
rect 118606 99592 118662 99648
rect 118514 75384 118570 75440
rect 118422 72936 118478 72992
rect 118422 34176 118478 34232
rect 118514 26832 118570 26888
rect 118422 6024 118478 6080
rect 118698 97144 118754 97200
rect 118790 94696 118846 94752
rect 118882 89936 118938 89992
rect 118606 3304 118662 3360
rect 121918 156576 121974 156632
rect 121458 155352 121514 155408
rect 121274 154672 121330 154728
rect 121458 154400 121514 154456
rect 121458 152496 121514 152552
rect 122286 155352 122342 155408
rect 123206 156576 123262 156632
rect 123206 154400 123262 154456
rect 127898 156032 127954 156088
rect 128082 152496 128138 152552
rect 131026 157120 131082 157176
rect 131118 154264 131174 154320
rect 136178 155488 136234 155544
rect 140870 155624 140926 155680
rect 142250 156168 142306 156224
rect 144918 152632 144974 152688
rect 146758 155216 146814 155272
rect 149150 155216 149206 155272
rect 149058 154536 149114 154592
rect 152462 157256 152518 157312
rect 153198 156712 153254 156768
rect 154578 155760 154634 155816
rect 161294 155216 161350 155272
rect 162858 156848 162914 156904
rect 170126 155896 170182 155952
rect 179602 156984 179658 157040
rect 179418 154808 179474 154864
rect 180430 155080 180486 155136
rect 186318 155352 186374 155408
rect 189078 152768 189134 152824
rect 190458 154944 190514 155000
rect 192114 152904 192170 152960
rect 200578 154672 200634 154728
rect 201866 156576 201922 156632
rect 204166 155352 204222 155408
rect 205178 152496 205234 152552
rect 207202 157120 207258 157176
rect 217782 155488 217838 155544
rect 221370 157256 221426 157312
rect 227258 155216 227314 155272
rect 231490 155624 231546 155680
rect 234342 155216 234398 155272
rect 251178 155352 251234 155408
rect 261666 155352 261722 155408
rect 262218 155488 262274 155544
rect 267554 155488 267610 155544
rect 271970 155624 272026 155680
rect 275926 155216 275982 155272
rect 277306 155080 277362 155136
rect 277398 154944 277454 155000
rect 292762 155352 292818 155408
rect 298190 155488 298246 155544
rect 494610 155896 494666 155952
rect 493966 155760 494022 155816
rect 497186 155624 497242 155680
rect 496542 155488 496598 155544
rect 499394 155352 499450 155408
rect 500866 155216 500922 155272
rect 506478 153176 506534 153232
rect 505650 151952 505706 152008
rect 510894 153312 510950 153368
rect 508870 153176 508926 153232
rect 512182 153448 512238 153504
rect 516690 153992 516746 154048
rect 516138 153856 516194 153912
rect 514758 153720 514814 153776
rect 513470 153584 513526 153640
rect 517978 154128 518034 154184
rect 519266 151816 519322 151872
rect 119526 2624 119582 2680
rect 119342 2352 119398 2408
rect 519726 148960 519782 149016
rect 119710 2488 119766 2544
rect 426346 3440 426402 3496
rect 520554 4664 520610 4720
rect 520646 4392 520702 4448
rect 522026 151000 522082 151056
rect 521842 150864 521898 150920
rect 521658 141752 521714 141808
rect 520830 121488 520886 121544
rect 520830 94560 520886 94616
rect 521750 108024 521806 108080
rect 521750 101360 521806 101416
rect 521658 7248 521714 7304
rect 521934 114824 521990 114880
rect 521934 87896 521990 87952
rect 521842 60968 521898 61024
rect 521658 4936 521714 4992
rect 522118 134952 522174 135008
rect 522210 128288 522266 128344
rect 522026 81232 522082 81288
rect 522026 74432 522082 74488
rect 522394 67768 522450 67824
rect 522118 47504 522174 47560
rect 522026 4800 522082 4856
rect 521934 4528 521990 4584
rect 522210 27376 522266 27432
rect 522578 34040 522634 34096
rect 522670 13912 522726 13968
rect 560942 155896 560998 155952
rect 559930 155760 559986 155816
rect 564806 155624 564862 155680
rect 563794 155488 563850 155544
rect 568670 155352 568726 155408
rect 570694 155216 570750 155272
rect 579434 152360 579490 152416
rect 550546 3304 550602 3360
<< metal3 >>
rect 0 157586 800 157616
rect 3141 157586 3207 157589
rect 0 157584 3207 157586
rect 0 157528 3146 157584
rect 3202 157528 3207 157584
rect 0 157526 3207 157528
rect 0 157496 800 157526
rect 3141 157523 3207 157526
rect 152457 157314 152523 157317
rect 221365 157314 221431 157317
rect 152457 157312 221431 157314
rect 152457 157256 152462 157312
rect 152518 157256 221370 157312
rect 221426 157256 221431 157312
rect 152457 157254 221431 157256
rect 152457 157251 152523 157254
rect 221365 157251 221431 157254
rect 131021 157178 131087 157181
rect 207197 157178 207263 157181
rect 131021 157176 207263 157178
rect 131021 157120 131026 157176
rect 131082 157120 207202 157176
rect 207258 157120 207263 157176
rect 131021 157118 207263 157120
rect 131021 157115 131087 157118
rect 207197 157115 207263 157118
rect 89161 157042 89227 157045
rect 179597 157042 179663 157045
rect 89161 157040 179663 157042
rect 89161 156984 89166 157040
rect 89222 156984 179602 157040
rect 179658 156984 179663 157040
rect 89161 156982 179663 156984
rect 89161 156979 89227 156982
rect 179597 156979 179663 156982
rect 64781 156906 64847 156909
rect 162853 156906 162919 156909
rect 64781 156904 162919 156906
rect 64781 156848 64786 156904
rect 64842 156848 162858 156904
rect 162914 156848 162919 156904
rect 64781 156846 162919 156848
rect 64781 156843 64847 156846
rect 162853 156843 162919 156846
rect 50153 156770 50219 156773
rect 153193 156770 153259 156773
rect 50153 156768 153259 156770
rect 50153 156712 50158 156768
rect 50214 156712 153198 156768
rect 153254 156712 153259 156768
rect 50153 156710 153259 156712
rect 50153 156707 50219 156710
rect 153193 156707 153259 156710
rect 3325 156634 3391 156637
rect 121913 156634 121979 156637
rect 3325 156632 121979 156634
rect 3325 156576 3330 156632
rect 3386 156576 121918 156632
rect 121974 156576 121979 156632
rect 3325 156574 121979 156576
rect 3325 156571 3391 156574
rect 121913 156571 121979 156574
rect 123201 156634 123267 156637
rect 201861 156634 201927 156637
rect 123201 156632 201927 156634
rect 123201 156576 123206 156632
rect 123262 156576 201866 156632
rect 201922 156576 201927 156632
rect 123201 156574 201927 156576
rect 123201 156571 123267 156574
rect 201861 156571 201927 156574
rect 34697 156226 34763 156229
rect 142245 156226 142311 156229
rect 34697 156224 142311 156226
rect 34697 156168 34702 156224
rect 34758 156168 142250 156224
rect 142306 156168 142311 156224
rect 34697 156166 142311 156168
rect 34697 156163 34763 156166
rect 142245 156163 142311 156166
rect 17861 156090 17927 156093
rect 127893 156090 127959 156093
rect 17861 156088 127959 156090
rect 17861 156032 17866 156088
rect 17922 156032 127898 156088
rect 127954 156032 127959 156088
rect 17861 156030 127959 156032
rect 17861 156027 17927 156030
rect 127893 156027 127959 156030
rect 75453 155954 75519 155957
rect 170121 155954 170187 155957
rect 75453 155952 170187 155954
rect 75453 155896 75458 155952
rect 75514 155896 170126 155952
rect 170182 155896 170187 155952
rect 75453 155894 170187 155896
rect 75453 155891 75519 155894
rect 170121 155891 170187 155894
rect 494605 155954 494671 155957
rect 560937 155954 561003 155957
rect 494605 155952 561003 155954
rect 494605 155896 494610 155952
rect 494666 155896 560942 155952
rect 560998 155896 561003 155952
rect 494605 155894 561003 155896
rect 494605 155891 494671 155894
rect 560937 155891 561003 155894
rect 52085 155818 52151 155821
rect 154573 155818 154639 155821
rect 52085 155816 154639 155818
rect 52085 155760 52090 155816
rect 52146 155760 154578 155816
rect 154634 155760 154639 155816
rect 52085 155758 154639 155760
rect 52085 155755 52151 155758
rect 154573 155755 154639 155758
rect 493961 155818 494027 155821
rect 559925 155818 559991 155821
rect 493961 155816 559991 155818
rect 493961 155760 493966 155816
rect 494022 155760 559930 155816
rect 559986 155760 559991 155816
rect 493961 155758 559991 155760
rect 493961 155755 494027 155758
rect 559925 155755 559991 155758
rect 36537 155682 36603 155685
rect 140865 155682 140931 155685
rect 36537 155680 140931 155682
rect 36537 155624 36542 155680
rect 36598 155624 140870 155680
rect 140926 155624 140931 155680
rect 36537 155622 140931 155624
rect 36537 155619 36603 155622
rect 140865 155619 140931 155622
rect 231485 155682 231551 155685
rect 271965 155682 272031 155685
rect 231485 155680 272031 155682
rect 231485 155624 231490 155680
rect 231546 155624 271970 155680
rect 272026 155624 272031 155680
rect 231485 155622 272031 155624
rect 231485 155619 231551 155622
rect 271965 155619 272031 155622
rect 497181 155682 497247 155685
rect 564801 155682 564867 155685
rect 497181 155680 564867 155682
rect 497181 155624 497186 155680
rect 497242 155624 564806 155680
rect 564862 155624 564867 155680
rect 497181 155622 564867 155624
rect 497181 155619 497247 155622
rect 564801 155619 564867 155622
rect 24761 155546 24827 155549
rect 136173 155546 136239 155549
rect 24761 155544 136239 155546
rect 24761 155488 24766 155544
rect 24822 155488 136178 155544
rect 136234 155488 136239 155544
rect 24761 155486 136239 155488
rect 24761 155483 24827 155486
rect 136173 155483 136239 155486
rect 217777 155546 217843 155549
rect 262213 155546 262279 155549
rect 217777 155544 262279 155546
rect 217777 155488 217782 155544
rect 217838 155488 262218 155544
rect 262274 155488 262279 155544
rect 217777 155486 262279 155488
rect 217777 155483 217843 155486
rect 262213 155483 262279 155486
rect 267549 155546 267615 155549
rect 298185 155546 298251 155549
rect 267549 155544 298251 155546
rect 267549 155488 267554 155544
rect 267610 155488 298190 155544
rect 298246 155488 298251 155544
rect 267549 155486 298251 155488
rect 267549 155483 267615 155486
rect 298185 155483 298251 155486
rect 496537 155546 496603 155549
rect 563789 155546 563855 155549
rect 496537 155544 563855 155546
rect 496537 155488 496542 155544
rect 496598 155488 563794 155544
rect 563850 155488 563855 155544
rect 496537 155486 563855 155488
rect 496537 155483 496603 155486
rect 563789 155483 563855 155486
rect 5257 155410 5323 155413
rect 121453 155410 121519 155413
rect 5257 155408 121519 155410
rect 5257 155352 5262 155408
rect 5318 155352 121458 155408
rect 121514 155352 121519 155408
rect 5257 155350 121519 155352
rect 5257 155347 5323 155350
rect 121453 155347 121519 155350
rect 122281 155410 122347 155413
rect 186313 155410 186379 155413
rect 122281 155408 186379 155410
rect 122281 155352 122286 155408
rect 122342 155352 186318 155408
rect 186374 155352 186379 155408
rect 122281 155350 186379 155352
rect 122281 155347 122347 155350
rect 186313 155347 186379 155350
rect 204161 155410 204227 155413
rect 251173 155410 251239 155413
rect 204161 155408 251239 155410
rect 204161 155352 204166 155408
rect 204222 155352 251178 155408
rect 251234 155352 251239 155408
rect 204161 155350 251239 155352
rect 204161 155347 204227 155350
rect 251173 155347 251239 155350
rect 261661 155410 261727 155413
rect 292757 155410 292823 155413
rect 261661 155408 292823 155410
rect 261661 155352 261666 155408
rect 261722 155352 292762 155408
rect 292818 155352 292823 155408
rect 261661 155350 292823 155352
rect 261661 155347 261727 155350
rect 292757 155347 292823 155350
rect 499389 155410 499455 155413
rect 568665 155410 568731 155413
rect 499389 155408 568731 155410
rect 499389 155352 499394 155408
rect 499450 155352 568670 155408
rect 568726 155352 568731 155408
rect 499389 155350 568731 155352
rect 499389 155347 499455 155350
rect 568665 155347 568731 155350
rect 1393 155274 1459 155277
rect 120625 155274 120691 155277
rect 1393 155272 120691 155274
rect 1393 155216 1398 155272
rect 1454 155216 120630 155272
rect 120686 155216 120691 155272
rect 1393 155214 120691 155216
rect 1393 155211 1459 155214
rect 120625 155211 120691 155214
rect 146753 155274 146819 155277
rect 149145 155274 149211 155277
rect 146753 155272 149211 155274
rect 146753 155216 146758 155272
rect 146814 155216 149150 155272
rect 149206 155216 149211 155272
rect 146753 155214 149211 155216
rect 146753 155211 146819 155214
rect 149145 155211 149211 155214
rect 161289 155274 161355 155277
rect 227253 155274 227319 155277
rect 161289 155272 227319 155274
rect 161289 155216 161294 155272
rect 161350 155216 227258 155272
rect 227314 155216 227319 155272
rect 161289 155214 227319 155216
rect 161289 155211 161355 155214
rect 227253 155211 227319 155214
rect 234337 155274 234403 155277
rect 275921 155274 275987 155277
rect 234337 155272 275987 155274
rect 234337 155216 234342 155272
rect 234398 155216 275926 155272
rect 275982 155216 275987 155272
rect 234337 155214 275987 155216
rect 234337 155211 234403 155214
rect 275921 155211 275987 155214
rect 500861 155274 500927 155277
rect 570689 155274 570755 155277
rect 500861 155272 570755 155274
rect 500861 155216 500866 155272
rect 500922 155216 570694 155272
rect 570750 155216 570755 155272
rect 500861 155214 570755 155216
rect 500861 155211 500927 155214
rect 570689 155211 570755 155214
rect 91093 155138 91159 155141
rect 180425 155138 180491 155141
rect 91093 155136 180491 155138
rect 91093 155080 91098 155136
rect 91154 155080 180430 155136
rect 180486 155080 180491 155136
rect 91093 155078 180491 155080
rect 91093 155075 91159 155078
rect 180425 155075 180491 155078
rect 277301 155138 277367 155141
rect 277301 155136 277410 155138
rect 277301 155080 277306 155136
rect 277362 155080 277410 155136
rect 277301 155075 277410 155080
rect 277350 155005 277410 155075
rect 105721 155002 105787 155005
rect 190453 155002 190519 155005
rect 105721 155000 190519 155002
rect 105721 154944 105726 155000
rect 105782 154944 190458 155000
rect 190514 154944 190519 155000
rect 105721 154942 190519 154944
rect 277350 155000 277459 155005
rect 277350 154944 277398 155000
rect 277454 154944 277459 155000
rect 277350 154942 277459 154944
rect 105721 154939 105787 154942
rect 190453 154939 190519 154942
rect 277393 154939 277459 154942
rect 97901 154866 97967 154869
rect 179413 154866 179479 154869
rect 97901 154864 179479 154866
rect 97901 154808 97906 154864
rect 97962 154808 179418 154864
rect 179474 154808 179479 154864
rect 97901 154806 179479 154808
rect 97901 154803 97967 154806
rect 179413 154803 179479 154806
rect 121269 154730 121335 154733
rect 200573 154730 200639 154733
rect 121269 154728 200639 154730
rect 121269 154672 121274 154728
rect 121330 154672 200578 154728
rect 200634 154672 200639 154728
rect 121269 154670 200639 154672
rect 121269 154667 121335 154670
rect 200573 154667 200639 154670
rect 70577 154594 70643 154597
rect 149053 154594 149119 154597
rect 70577 154592 149119 154594
rect 70577 154536 70582 154592
rect 70638 154536 149058 154592
rect 149114 154536 149119 154592
rect 70577 154534 149119 154536
rect 70577 154531 70643 154534
rect 149053 154531 149119 154534
rect 106181 154458 106247 154461
rect 120073 154458 120139 154461
rect 106181 154456 120139 154458
rect 106181 154400 106186 154456
rect 106242 154400 120078 154456
rect 120134 154400 120139 154456
rect 106181 154398 120139 154400
rect 106181 154395 106247 154398
rect 120073 154395 120139 154398
rect 121453 154458 121519 154461
rect 123201 154458 123267 154461
rect 121453 154456 123267 154458
rect 121453 154400 121458 154456
rect 121514 154400 123206 154456
rect 123262 154400 123267 154456
rect 121453 154398 123267 154400
rect 121453 154395 121519 154398
rect 123201 154395 123267 154398
rect 17033 154322 17099 154325
rect 131113 154322 131179 154325
rect 17033 154320 131179 154322
rect 17033 154264 17038 154320
rect 17094 154264 131118 154320
rect 131174 154264 131179 154320
rect 17033 154262 131179 154264
rect 17033 154259 17099 154262
rect 131113 154259 131179 154262
rect 91921 154186 91987 154189
rect 517973 154186 518039 154189
rect 91921 154184 518039 154186
rect 91921 154128 91926 154184
rect 91982 154128 517978 154184
rect 518034 154128 518039 154184
rect 91921 154126 518039 154128
rect 91921 154123 91987 154126
rect 517973 154123 518039 154126
rect 88057 154050 88123 154053
rect 516685 154050 516751 154053
rect 88057 154048 516751 154050
rect 88057 153992 88062 154048
rect 88118 153992 516690 154048
rect 516746 153992 516751 154048
rect 88057 153990 516751 153992
rect 88057 153987 88123 153990
rect 516685 153987 516751 153990
rect 81157 153914 81223 153917
rect 516133 153914 516199 153917
rect 81157 153912 516199 153914
rect 81157 153856 81162 153912
rect 81218 153856 516138 153912
rect 516194 153856 516199 153912
rect 81157 153854 516199 153856
rect 81157 153851 81223 153854
rect 516133 153851 516199 153854
rect 50613 153778 50679 153781
rect 514753 153778 514819 153781
rect 50613 153776 514819 153778
rect 50613 153720 50618 153776
rect 50674 153720 514758 153776
rect 514814 153720 514819 153776
rect 50613 153718 514819 153720
rect 50613 153715 50679 153718
rect 514753 153715 514819 153718
rect 39849 153642 39915 153645
rect 513465 153642 513531 153645
rect 39849 153640 513531 153642
rect 39849 153584 39854 153640
rect 39910 153584 513470 153640
rect 513526 153584 513531 153640
rect 39849 153582 513531 153584
rect 39849 153579 39915 153582
rect 513465 153579 513531 153582
rect 30005 153506 30071 153509
rect 512177 153506 512243 153509
rect 30005 153504 512243 153506
rect 30005 153448 30010 153504
rect 30066 153448 512182 153504
rect 512238 153448 512243 153504
rect 30005 153446 512243 153448
rect 30005 153443 30071 153446
rect 512177 153443 512243 153446
rect 9397 153372 9463 153373
rect 9397 153370 9444 153372
rect 9352 153368 9444 153370
rect 9352 153312 9402 153368
rect 9352 153310 9444 153312
rect 9397 153308 9444 153310
rect 9508 153308 9514 153372
rect 26601 153370 26667 153373
rect 510889 153370 510955 153373
rect 26601 153368 510955 153370
rect 26601 153312 26606 153368
rect 26662 153312 510894 153368
rect 510950 153312 510955 153368
rect 26601 153310 510955 153312
rect 9397 153307 9463 153308
rect 26601 153307 26667 153310
rect 510889 153307 510955 153310
rect 19701 153234 19767 153237
rect 506473 153236 506539 153237
rect 19701 153232 506306 153234
rect 19701 153176 19706 153232
rect 19762 153176 506306 153232
rect 19701 153174 506306 153176
rect 19701 153171 19767 153174
rect 506246 153098 506306 153174
rect 506422 153172 506428 153236
rect 506492 153234 506539 153236
rect 508865 153234 508931 153237
rect 506492 153232 506584 153234
rect 506534 153176 506584 153232
rect 506492 153174 506584 153176
rect 506798 153232 508931 153234
rect 506798 153176 508870 153232
rect 508926 153176 508931 153232
rect 506798 153174 508931 153176
rect 506492 153172 506539 153174
rect 506473 153171 506539 153172
rect 506798 153098 506858 153174
rect 508865 153171 508931 153174
rect 506246 153038 506858 153098
rect 0 152962 800 152992
rect 3233 152962 3299 152965
rect 0 152960 3299 152962
rect 0 152904 3238 152960
rect 3294 152904 3299 152960
rect 0 152902 3299 152904
rect 0 152872 800 152902
rect 3233 152899 3299 152902
rect 108665 152962 108731 152965
rect 192109 152962 192175 152965
rect 108665 152960 192175 152962
rect 108665 152904 108670 152960
rect 108726 152904 192114 152960
rect 192170 152904 192175 152960
rect 108665 152902 192175 152904
rect 108665 152899 108731 152902
rect 192109 152899 192175 152902
rect 103789 152826 103855 152829
rect 189073 152826 189139 152829
rect 103789 152824 189139 152826
rect 103789 152768 103794 152824
rect 103850 152768 189078 152824
rect 189134 152768 189139 152824
rect 103789 152766 189139 152768
rect 103789 152763 103855 152766
rect 189073 152763 189139 152766
rect 37457 152690 37523 152693
rect 144913 152690 144979 152693
rect 37457 152688 144979 152690
rect 37457 152632 37462 152688
rect 37518 152632 144918 152688
rect 144974 152632 144979 152688
rect 37457 152630 144979 152632
rect 37457 152627 37523 152630
rect 144913 152627 144979 152630
rect 2405 152554 2471 152557
rect 121453 152554 121519 152557
rect 2405 152552 121519 152554
rect 2405 152496 2410 152552
rect 2466 152496 121458 152552
rect 121514 152496 121519 152552
rect 2405 152494 121519 152496
rect 2405 152491 2471 152494
rect 121453 152491 121519 152494
rect 128077 152554 128143 152557
rect 205173 152554 205239 152557
rect 128077 152552 205239 152554
rect 128077 152496 128082 152552
rect 128138 152496 205178 152552
rect 205234 152496 205239 152552
rect 128077 152494 205239 152496
rect 128077 152491 128143 152494
rect 205173 152491 205239 152494
rect 3141 152418 3207 152421
rect 115749 152418 115815 152421
rect 3141 152416 115815 152418
rect 3141 152360 3146 152416
rect 3202 152360 115754 152416
rect 115810 152360 115815 152416
rect 3141 152358 115815 152360
rect 3141 152355 3207 152358
rect 115749 152355 115815 152358
rect 118693 152418 118759 152421
rect 579429 152418 579495 152421
rect 118693 152416 579495 152418
rect 118693 152360 118698 152416
rect 118754 152360 579434 152416
rect 579490 152360 579495 152416
rect 118693 152358 579495 152360
rect 118693 152355 118759 152358
rect 579429 152355 579495 152358
rect 119521 152010 119587 152013
rect 505645 152010 505711 152013
rect 119521 152008 505711 152010
rect 119521 151952 119526 152008
rect 119582 151952 505650 152008
rect 505706 151952 505711 152008
rect 119521 151950 505711 151952
rect 119521 151947 119587 151950
rect 505645 151947 505711 151950
rect 102041 151874 102107 151877
rect 519261 151874 519327 151877
rect 102041 151872 519327 151874
rect 102041 151816 102046 151872
rect 102102 151816 519266 151872
rect 519322 151816 519327 151872
rect 102041 151814 519327 151816
rect 102041 151811 102107 151814
rect 519261 151811 519327 151814
rect 26190 151542 45570 151602
rect 23105 151330 23171 151333
rect 26190 151330 26250 151542
rect 33501 151466 33567 151469
rect 33501 151464 41338 151466
rect 33501 151408 33506 151464
rect 33562 151408 41338 151464
rect 33501 151406 41338 151408
rect 33501 151403 33567 151406
rect 23105 151328 26250 151330
rect 23105 151272 23110 151328
rect 23166 151272 26250 151328
rect 23105 151270 26250 151272
rect 36905 151330 36971 151333
rect 36905 151328 41154 151330
rect 36905 151272 36910 151328
rect 36966 151272 41154 151328
rect 36905 151270 41154 151272
rect 23105 151267 23171 151270
rect 36905 151267 36971 151270
rect 41094 150650 41154 151270
rect 41278 151194 41338 151406
rect 45510 151330 45570 151542
rect 51030 151542 60750 151602
rect 51030 151330 51090 151542
rect 45510 151270 51090 151330
rect 53054 151406 57990 151466
rect 41278 151134 45570 151194
rect 45510 150922 45570 151134
rect 53054 150922 53114 151406
rect 53925 151328 53991 151333
rect 53925 151272 53930 151328
rect 53986 151272 53991 151328
rect 53925 151267 53991 151272
rect 53928 151058 53988 151267
rect 57930 151058 57990 151406
rect 60690 151330 60750 151542
rect 70350 151542 92674 151602
rect 70350 151330 70410 151542
rect 92062 151406 92490 151466
rect 60690 151270 70410 151330
rect 71313 151330 71379 151333
rect 71313 151328 75378 151330
rect 71313 151272 71318 151328
rect 71374 151272 75378 151328
rect 71313 151270 75378 151272
rect 71313 151267 71379 151270
rect 75318 151194 75378 151270
rect 92062 151194 92122 151406
rect 92197 151330 92263 151333
rect 92197 151328 92306 151330
rect 92197 151272 92202 151328
rect 92258 151272 92306 151328
rect 92197 151267 92306 151272
rect 75318 151134 92122 151194
rect 92246 151058 92306 151267
rect 92430 151194 92490 151406
rect 92614 151330 92674 151542
rect 98821 151466 98887 151469
rect 112437 151466 112503 151469
rect 98821 151464 112503 151466
rect 98821 151408 98826 151464
rect 98882 151408 112442 151464
rect 112498 151408 112503 151464
rect 98821 151406 112503 151408
rect 98821 151403 98887 151406
rect 112437 151403 112503 151406
rect 118141 151330 118207 151333
rect 92614 151328 118207 151330
rect 92614 151272 118146 151328
rect 118202 151272 118207 151328
rect 92614 151270 118207 151272
rect 118141 151267 118207 151270
rect 116577 151194 116643 151197
rect 92430 151192 116643 151194
rect 92430 151136 116582 151192
rect 116638 151136 116643 151192
rect 92430 151134 116643 151136
rect 116577 151131 116643 151134
rect 522021 151058 522087 151061
rect 53928 150998 55874 151058
rect 57930 150998 60750 151058
rect 92246 151056 522087 151058
rect 92246 151000 522026 151056
rect 522082 151000 522087 151056
rect 92246 150998 522087 151000
rect 45510 150862 53114 150922
rect 55814 150786 55874 150998
rect 60690 150922 60750 150998
rect 522021 150995 522087 150998
rect 521837 150922 521903 150925
rect 60690 150920 521903 150922
rect 60690 150864 521842 150920
rect 521898 150864 521903 150920
rect 60690 150862 521903 150864
rect 521837 150859 521903 150862
rect 117957 150786 118023 150789
rect 55814 150784 118023 150786
rect 55814 150728 117962 150784
rect 118018 150728 118023 150784
rect 55814 150726 118023 150728
rect 117957 150723 118023 150726
rect 113817 150650 113883 150653
rect 41094 150648 113883 150650
rect 41094 150592 113822 150648
rect 113878 150592 113883 150648
rect 41094 150590 113883 150592
rect 113817 150587 113883 150590
rect 117773 150650 117839 150653
rect 117773 150648 120060 150650
rect 117773 150592 117778 150648
rect 117834 150592 120060 150648
rect 117773 150590 120060 150592
rect 117773 150587 117839 150590
rect 112437 150514 112503 150517
rect 115197 150514 115263 150517
rect 112437 150512 115263 150514
rect 112437 150456 112442 150512
rect 112498 150456 115202 150512
rect 115258 150456 115263 150512
rect 112437 150454 115263 150456
rect 112437 150451 112503 150454
rect 115197 150451 115263 150454
rect 3325 149970 3391 149973
rect 118509 149970 118575 149973
rect 3325 149968 118575 149970
rect 3325 149912 3330 149968
rect 3386 149912 118514 149968
rect 118570 149912 118575 149968
rect 3325 149910 118575 149912
rect 3325 149907 3391 149910
rect 118509 149907 118575 149910
rect 519721 149018 519787 149021
rect 519678 149016 519787 149018
rect 519678 148960 519726 149016
rect 519782 148960 519787 149016
rect 519678 148955 519787 148960
rect 0 148474 800 148504
rect 3509 148474 3575 148477
rect 0 148472 3575 148474
rect 0 148416 3514 148472
rect 3570 148416 3575 148472
rect 519678 148444 519738 148955
rect 0 148414 3575 148416
rect 0 148384 800 148414
rect 3509 148411 3575 148414
rect 117681 148202 117747 148205
rect 117681 148200 120060 148202
rect 117681 148144 117686 148200
rect 117742 148144 120060 148200
rect 117681 148142 120060 148144
rect 117681 148139 117747 148142
rect 117221 146162 117287 146165
rect 113804 146160 117287 146162
rect 113804 146104 117226 146160
rect 117282 146104 117287 146160
rect 113804 146102 117287 146104
rect 117221 146099 117287 146102
rect 117313 145754 117379 145757
rect 117313 145752 120060 145754
rect 117313 145696 117318 145752
rect 117374 145696 120060 145752
rect 117313 145694 120060 145696
rect 117313 145691 117379 145694
rect 0 143850 800 143880
rect 2957 143850 3023 143853
rect 0 143848 3023 143850
rect 0 143792 2962 143848
rect 3018 143792 3023 143848
rect 0 143790 3023 143792
rect 0 143760 800 143790
rect 2957 143787 3023 143790
rect 117313 143306 117379 143309
rect 117313 143304 120060 143306
rect 117313 143248 117318 143304
rect 117374 143248 120060 143304
rect 117313 143246 120060 143248
rect 117313 143243 117379 143246
rect 521653 141810 521719 141813
rect 519892 141808 521719 141810
rect 519892 141752 521658 141808
rect 521714 141752 521719 141808
rect 519892 141750 521719 141752
rect 521653 141747 521719 141750
rect 117313 140858 117379 140861
rect 117313 140856 120060 140858
rect 117313 140800 117318 140856
rect 117374 140800 120060 140856
rect 117313 140798 120060 140800
rect 117313 140795 117379 140798
rect 0 139362 800 139392
rect 3233 139362 3299 139365
rect 0 139360 3299 139362
rect 0 139304 3238 139360
rect 3294 139304 3299 139360
rect 0 139302 3299 139304
rect 0 139272 800 139302
rect 3233 139299 3299 139302
rect 117681 138410 117747 138413
rect 117681 138408 120060 138410
rect 117681 138352 117686 138408
rect 117742 138352 120060 138408
rect 117681 138350 120060 138352
rect 117681 138347 117747 138350
rect 118049 136098 118115 136101
rect 118049 136096 120060 136098
rect 118049 136040 118054 136096
rect 118110 136040 120060 136096
rect 118049 136038 120060 136040
rect 118049 136035 118115 136038
rect 522113 135010 522179 135013
rect 519892 135008 522179 135010
rect 519892 134952 522118 135008
rect 522174 134952 522179 135008
rect 519892 134950 522179 134952
rect 522113 134947 522179 134950
rect 0 134738 800 134768
rect 3325 134738 3391 134741
rect 116669 134738 116735 134741
rect 0 134736 3391 134738
rect 0 134680 3330 134736
rect 3386 134680 3391 134736
rect 0 134678 3391 134680
rect 113804 134736 116735 134738
rect 113804 134680 116674 134736
rect 116730 134680 116735 134736
rect 113804 134678 116735 134680
rect 0 134648 800 134678
rect 3325 134675 3391 134678
rect 116669 134675 116735 134678
rect 117313 133650 117379 133653
rect 117313 133648 120060 133650
rect 117313 133592 117318 133648
rect 117374 133592 120060 133648
rect 117313 133590 120060 133592
rect 117313 133587 117379 133590
rect 116761 131202 116827 131205
rect 116761 131200 120060 131202
rect 116761 131144 116766 131200
rect 116822 131144 120060 131200
rect 116761 131142 120060 131144
rect 116761 131139 116827 131142
rect 0 130114 800 130144
rect 3969 130114 4035 130117
rect 0 130112 4035 130114
rect 0 130056 3974 130112
rect 4030 130056 4035 130112
rect 0 130054 4035 130056
rect 0 130024 800 130054
rect 3969 130051 4035 130054
rect 117129 128754 117195 128757
rect 117129 128752 120060 128754
rect 117129 128696 117134 128752
rect 117190 128696 120060 128752
rect 117129 128694 120060 128696
rect 117129 128691 117195 128694
rect 522205 128346 522271 128349
rect 519892 128344 522271 128346
rect 519892 128288 522210 128344
rect 522266 128288 522271 128344
rect 519892 128286 522271 128288
rect 522205 128283 522271 128286
rect 118049 126306 118115 126309
rect 118049 126304 120060 126306
rect 118049 126248 118054 126304
rect 118110 126248 120060 126304
rect 118049 126246 120060 126248
rect 118049 126243 118115 126246
rect 0 125626 800 125656
rect 3877 125626 3943 125629
rect 0 125624 3943 125626
rect 0 125568 3882 125624
rect 3938 125568 3943 125624
rect 0 125566 3943 125568
rect 0 125536 800 125566
rect 3877 125563 3943 125566
rect 118233 123858 118299 123861
rect 118233 123856 120060 123858
rect 118233 123800 118238 123856
rect 118294 123800 120060 123856
rect 118233 123798 120060 123800
rect 118233 123795 118299 123798
rect 116945 123314 117011 123317
rect 113804 123312 117011 123314
rect 113804 123256 116950 123312
rect 117006 123256 117011 123312
rect 113804 123254 117011 123256
rect 116945 123251 117011 123254
rect 116853 121546 116919 121549
rect 520825 121546 520891 121549
rect 116853 121544 120060 121546
rect 116853 121488 116858 121544
rect 116914 121488 120060 121544
rect 116853 121486 120060 121488
rect 519892 121544 520891 121546
rect 519892 121488 520830 121544
rect 520886 121488 520891 121544
rect 519892 121486 520891 121488
rect 116853 121483 116919 121486
rect 520825 121483 520891 121486
rect 0 121002 800 121032
rect 3785 121002 3851 121005
rect 0 121000 3851 121002
rect 0 120944 3790 121000
rect 3846 120944 3851 121000
rect 0 120942 3851 120944
rect 0 120912 800 120942
rect 3785 120939 3851 120942
rect 118325 119098 118391 119101
rect 118325 119096 120060 119098
rect 118325 119040 118330 119096
rect 118386 119040 120060 119096
rect 118325 119038 120060 119040
rect 118325 119035 118391 119038
rect 117497 116650 117563 116653
rect 117497 116648 120060 116650
rect 117497 116592 117502 116648
rect 117558 116592 120060 116648
rect 117497 116590 120060 116592
rect 117497 116587 117563 116590
rect 0 116514 800 116544
rect 3693 116514 3759 116517
rect 0 116512 3759 116514
rect 0 116456 3698 116512
rect 3754 116456 3759 116512
rect 0 116454 3759 116456
rect 0 116424 800 116454
rect 3693 116451 3759 116454
rect 521929 114882 521995 114885
rect 519892 114880 521995 114882
rect 519892 114824 521934 114880
rect 521990 114824 521995 114880
rect 519892 114822 521995 114824
rect 521929 114819 521995 114822
rect 118693 114202 118759 114205
rect 118693 114200 120060 114202
rect 118693 114144 118698 114200
rect 118754 114144 120060 114200
rect 118693 114142 120060 114144
rect 118693 114139 118759 114142
rect 116853 112026 116919 112029
rect 113804 112024 116919 112026
rect 113804 111968 116858 112024
rect 116914 111968 116919 112024
rect 113804 111966 116919 111968
rect 116853 111963 116919 111966
rect 0 111890 800 111920
rect 3601 111890 3667 111893
rect 0 111888 3667 111890
rect 0 111832 3606 111888
rect 3662 111832 3667 111888
rect 0 111830 3667 111832
rect 0 111800 800 111830
rect 3601 111827 3667 111830
rect 116945 111754 117011 111757
rect 116945 111752 120060 111754
rect 116945 111696 116950 111752
rect 117006 111696 120060 111752
rect 116945 111694 120060 111696
rect 116945 111691 117011 111694
rect 117773 109306 117839 109309
rect 117773 109304 120060 109306
rect 117773 109248 117778 109304
rect 117834 109248 120060 109304
rect 117773 109246 120060 109248
rect 117773 109243 117839 109246
rect 521745 108082 521811 108085
rect 519892 108080 521811 108082
rect 519892 108024 521750 108080
rect 521806 108024 521811 108080
rect 519892 108022 521811 108024
rect 521745 108019 521811 108022
rect 0 107266 800 107296
rect 3509 107266 3575 107269
rect 0 107264 3575 107266
rect 0 107208 3514 107264
rect 3570 107208 3575 107264
rect 0 107206 3575 107208
rect 0 107176 800 107206
rect 3509 107203 3575 107206
rect 117129 106994 117195 106997
rect 117129 106992 120060 106994
rect 117129 106936 117134 106992
rect 117190 106936 120060 106992
rect 117129 106934 120060 106936
rect 117129 106931 117195 106934
rect 118601 104546 118667 104549
rect 118601 104544 120060 104546
rect 118601 104488 118606 104544
rect 118662 104488 120060 104544
rect 118601 104486 120060 104488
rect 118601 104483 118667 104486
rect 0 102778 800 102808
rect 3417 102778 3483 102781
rect 0 102776 3483 102778
rect 0 102720 3422 102776
rect 3478 102720 3483 102776
rect 0 102718 3483 102720
rect 0 102688 800 102718
rect 3417 102715 3483 102718
rect 117313 102098 117379 102101
rect 117313 102096 120060 102098
rect 117313 102040 117318 102096
rect 117374 102040 120060 102096
rect 117313 102038 120060 102040
rect 117313 102035 117379 102038
rect 521745 101418 521811 101421
rect 519892 101416 521811 101418
rect 519892 101360 521750 101416
rect 521806 101360 521811 101416
rect 519892 101358 521811 101360
rect 521745 101355 521811 101358
rect 117313 100874 117379 100877
rect 117270 100872 117379 100874
rect 117270 100816 117318 100872
rect 117374 100816 117379 100872
rect 117270 100811 117379 100816
rect 117270 100738 117330 100811
rect 113774 100678 117330 100738
rect 113774 100572 113834 100678
rect 118601 99650 118667 99653
rect 118601 99648 120060 99650
rect 118601 99592 118606 99648
rect 118662 99592 120060 99648
rect 118601 99590 120060 99592
rect 118601 99587 118667 99590
rect 0 98154 800 98184
rect 3785 98154 3851 98157
rect 0 98152 3851 98154
rect 0 98096 3790 98152
rect 3846 98096 3851 98152
rect 0 98094 3851 98096
rect 0 98064 800 98094
rect 3785 98091 3851 98094
rect 118693 97202 118759 97205
rect 118693 97200 120060 97202
rect 118693 97144 118698 97200
rect 118754 97144 120060 97200
rect 118693 97142 120060 97144
rect 118693 97139 118759 97142
rect 118785 94754 118851 94757
rect 118785 94752 120060 94754
rect 118785 94696 118790 94752
rect 118846 94696 120060 94752
rect 118785 94694 120060 94696
rect 118785 94691 118851 94694
rect 520825 94618 520891 94621
rect 519892 94616 520891 94618
rect 519892 94560 520830 94616
rect 520886 94560 520891 94616
rect 519892 94558 520891 94560
rect 520825 94555 520891 94558
rect 0 93666 800 93696
rect 3417 93666 3483 93669
rect 0 93664 3483 93666
rect 0 93608 3422 93664
rect 3478 93608 3483 93664
rect 0 93606 3483 93608
rect 0 93576 800 93606
rect 3417 93603 3483 93606
rect 117221 92442 117287 92445
rect 117221 92440 120060 92442
rect 117221 92384 117226 92440
rect 117282 92384 120060 92440
rect 117221 92382 120060 92384
rect 117221 92379 117287 92382
rect 118877 89994 118943 89997
rect 118877 89992 120060 89994
rect 118877 89936 118882 89992
rect 118938 89936 120060 89992
rect 118877 89934 120060 89936
rect 118877 89931 118943 89934
rect 116485 89178 116551 89181
rect 113804 89176 116551 89178
rect 113804 89120 116490 89176
rect 116546 89120 116551 89176
rect 113804 89118 116551 89120
rect 116485 89115 116551 89118
rect 0 89042 800 89072
rect 3693 89042 3759 89045
rect 0 89040 3759 89042
rect 0 88984 3698 89040
rect 3754 88984 3759 89040
rect 0 88982 3759 88984
rect 0 88952 800 88982
rect 3693 88979 3759 88982
rect 521929 87954 521995 87957
rect 519892 87952 521995 87954
rect 519892 87896 521934 87952
rect 521990 87896 521995 87952
rect 519892 87894 521995 87896
rect 521929 87891 521995 87894
rect 117681 87546 117747 87549
rect 117681 87544 120060 87546
rect 117681 87488 117686 87544
rect 117742 87488 120060 87544
rect 117681 87486 120060 87488
rect 117681 87483 117747 87486
rect 117865 85098 117931 85101
rect 117865 85096 120060 85098
rect 117865 85040 117870 85096
rect 117926 85040 120060 85096
rect 117865 85038 120060 85040
rect 117865 85035 117931 85038
rect 0 84418 800 84448
rect 3601 84418 3667 84421
rect 0 84416 3667 84418
rect 0 84360 3606 84416
rect 3662 84360 3667 84416
rect 0 84358 3667 84360
rect 0 84328 800 84358
rect 3601 84355 3667 84358
rect 117037 82650 117103 82653
rect 117037 82648 120060 82650
rect 117037 82592 117042 82648
rect 117098 82592 120060 82648
rect 117037 82590 120060 82592
rect 117037 82587 117103 82590
rect 522021 81290 522087 81293
rect 519892 81288 522087 81290
rect 519892 81232 522026 81288
rect 522082 81232 522087 81288
rect 519892 81230 522087 81232
rect 522021 81227 522087 81230
rect 117313 80202 117379 80205
rect 117313 80200 120060 80202
rect 117313 80144 117318 80200
rect 117374 80144 120060 80200
rect 117313 80142 120060 80144
rect 117313 80139 117379 80142
rect 0 79930 800 79960
rect 3877 79930 3943 79933
rect 0 79928 3943 79930
rect 0 79872 3882 79928
rect 3938 79872 3943 79928
rect 0 79870 3943 79872
rect 0 79840 800 79870
rect 3877 79867 3943 79870
rect 117446 77890 117452 77892
rect 113804 77830 117452 77890
rect 117446 77828 117452 77830
rect 117516 77828 117522 77892
rect 117681 77890 117747 77893
rect 117681 77888 120060 77890
rect 117681 77832 117686 77888
rect 117742 77832 120060 77888
rect 117681 77830 120060 77832
rect 117681 77827 117747 77830
rect 118509 75442 118575 75445
rect 118509 75440 120060 75442
rect 118509 75384 118514 75440
rect 118570 75384 120060 75440
rect 118509 75382 120060 75384
rect 118509 75379 118575 75382
rect 0 75306 800 75336
rect 3509 75306 3575 75309
rect 0 75304 3575 75306
rect 0 75248 3514 75304
rect 3570 75248 3575 75304
rect 0 75246 3575 75248
rect 0 75216 800 75246
rect 3509 75243 3575 75246
rect 522021 74490 522087 74493
rect 519892 74488 522087 74490
rect 519892 74432 522026 74488
rect 522082 74432 522087 74488
rect 519892 74430 522087 74432
rect 522021 74427 522087 74430
rect 118417 72994 118483 72997
rect 118417 72992 120060 72994
rect 118417 72936 118422 72992
rect 118478 72936 120060 72992
rect 118417 72934 120060 72936
rect 118417 72931 118483 72934
rect 0 70818 800 70848
rect 3969 70818 4035 70821
rect 0 70816 4035 70818
rect 0 70760 3974 70816
rect 4030 70760 4035 70816
rect 0 70758 4035 70760
rect 0 70728 800 70758
rect 3969 70755 4035 70758
rect 117313 70546 117379 70549
rect 117313 70544 120060 70546
rect 117313 70488 117318 70544
rect 117374 70488 120060 70544
rect 117313 70486 120060 70488
rect 117313 70483 117379 70486
rect 117313 68098 117379 68101
rect 117313 68096 120060 68098
rect 117313 68040 117318 68096
rect 117374 68040 120060 68096
rect 117313 68038 120060 68040
rect 117313 68035 117379 68038
rect 522389 67826 522455 67829
rect 519892 67824 522455 67826
rect 519892 67768 522394 67824
rect 522450 67768 522455 67824
rect 519892 67766 522455 67768
rect 522389 67763 522455 67766
rect 116393 66466 116459 66469
rect 113804 66464 116459 66466
rect 113804 66408 116398 66464
rect 116454 66408 116459 66464
rect 113804 66406 116459 66408
rect 116393 66403 116459 66406
rect 0 66194 800 66224
rect 3325 66194 3391 66197
rect 0 66192 3391 66194
rect 0 66136 3330 66192
rect 3386 66136 3391 66192
rect 0 66134 3391 66136
rect 0 66104 800 66134
rect 3325 66131 3391 66134
rect 117313 65650 117379 65653
rect 117313 65648 120060 65650
rect 117313 65592 117318 65648
rect 117374 65592 120060 65648
rect 117313 65590 120060 65592
rect 117313 65587 117379 65590
rect 117865 63338 117931 63341
rect 117865 63336 120060 63338
rect 117865 63280 117870 63336
rect 117926 63280 120060 63336
rect 117865 63278 120060 63280
rect 117865 63275 117931 63278
rect 0 61570 800 61600
rect 3233 61570 3299 61573
rect 0 61568 3299 61570
rect 0 61512 3238 61568
rect 3294 61512 3299 61568
rect 0 61510 3299 61512
rect 0 61480 800 61510
rect 3233 61507 3299 61510
rect 521837 61026 521903 61029
rect 519892 61024 521903 61026
rect 519892 60968 521842 61024
rect 521898 60968 521903 61024
rect 519892 60966 521903 60968
rect 521837 60963 521903 60966
rect 117773 60890 117839 60893
rect 117773 60888 120060 60890
rect 117773 60832 117778 60888
rect 117834 60832 120060 60888
rect 117773 60830 120060 60832
rect 117773 60827 117839 60830
rect 117313 58442 117379 58445
rect 117313 58440 120060 58442
rect 117313 58384 117318 58440
rect 117374 58384 120060 58440
rect 117313 58382 120060 58384
rect 117313 58379 117379 58382
rect 0 57082 800 57112
rect 2773 57082 2839 57085
rect 0 57080 2839 57082
rect 0 57024 2778 57080
rect 2834 57024 2839 57080
rect 0 57022 2839 57024
rect 0 56992 800 57022
rect 2773 57019 2839 57022
rect 117313 55994 117379 55997
rect 117313 55992 120060 55994
rect 117313 55936 117318 55992
rect 117374 55936 120060 55992
rect 117313 55934 120060 55936
rect 117313 55931 117379 55934
rect 116526 55042 116532 55044
rect 113804 54982 116532 55042
rect 116526 54980 116532 54982
rect 116596 54980 116602 55044
rect 521878 54362 521884 54364
rect 519892 54302 521884 54362
rect 521878 54300 521884 54302
rect 521948 54300 521954 54364
rect 117313 53546 117379 53549
rect 117313 53544 120060 53546
rect 117313 53488 117318 53544
rect 117374 53488 120060 53544
rect 117313 53486 120060 53488
rect 117313 53483 117379 53486
rect 0 52458 800 52488
rect 3141 52458 3207 52461
rect 0 52456 3207 52458
rect 0 52400 3146 52456
rect 3202 52400 3207 52456
rect 0 52398 3207 52400
rect 0 52368 800 52398
rect 3141 52395 3207 52398
rect 117221 51098 117287 51101
rect 117221 51096 120060 51098
rect 117221 51040 117226 51096
rect 117282 51040 120060 51096
rect 117221 51038 120060 51040
rect 117221 51035 117287 51038
rect 117313 48786 117379 48789
rect 117313 48784 120060 48786
rect 117313 48728 117318 48784
rect 117374 48728 120060 48784
rect 117313 48726 120060 48728
rect 117313 48723 117379 48726
rect 0 47970 800 48000
rect 3049 47970 3115 47973
rect 0 47968 3115 47970
rect 0 47912 3054 47968
rect 3110 47912 3115 47968
rect 0 47910 3115 47912
rect 0 47880 800 47910
rect 3049 47907 3115 47910
rect 522113 47562 522179 47565
rect 519892 47560 522179 47562
rect 519892 47504 522118 47560
rect 522174 47504 522179 47560
rect 519892 47502 522179 47504
rect 522113 47499 522179 47502
rect 117865 46338 117931 46341
rect 117865 46336 120060 46338
rect 117865 46280 117870 46336
rect 117926 46280 120060 46336
rect 117865 46278 120060 46280
rect 117865 46275 117931 46278
rect 117221 43890 117287 43893
rect 117221 43888 120060 43890
rect 117221 43832 117226 43888
rect 117282 43832 120060 43888
rect 117221 43830 120060 43832
rect 117221 43827 117287 43830
rect 117129 43754 117195 43757
rect 113804 43752 117195 43754
rect 113804 43696 117134 43752
rect 117190 43696 117195 43752
rect 113804 43694 117195 43696
rect 117129 43691 117195 43694
rect 0 43346 800 43376
rect 2957 43346 3023 43349
rect 0 43344 3023 43346
rect 0 43288 2962 43344
rect 3018 43288 3023 43344
rect 0 43286 3023 43288
rect 0 43256 800 43286
rect 2957 43283 3023 43286
rect 117313 41442 117379 41445
rect 117313 41440 120060 41442
rect 117313 41384 117318 41440
rect 117374 41384 120060 41440
rect 117313 41382 120060 41384
rect 117313 41379 117379 41382
rect 522246 40898 522252 40900
rect 519892 40838 522252 40898
rect 522246 40836 522252 40838
rect 522316 40836 522322 40900
rect 117313 38994 117379 38997
rect 117313 38992 120060 38994
rect 117313 38936 117318 38992
rect 117374 38936 120060 38992
rect 117313 38934 120060 38936
rect 117313 38931 117379 38934
rect 0 38722 800 38752
rect 2865 38722 2931 38725
rect 0 38720 2931 38722
rect 0 38664 2870 38720
rect 2926 38664 2931 38720
rect 0 38662 2931 38664
rect 0 38632 800 38662
rect 2865 38659 2931 38662
rect 117313 36546 117379 36549
rect 117313 36544 120060 36546
rect 117313 36488 117318 36544
rect 117374 36488 120060 36544
rect 117313 36486 120060 36488
rect 117313 36483 117379 36486
rect 0 34234 800 34264
rect 3785 34234 3851 34237
rect 0 34232 3851 34234
rect 0 34176 3790 34232
rect 3846 34176 3851 34232
rect 0 34174 3851 34176
rect 0 34144 800 34174
rect 3785 34171 3851 34174
rect 118417 34234 118483 34237
rect 118417 34232 120060 34234
rect 118417 34176 118422 34232
rect 118478 34176 120060 34232
rect 118417 34174 120060 34176
rect 118417 34171 118483 34174
rect 522573 34098 522639 34101
rect 519892 34096 522639 34098
rect 519892 34040 522578 34096
rect 522634 34040 522639 34096
rect 519892 34038 522639 34040
rect 522573 34035 522639 34038
rect 117037 32330 117103 32333
rect 113804 32328 117103 32330
rect 113804 32272 117042 32328
rect 117098 32272 117103 32328
rect 113804 32270 117103 32272
rect 117037 32267 117103 32270
rect 117313 31786 117379 31789
rect 117313 31784 120060 31786
rect 117313 31728 117318 31784
rect 117374 31728 120060 31784
rect 117313 31726 120060 31728
rect 117313 31723 117379 31726
rect 0 29610 800 29640
rect 2773 29610 2839 29613
rect 0 29608 2839 29610
rect 0 29552 2778 29608
rect 2834 29552 2839 29608
rect 0 29550 2839 29552
rect 0 29520 800 29550
rect 2773 29547 2839 29550
rect 117313 29338 117379 29341
rect 117313 29336 120060 29338
rect 117313 29280 117318 29336
rect 117374 29280 120060 29336
rect 117313 29278 120060 29280
rect 117313 29275 117379 29278
rect 522205 27434 522271 27437
rect 519892 27432 522271 27434
rect 519892 27376 522210 27432
rect 522266 27376 522271 27432
rect 519892 27374 522271 27376
rect 522205 27371 522271 27374
rect 118509 26890 118575 26893
rect 118509 26888 120060 26890
rect 118509 26832 118514 26888
rect 118570 26832 120060 26888
rect 118509 26830 120060 26832
rect 118509 26827 118575 26830
rect 0 25122 800 25152
rect 3693 25122 3759 25125
rect 0 25120 3759 25122
rect 0 25064 3698 25120
rect 3754 25064 3759 25120
rect 0 25062 3759 25064
rect 0 25032 800 25062
rect 3693 25059 3759 25062
rect 117865 24442 117931 24445
rect 117865 24440 120060 24442
rect 117865 24384 117870 24440
rect 117926 24384 120060 24440
rect 117865 24382 120060 24384
rect 117865 24379 117931 24382
rect 117773 21994 117839 21997
rect 117773 21992 120060 21994
rect 117773 21936 117778 21992
rect 117834 21936 120060 21992
rect 117773 21934 120060 21936
rect 117773 21931 117839 21934
rect 117262 20906 117268 20908
rect 113804 20846 117268 20906
rect 117262 20844 117268 20846
rect 117332 20844 117338 20908
rect 0 20498 800 20528
rect 3601 20498 3667 20501
rect 0 20496 3667 20498
rect 0 20440 3606 20496
rect 3662 20440 3667 20496
rect 0 20438 3667 20440
rect 0 20408 800 20438
rect 3601 20435 3667 20438
rect 519862 20090 519922 20604
rect 520222 20090 520228 20092
rect 519862 20030 520228 20090
rect 520222 20028 520228 20030
rect 520292 20028 520298 20092
rect 117129 19682 117195 19685
rect 117129 19680 120060 19682
rect 117129 19624 117134 19680
rect 117190 19624 120060 19680
rect 117129 19622 120060 19624
rect 117129 19619 117195 19622
rect 117497 17234 117563 17237
rect 117497 17232 120060 17234
rect 117497 17176 117502 17232
rect 117558 17176 120060 17232
rect 117497 17174 120060 17176
rect 117497 17171 117563 17174
rect 0 15874 800 15904
rect 3877 15874 3943 15877
rect 0 15872 3943 15874
rect 0 15816 3882 15872
rect 3938 15816 3943 15872
rect 0 15814 3943 15816
rect 0 15784 800 15814
rect 3877 15811 3943 15814
rect 117313 14786 117379 14789
rect 117313 14784 120060 14786
rect 117313 14728 117318 14784
rect 117374 14728 120060 14784
rect 117313 14726 120060 14728
rect 117313 14723 117379 14726
rect 522665 13970 522731 13973
rect 519892 13968 522731 13970
rect 519892 13912 522670 13968
rect 522726 13912 522731 13968
rect 519892 13910 522731 13912
rect 522665 13907 522731 13910
rect 117221 12338 117287 12341
rect 117221 12336 120060 12338
rect 117221 12280 117226 12336
rect 117282 12280 120060 12336
rect 117221 12278 120060 12280
rect 117221 12275 117287 12278
rect 0 11386 800 11416
rect 3969 11386 4035 11389
rect 0 11384 4035 11386
rect 0 11328 3974 11384
rect 4030 11328 4035 11384
rect 0 11326 4035 11328
rect 0 11296 800 11326
rect 3969 11323 4035 11326
rect 117313 9890 117379 9893
rect 117313 9888 120060 9890
rect 117313 9832 117318 9888
rect 117374 9832 120060 9888
rect 117313 9830 120060 9832
rect 117313 9827 117379 9830
rect 116025 9618 116091 9621
rect 113804 9616 116091 9618
rect 113804 9560 116030 9616
rect 116086 9560 116091 9616
rect 113804 9558 116091 9560
rect 116025 9555 116091 9558
rect 117313 7442 117379 7445
rect 117313 7440 120060 7442
rect 117313 7384 117318 7440
rect 117374 7384 120060 7440
rect 117313 7382 120060 7384
rect 117313 7379 117379 7382
rect 521653 7306 521719 7309
rect 519892 7304 521719 7306
rect 519892 7248 521658 7304
rect 521714 7248 521719 7304
rect 519892 7246 521719 7248
rect 521653 7243 521719 7246
rect 0 6762 800 6792
rect 3233 6762 3299 6765
rect 0 6760 3299 6762
rect 0 6704 3238 6760
rect 3294 6704 3299 6760
rect 0 6702 3299 6704
rect 0 6672 800 6702
rect 3233 6699 3299 6702
rect 4797 6082 4863 6085
rect 118417 6082 118483 6085
rect 4797 6080 118483 6082
rect 4797 6024 4802 6080
rect 4858 6024 118422 6080
rect 118478 6024 118483 6080
rect 4797 6022 118483 6024
rect 4797 6019 4863 6022
rect 118417 6019 118483 6022
rect 117313 5130 117379 5133
rect 117313 5128 120060 5130
rect 117313 5072 117318 5128
rect 117374 5072 120060 5128
rect 117313 5070 120060 5072
rect 117313 5067 117379 5070
rect 3601 4994 3667 4997
rect 521653 4994 521719 4997
rect 3601 4992 521719 4994
rect 3601 4936 3606 4992
rect 3662 4936 521658 4992
rect 521714 4936 521719 4992
rect 3601 4934 521719 4936
rect 3601 4931 3667 4934
rect 521653 4931 521719 4934
rect 522021 4858 522087 4861
rect 45510 4856 522087 4858
rect 45510 4800 522026 4856
rect 522082 4800 522087 4856
rect 45510 4798 522087 4800
rect 39297 4586 39363 4589
rect 45510 4586 45570 4798
rect 522021 4795 522087 4798
rect 520549 4722 520615 4725
rect 50294 4720 520615 4722
rect 50294 4664 520554 4720
rect 520610 4664 520615 4720
rect 50294 4662 520615 4664
rect 39297 4584 45570 4586
rect 39297 4528 39302 4584
rect 39358 4528 45570 4584
rect 39297 4526 45570 4528
rect 45921 4586 45987 4589
rect 50294 4586 50354 4662
rect 520549 4659 520615 4662
rect 45921 4584 50354 4586
rect 45921 4528 45926 4584
rect 45982 4528 50354 4584
rect 45921 4526 50354 4528
rect 52453 4586 52519 4589
rect 521929 4586 521995 4589
rect 52453 4584 521995 4586
rect 52453 4528 52458 4584
rect 52514 4528 521934 4584
rect 521990 4528 521995 4584
rect 52453 4526 521995 4528
rect 39297 4523 39363 4526
rect 45921 4523 45987 4526
rect 52453 4523 52519 4526
rect 521929 4523 521995 4526
rect 75821 4450 75887 4453
rect 520641 4450 520707 4453
rect 75821 4448 520707 4450
rect 75821 4392 75826 4448
rect 75882 4392 520646 4448
rect 520702 4392 520707 4448
rect 75821 4390 520707 4392
rect 75821 4387 75887 4390
rect 520641 4387 520707 4390
rect 116945 3498 117011 3501
rect 426341 3498 426407 3501
rect 116945 3496 426407 3498
rect 116945 3440 116950 3496
rect 117006 3440 426346 3496
rect 426402 3440 426407 3496
rect 116945 3438 426407 3440
rect 116945 3435 117011 3438
rect 426341 3435 426407 3438
rect 118601 3362 118667 3365
rect 550541 3362 550607 3365
rect 118601 3360 550607 3362
rect 118601 3304 118606 3360
rect 118662 3304 550546 3360
rect 550602 3304 550607 3360
rect 118601 3302 550607 3304
rect 118601 3299 118667 3302
rect 550541 3299 550607 3302
rect 5993 2682 6059 2685
rect 119521 2682 119587 2685
rect 5993 2680 119587 2682
rect 5993 2624 5998 2680
rect 6054 2624 119526 2680
rect 119582 2624 119587 2680
rect 5993 2622 119587 2624
rect 5993 2619 6059 2622
rect 119521 2619 119587 2622
rect 12341 2546 12407 2549
rect 119705 2546 119771 2549
rect 12341 2544 119771 2546
rect 12341 2488 12346 2544
rect 12402 2488 119710 2544
rect 119766 2488 119771 2544
rect 12341 2486 119771 2488
rect 12341 2483 12407 2486
rect 119705 2483 119771 2486
rect 28901 2410 28967 2413
rect 119337 2410 119403 2413
rect 28901 2408 119403 2410
rect 28901 2352 28906 2408
rect 28962 2352 119342 2408
rect 119398 2352 119403 2408
rect 28901 2350 119403 2352
rect 28901 2347 28967 2350
rect 119337 2347 119403 2350
rect 0 2274 800 2304
rect 2957 2274 3023 2277
rect 0 2272 3023 2274
rect 0 2216 2962 2272
rect 3018 2216 3023 2272
rect 0 2214 3023 2216
rect 0 2184 800 2214
rect 2957 2211 3023 2214
<< via3 >>
rect 9444 153368 9508 153372
rect 9444 153312 9458 153368
rect 9458 153312 9508 153368
rect 9444 153308 9508 153312
rect 506428 153232 506492 153236
rect 506428 153176 506478 153232
rect 506478 153176 506492 153232
rect 506428 153172 506492 153176
rect 117452 77828 117516 77892
rect 116532 54980 116596 55044
rect 521884 54300 521948 54364
rect 522252 40836 522316 40900
rect 117268 20844 117332 20908
rect 520228 20028 520292 20092
<< metal4 >>
rect 4208 154000 4528 157760
rect 9208 154000 9528 157760
rect 14208 154000 14528 157760
rect 19208 154000 19528 157760
rect 24208 154000 24528 157760
rect 29208 154000 29528 157760
rect 34208 154000 34528 157760
rect 39208 154000 39528 157760
rect 44208 154000 44528 157760
rect 49208 154000 49528 157760
rect 54208 154000 54528 157760
rect 59208 154000 59528 157760
rect 64208 154000 64528 157760
rect 69208 154000 69528 157760
rect 74208 154000 74528 157760
rect 79208 154000 79528 157760
rect 84208 154000 84528 157760
rect 89208 154000 89528 157760
rect 94208 154000 94528 157760
rect 99208 154000 99528 157760
rect 104208 154000 104528 157760
rect 109208 154000 109528 157760
rect 114208 154000 114528 157760
rect 119208 154000 119528 157760
rect 124208 154000 124528 157760
rect 129208 154000 129528 157760
rect 134208 154000 134528 157760
rect 139208 154000 139528 157760
rect 144208 154000 144528 157760
rect 149208 154000 149528 157760
rect 154208 154000 154528 157760
rect 159208 154000 159528 157760
rect 164208 154000 164528 157760
rect 169208 154000 169528 157760
rect 174208 154000 174528 157760
rect 179208 154000 179528 157760
rect 184208 154000 184528 157760
rect 189208 154000 189528 157760
rect 194208 154000 194528 157760
rect 199208 154000 199528 157760
rect 204208 154000 204528 157760
rect 209208 154000 209528 157760
rect 214208 154000 214528 157760
rect 219208 154000 219528 157760
rect 224208 154000 224528 157760
rect 229208 154000 229528 157760
rect 234208 154000 234528 157760
rect 239208 154000 239528 157760
rect 244208 154000 244528 157760
rect 249208 154000 249528 157760
rect 254208 154000 254528 157760
rect 259208 154000 259528 157760
rect 264208 154000 264528 157760
rect 269208 154000 269528 157760
rect 274208 154000 274528 157760
rect 279208 154000 279528 157760
rect 284208 154000 284528 157760
rect 289208 154000 289528 157760
rect 294208 154000 294528 157760
rect 299208 154000 299528 157760
rect 304208 154000 304528 157760
rect 309208 154000 309528 157760
rect 314208 154000 314528 157760
rect 319208 154000 319528 157760
rect 324208 154000 324528 157760
rect 329208 154000 329528 157760
rect 334208 154000 334528 157760
rect 339208 154000 339528 157760
rect 344208 154000 344528 157760
rect 349208 154000 349528 157760
rect 354208 154000 354528 157760
rect 359208 154000 359528 157760
rect 364208 154000 364528 157760
rect 369208 154000 369528 157760
rect 374208 154000 374528 157760
rect 379208 154000 379528 157760
rect 384208 154000 384528 157760
rect 389208 154000 389528 157760
rect 394208 154000 394528 157760
rect 399208 154000 399528 157760
rect 404208 154000 404528 157760
rect 409208 154000 409528 157760
rect 414208 154000 414528 157760
rect 419208 154000 419528 157760
rect 424208 154000 424528 157760
rect 429208 154000 429528 157760
rect 434208 154000 434528 157760
rect 439208 154000 439528 157760
rect 444208 154000 444528 157760
rect 449208 154000 449528 157760
rect 454208 154000 454528 157760
rect 459208 154000 459528 157760
rect 464208 154000 464528 157760
rect 469208 154000 469528 157760
rect 474208 154000 474528 157760
rect 479208 154000 479528 157760
rect 484208 154000 484528 157760
rect 489208 154000 489528 157760
rect 494208 154000 494528 157760
rect 499208 154000 499528 157760
rect 504208 154000 504528 157760
rect 509208 154000 509528 157760
rect 514208 154000 514528 157760
rect 519208 154000 519528 157760
rect 506427 153172 506428 153222
rect 506492 153172 506493 153222
rect 506427 153171 506493 153172
rect 524208 135624 524528 157760
rect 524208 135388 524250 135624
rect 524486 135388 524528 135624
rect 524208 109624 524528 135388
rect 524208 109388 524250 109624
rect 524486 109388 524528 109624
rect 524208 83624 524528 109388
rect 524208 83388 524250 83624
rect 524486 83388 524528 83624
rect 117451 77892 117517 77893
rect 117451 77828 117452 77892
rect 117516 77828 117517 77892
rect 117451 77827 117517 77828
rect 117454 75258 117514 77827
rect 116534 55045 116594 62102
rect 116531 55044 116597 55045
rect 116531 54980 116532 55044
rect 116596 54980 116597 55044
rect 116531 54979 116597 54980
rect 521886 54365 521946 73662
rect 521883 54364 521949 54365
rect 521883 54300 521884 54364
rect 521948 54300 521949 54364
rect 521883 54299 521949 54300
rect 522254 40901 522314 60742
rect 524208 57624 524528 83388
rect 524208 57388 524250 57624
rect 524486 57388 524528 57624
rect 522251 40900 522317 40901
rect 522251 40836 522252 40900
rect 522316 40836 522317 40900
rect 522251 40835 522317 40836
rect 524208 31624 524528 57388
rect 524208 31388 524250 31624
rect 524486 31388 524528 31624
rect 117267 20908 117333 20909
rect 117267 20844 117268 20908
rect 117332 20844 117333 20908
rect 117267 20843 117333 20844
rect 117270 20178 117330 20843
rect 524208 5624 524528 31388
rect 524208 5388 524250 5624
rect 524486 5388 524528 5624
rect 524208 2176 524528 5388
rect 529208 148624 529528 157760
rect 529208 148388 529250 148624
rect 529486 148388 529528 148624
rect 529208 122624 529528 148388
rect 529208 122388 529250 122624
rect 529486 122388 529528 122624
rect 529208 96624 529528 122388
rect 529208 96388 529250 96624
rect 529486 96388 529528 96624
rect 529208 70624 529528 96388
rect 529208 70388 529250 70624
rect 529486 70388 529528 70624
rect 529208 44624 529528 70388
rect 529208 44388 529250 44624
rect 529486 44388 529528 44624
rect 529208 18624 529528 44388
rect 529208 18388 529250 18624
rect 529486 18388 529528 18624
rect 529208 2176 529528 18388
rect 534208 135624 534528 157760
rect 534208 135388 534250 135624
rect 534486 135388 534528 135624
rect 534208 109624 534528 135388
rect 534208 109388 534250 109624
rect 534486 109388 534528 109624
rect 534208 83624 534528 109388
rect 534208 83388 534250 83624
rect 534486 83388 534528 83624
rect 534208 57624 534528 83388
rect 534208 57388 534250 57624
rect 534486 57388 534528 57624
rect 534208 31624 534528 57388
rect 534208 31388 534250 31624
rect 534486 31388 534528 31624
rect 534208 5624 534528 31388
rect 534208 5388 534250 5624
rect 534486 5388 534528 5624
rect 534208 2176 534528 5388
rect 539208 148624 539528 157760
rect 539208 148388 539250 148624
rect 539486 148388 539528 148624
rect 539208 122624 539528 148388
rect 539208 122388 539250 122624
rect 539486 122388 539528 122624
rect 539208 96624 539528 122388
rect 539208 96388 539250 96624
rect 539486 96388 539528 96624
rect 539208 70624 539528 96388
rect 539208 70388 539250 70624
rect 539486 70388 539528 70624
rect 539208 44624 539528 70388
rect 539208 44388 539250 44624
rect 539486 44388 539528 44624
rect 539208 18624 539528 44388
rect 539208 18388 539250 18624
rect 539486 18388 539528 18624
rect 539208 2176 539528 18388
rect 544208 135624 544528 157760
rect 544208 135388 544250 135624
rect 544486 135388 544528 135624
rect 544208 109624 544528 135388
rect 544208 109388 544250 109624
rect 544486 109388 544528 109624
rect 544208 83624 544528 109388
rect 544208 83388 544250 83624
rect 544486 83388 544528 83624
rect 544208 57624 544528 83388
rect 544208 57388 544250 57624
rect 544486 57388 544528 57624
rect 544208 31624 544528 57388
rect 544208 31388 544250 31624
rect 544486 31388 544528 31624
rect 544208 5624 544528 31388
rect 544208 5388 544250 5624
rect 544486 5388 544528 5624
rect 544208 2176 544528 5388
rect 549208 148624 549528 157760
rect 549208 148388 549250 148624
rect 549486 148388 549528 148624
rect 549208 122624 549528 148388
rect 549208 122388 549250 122624
rect 549486 122388 549528 122624
rect 549208 96624 549528 122388
rect 549208 96388 549250 96624
rect 549486 96388 549528 96624
rect 549208 70624 549528 96388
rect 549208 70388 549250 70624
rect 549486 70388 549528 70624
rect 549208 44624 549528 70388
rect 549208 44388 549250 44624
rect 549486 44388 549528 44624
rect 549208 18624 549528 44388
rect 549208 18388 549250 18624
rect 549486 18388 549528 18624
rect 549208 2176 549528 18388
rect 554208 135624 554528 157760
rect 554208 135388 554250 135624
rect 554486 135388 554528 135624
rect 554208 109624 554528 135388
rect 554208 109388 554250 109624
rect 554486 109388 554528 109624
rect 554208 83624 554528 109388
rect 554208 83388 554250 83624
rect 554486 83388 554528 83624
rect 554208 57624 554528 83388
rect 554208 57388 554250 57624
rect 554486 57388 554528 57624
rect 554208 31624 554528 57388
rect 554208 31388 554250 31624
rect 554486 31388 554528 31624
rect 554208 5624 554528 31388
rect 554208 5388 554250 5624
rect 554486 5388 554528 5624
rect 554208 2176 554528 5388
rect 559208 148624 559528 157760
rect 559208 148388 559250 148624
rect 559486 148388 559528 148624
rect 559208 122624 559528 148388
rect 559208 122388 559250 122624
rect 559486 122388 559528 122624
rect 559208 96624 559528 122388
rect 559208 96388 559250 96624
rect 559486 96388 559528 96624
rect 559208 70624 559528 96388
rect 559208 70388 559250 70624
rect 559486 70388 559528 70624
rect 559208 44624 559528 70388
rect 559208 44388 559250 44624
rect 559486 44388 559528 44624
rect 559208 18624 559528 44388
rect 559208 18388 559250 18624
rect 559486 18388 559528 18624
rect 559208 2176 559528 18388
rect 564208 135624 564528 157760
rect 564208 135388 564250 135624
rect 564486 135388 564528 135624
rect 564208 109624 564528 135388
rect 564208 109388 564250 109624
rect 564486 109388 564528 109624
rect 564208 83624 564528 109388
rect 564208 83388 564250 83624
rect 564486 83388 564528 83624
rect 564208 57624 564528 83388
rect 564208 57388 564250 57624
rect 564486 57388 564528 57624
rect 564208 31624 564528 57388
rect 564208 31388 564250 31624
rect 564486 31388 564528 31624
rect 564208 5624 564528 31388
rect 564208 5388 564250 5624
rect 564486 5388 564528 5624
rect 564208 2176 564528 5388
rect 569208 148624 569528 157760
rect 569208 148388 569250 148624
rect 569486 148388 569528 148624
rect 569208 122624 569528 148388
rect 569208 122388 569250 122624
rect 569486 122388 569528 122624
rect 569208 96624 569528 122388
rect 569208 96388 569250 96624
rect 569486 96388 569528 96624
rect 569208 70624 569528 96388
rect 569208 70388 569250 70624
rect 569486 70388 569528 70624
rect 569208 44624 569528 70388
rect 569208 44388 569250 44624
rect 569486 44388 569528 44624
rect 569208 18624 569528 44388
rect 569208 18388 569250 18624
rect 569486 18388 569528 18624
rect 569208 2176 569528 18388
rect 574208 135624 574528 157760
rect 574208 135388 574250 135624
rect 574486 135388 574528 135624
rect 574208 109624 574528 135388
rect 574208 109388 574250 109624
rect 574486 109388 574528 109624
rect 574208 83624 574528 109388
rect 574208 83388 574250 83624
rect 574486 83388 574528 83624
rect 574208 57624 574528 83388
rect 574208 57388 574250 57624
rect 574486 57388 574528 57624
rect 574208 31624 574528 57388
rect 574208 31388 574250 31624
rect 574486 31388 574528 31624
rect 574208 5624 574528 31388
rect 574208 5388 574250 5624
rect 574486 5388 574528 5624
rect 574208 2176 574528 5388
<< via4 >>
rect 9358 153372 9594 153458
rect 9358 153308 9444 153372
rect 9444 153308 9508 153372
rect 9508 153308 9594 153372
rect 9358 153222 9594 153308
rect 506342 153236 506578 153458
rect 506342 153222 506428 153236
rect 506428 153222 506492 153236
rect 506492 153222 506578 153236
rect 524250 135388 524486 135624
rect 524250 109388 524486 109624
rect 524250 83388 524486 83624
rect 117366 75022 117602 75258
rect 521798 73662 522034 73898
rect 116446 62102 116682 62338
rect 522166 60742 522402 60978
rect 524250 57388 524486 57624
rect 524250 31388 524486 31624
rect 117182 19942 117418 20178
rect 520142 20092 520378 20178
rect 520142 20028 520228 20092
rect 520228 20028 520292 20092
rect 520292 20028 520378 20092
rect 520142 19942 520378 20028
rect 524250 5388 524486 5624
rect 529250 148388 529486 148624
rect 529250 122388 529486 122624
rect 529250 96388 529486 96624
rect 529250 70388 529486 70624
rect 529250 44388 529486 44624
rect 529250 18388 529486 18624
rect 534250 135388 534486 135624
rect 534250 109388 534486 109624
rect 534250 83388 534486 83624
rect 534250 57388 534486 57624
rect 534250 31388 534486 31624
rect 534250 5388 534486 5624
rect 539250 148388 539486 148624
rect 539250 122388 539486 122624
rect 539250 96388 539486 96624
rect 539250 70388 539486 70624
rect 539250 44388 539486 44624
rect 539250 18388 539486 18624
rect 544250 135388 544486 135624
rect 544250 109388 544486 109624
rect 544250 83388 544486 83624
rect 544250 57388 544486 57624
rect 544250 31388 544486 31624
rect 544250 5388 544486 5624
rect 549250 148388 549486 148624
rect 549250 122388 549486 122624
rect 549250 96388 549486 96624
rect 549250 70388 549486 70624
rect 549250 44388 549486 44624
rect 549250 18388 549486 18624
rect 554250 135388 554486 135624
rect 554250 109388 554486 109624
rect 554250 83388 554486 83624
rect 554250 57388 554486 57624
rect 554250 31388 554486 31624
rect 554250 5388 554486 5624
rect 559250 148388 559486 148624
rect 559250 122388 559486 122624
rect 559250 96388 559486 96624
rect 559250 70388 559486 70624
rect 559250 44388 559486 44624
rect 559250 18388 559486 18624
rect 564250 135388 564486 135624
rect 564250 109388 564486 109624
rect 564250 83388 564486 83624
rect 564250 57388 564486 57624
rect 564250 31388 564486 31624
rect 564250 5388 564486 5624
rect 569250 148388 569486 148624
rect 569250 122388 569486 122624
rect 569250 96388 569486 96624
rect 569250 70388 569486 70624
rect 569250 44388 569486 44624
rect 569250 18388 569486 18624
rect 574250 135388 574486 135624
rect 574250 109388 574486 109624
rect 574250 83388 574486 83624
rect 574250 57388 574486 57624
rect 574250 31388 574486 31624
rect 574250 5388 574486 5624
<< metal5 >>
rect 9316 153458 506620 153500
rect 9316 153222 9358 153458
rect 9594 153222 506342 153458
rect 506578 153222 506620 153458
rect 9316 153180 506620 153222
rect 1104 148346 2000 148666
rect 116000 148346 118000 148666
rect 522000 148624 578864 148666
rect 522000 148388 529250 148624
rect 529486 148388 539250 148624
rect 539486 148388 549250 148624
rect 549486 148388 559250 148624
rect 559486 148388 569250 148624
rect 569486 148388 578864 148624
rect 522000 148346 578864 148388
rect 1104 135346 2000 135666
rect 116000 135346 118000 135666
rect 522000 135624 578864 135666
rect 522000 135388 524250 135624
rect 524486 135388 534250 135624
rect 534486 135388 544250 135624
rect 544486 135388 554250 135624
rect 554486 135388 564250 135624
rect 564486 135388 574250 135624
rect 574486 135388 578864 135624
rect 522000 135346 578864 135388
rect 1104 122346 2000 122666
rect 116000 122346 118000 122666
rect 522000 122624 578864 122666
rect 522000 122388 529250 122624
rect 529486 122388 539250 122624
rect 539486 122388 549250 122624
rect 549486 122388 559250 122624
rect 559486 122388 569250 122624
rect 569486 122388 578864 122624
rect 522000 122346 578864 122388
rect 1104 109346 2000 109666
rect 116000 109346 118000 109666
rect 522000 109624 578864 109666
rect 522000 109388 524250 109624
rect 524486 109388 534250 109624
rect 534486 109388 544250 109624
rect 544486 109388 554250 109624
rect 554486 109388 564250 109624
rect 564486 109388 574250 109624
rect 574486 109388 578864 109624
rect 522000 109346 578864 109388
rect 1104 96346 2000 96666
rect 116000 96346 118000 96666
rect 522000 96624 578864 96666
rect 522000 96388 529250 96624
rect 529486 96388 539250 96624
rect 539486 96388 549250 96624
rect 549486 96388 559250 96624
rect 559486 96388 569250 96624
rect 569486 96388 578864 96624
rect 522000 96346 578864 96388
rect 1104 83346 2000 83666
rect 116000 83346 118000 83666
rect 522000 83624 578864 83666
rect 522000 83388 524250 83624
rect 524486 83388 534250 83624
rect 534486 83388 544250 83624
rect 544486 83388 554250 83624
rect 554486 83388 564250 83624
rect 564486 83388 574250 83624
rect 574486 83388 578864 83624
rect 522000 83346 578864 83388
rect 117324 75258 123348 75300
rect 117324 75022 117366 75258
rect 117602 75022 123348 75258
rect 117324 74980 123348 75022
rect 123028 74620 123348 74980
rect 123028 74300 393276 74620
rect 392956 73940 393276 74300
rect 392956 73898 522076 73940
rect 392956 73662 521798 73898
rect 522034 73662 522076 73898
rect 392956 73620 522076 73662
rect 1104 70346 2000 70666
rect 116000 70346 118000 70666
rect 522000 70624 578864 70666
rect 522000 70388 529250 70624
rect 529486 70388 539250 70624
rect 539486 70388 549250 70624
rect 549486 70388 559250 70624
rect 559486 70388 569250 70624
rect 569486 70388 578864 70624
rect 522000 70346 578864 70388
rect 116404 62338 123164 62380
rect 116404 62102 116446 62338
rect 116682 62102 123164 62338
rect 116404 62060 123164 62102
rect 122844 61700 123164 62060
rect 122844 61380 393276 61700
rect 392956 60340 393276 61380
rect 520100 60978 522444 61020
rect 520100 60742 522166 60978
rect 522402 60742 522444 60978
rect 520100 60700 522444 60742
rect 520100 60340 520420 60700
rect 392956 60020 520420 60340
rect 1104 57346 2000 57666
rect 116000 57346 118000 57666
rect 522000 57624 578864 57666
rect 522000 57388 524250 57624
rect 524486 57388 534250 57624
rect 534486 57388 544250 57624
rect 544486 57388 554250 57624
rect 554486 57388 564250 57624
rect 564486 57388 574250 57624
rect 574486 57388 578864 57624
rect 522000 57346 578864 57388
rect 1104 44346 2000 44666
rect 116000 44346 118000 44666
rect 522000 44624 578864 44666
rect 522000 44388 529250 44624
rect 529486 44388 539250 44624
rect 539486 44388 549250 44624
rect 549486 44388 559250 44624
rect 559486 44388 569250 44624
rect 569486 44388 578864 44624
rect 522000 44346 578864 44388
rect 1104 31346 2000 31666
rect 116000 31346 118000 31666
rect 522000 31624 578864 31666
rect 522000 31388 524250 31624
rect 524486 31388 534250 31624
rect 534486 31388 544250 31624
rect 544486 31388 554250 31624
rect 554486 31388 564250 31624
rect 564486 31388 574250 31624
rect 574486 31388 578864 31624
rect 522000 31346 578864 31388
rect 117140 20178 520420 20220
rect 117140 19942 117182 20178
rect 117418 19942 520142 20178
rect 520378 19942 520420 20178
rect 117140 19900 520420 19942
rect 1104 18346 2000 18666
rect 116000 18346 118000 18666
rect 522000 18624 578864 18666
rect 522000 18388 529250 18624
rect 529486 18388 539250 18624
rect 539486 18388 549250 18624
rect 549486 18388 559250 18624
rect 559486 18388 569250 18624
rect 569486 18388 578864 18624
rect 522000 18346 578864 18388
rect 1104 5346 2000 5666
rect 116000 5346 118000 5666
rect 522000 5624 578864 5666
rect 522000 5388 524250 5624
rect 524486 5388 534250 5624
rect 534486 5388 544250 5624
rect 544486 5388 554250 5624
rect 554486 5388 564250 5624
rect 564486 5388 574250 5624
rect 574486 5388 578864 5624
rect 522000 5346 578864 5388
use mgmt_core  core
timestamp 1638169271
transform 1 0 120000 0 1 4000
box 0 0 400000 148000
use DFFRAM  DFFRAM
timestamp 1638169271
transform 1 0 4000 0 1 4000
box 4 0 110000 148000
<< labels >>
rlabel metal5 s 1104 18346 2000 18666 6 VGND
port 0 nsew ground input
rlabel metal5 s 116000 18346 118000 18666 6 VGND
port 0 nsew ground input
rlabel metal5 s 522000 18346 578864 18666 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 44346 2000 44666 6 VGND
port 0 nsew ground input
rlabel metal5 s 116000 44346 118000 44666 6 VGND
port 0 nsew ground input
rlabel metal5 s 522000 44346 578864 44666 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 70346 2000 70666 6 VGND
port 0 nsew ground input
rlabel metal5 s 116000 70346 118000 70666 6 VGND
port 0 nsew ground input
rlabel metal5 s 522000 70346 578864 70666 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 96346 2000 96666 6 VGND
port 0 nsew ground input
rlabel metal5 s 116000 96346 118000 96666 6 VGND
port 0 nsew ground input
rlabel metal5 s 522000 96346 578864 96666 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 122346 2000 122666 6 VGND
port 0 nsew ground input
rlabel metal5 s 116000 122346 118000 122666 6 VGND
port 0 nsew ground input
rlabel metal5 s 522000 122346 578864 122666 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 148346 2000 148666 6 VGND
port 0 nsew ground input
rlabel metal5 s 116000 148346 118000 148666 6 VGND
port 0 nsew ground input
rlabel metal5 s 522000 148346 578864 148666 6 VGND
port 0 nsew ground input
rlabel metal4 s 9208 154000 9528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 19208 154000 19528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 29208 154000 29528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 39208 154000 39528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 49208 154000 49528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 59208 154000 59528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 69208 154000 69528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 79208 154000 79528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 89208 154000 89528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 99208 154000 99528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 109208 154000 109528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 119208 154000 119528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 129208 154000 129528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 139208 154000 139528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 149208 154000 149528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 159208 154000 159528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 169208 154000 169528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 179208 154000 179528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 189208 154000 189528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 199208 154000 199528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 209208 154000 209528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 219208 154000 219528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 229208 154000 229528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 239208 154000 239528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 249208 154000 249528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 259208 154000 259528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 269208 154000 269528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 279208 154000 279528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 289208 154000 289528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 299208 154000 299528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 309208 154000 309528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 319208 154000 319528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 329208 154000 329528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 339208 154000 339528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 349208 154000 349528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 359208 154000 359528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 369208 154000 369528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 379208 154000 379528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 389208 154000 389528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 399208 154000 399528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 409208 154000 409528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 419208 154000 419528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 429208 154000 429528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 439208 154000 439528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 449208 154000 449528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 459208 154000 459528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 469208 154000 469528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 479208 154000 479528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 489208 154000 489528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 499208 154000 499528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 509208 154000 509528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 519208 154000 519528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 529208 2176 529528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 539208 2176 539528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 549208 2176 549528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 559208 2176 559528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 569208 2176 569528 157760 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 5346 2000 5666 6 VPWR
port 1 nsew power input
rlabel metal5 s 116000 5346 118000 5666 6 VPWR
port 1 nsew power input
rlabel metal5 s 522000 5346 578864 5666 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 31346 2000 31666 6 VPWR
port 1 nsew power input
rlabel metal5 s 116000 31346 118000 31666 6 VPWR
port 1 nsew power input
rlabel metal5 s 522000 31346 578864 31666 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 57346 2000 57666 6 VPWR
port 1 nsew power input
rlabel metal5 s 116000 57346 118000 57666 6 VPWR
port 1 nsew power input
rlabel metal5 s 522000 57346 578864 57666 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 83346 2000 83666 6 VPWR
port 1 nsew power input
rlabel metal5 s 116000 83346 118000 83666 6 VPWR
port 1 nsew power input
rlabel metal5 s 522000 83346 578864 83666 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 109346 2000 109666 6 VPWR
port 1 nsew power input
rlabel metal5 s 116000 109346 118000 109666 6 VPWR
port 1 nsew power input
rlabel metal5 s 522000 109346 578864 109666 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 135346 2000 135666 6 VPWR
port 1 nsew power input
rlabel metal5 s 116000 135346 118000 135666 6 VPWR
port 1 nsew power input
rlabel metal5 s 522000 135346 578864 135666 6 VPWR
port 1 nsew power input
rlabel metal4 s 4208 154000 4528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 14208 154000 14528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 24208 154000 24528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 34208 154000 34528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 44208 154000 44528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 54208 154000 54528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 64208 154000 64528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 74208 154000 74528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 84208 154000 84528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 94208 154000 94528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 104208 154000 104528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 114208 154000 114528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 124208 154000 124528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 134208 154000 134528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 144208 154000 144528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 154208 154000 154528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 164208 154000 164528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 174208 154000 174528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 184208 154000 184528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 194208 154000 194528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 204208 154000 204528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 214208 154000 214528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 224208 154000 224528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 234208 154000 234528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 244208 154000 244528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 254208 154000 254528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 264208 154000 264528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 274208 154000 274528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 284208 154000 284528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 294208 154000 294528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 304208 154000 304528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 314208 154000 314528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 324208 154000 324528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 334208 154000 334528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 344208 154000 344528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 354208 154000 354528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 364208 154000 364528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 374208 154000 374528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 384208 154000 384528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 394208 154000 394528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 404208 154000 404528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 414208 154000 414528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 424208 154000 424528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 434208 154000 434528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 444208 154000 444528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 454208 154000 454528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 464208 154000 464528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 474208 154000 474528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 484208 154000 484528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 494208 154000 494528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 504208 154000 504528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 514208 154000 514528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 524208 2176 524528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 534208 2176 534528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 544208 2176 544528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 554208 2176 554528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 564208 2176 564528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 574208 2176 574528 157760 6 VPWR
port 1 nsew power input
rlabel metal2 s 478 159200 534 160000 6 core_clk
port 2 nsew signal input
rlabel metal2 s 1398 159200 1454 160000 6 core_rstn
port 3 nsew signal input
rlabel metal2 s 508042 0 508098 800 6 debug_in
port 4 nsew signal input
rlabel metal2 s 513378 0 513434 800 6 debug_mode
port 5 nsew signal tristate
rlabel metal2 s 523958 0 524014 800 6 debug_oeb
port 6 nsew signal tristate
rlabel metal2 s 518622 0 518678 800 6 debug_out
port 7 nsew signal tristate
rlabel metal2 s 39762 0 39818 800 6 flash_clk
port 8 nsew signal tristate
rlabel metal2 s 34518 0 34574 800 6 flash_csb
port 9 nsew signal tristate
rlabel metal2 s 45098 0 45154 800 6 flash_io0_di
port 10 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 flash_io0_do
port 11 nsew signal tristate
rlabel metal2 s 55770 0 55826 800 6 flash_io0_oeb
port 12 nsew signal tristate
rlabel metal2 s 61106 0 61162 800 6 flash_io1_di
port 13 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 flash_io1_do
port 14 nsew signal tristate
rlabel metal2 s 71686 0 71742 800 6 flash_io1_oeb
port 15 nsew signal tristate
rlabel metal2 s 77022 0 77078 800 6 flash_io2_di
port 16 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 flash_io2_do
port 17 nsew signal tristate
rlabel metal3 s 0 6672 800 6792 6 flash_io2_oeb
port 18 nsew signal tristate
rlabel metal2 s 87694 0 87750 800 6 flash_io3_di
port 19 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 flash_io3_do
port 20 nsew signal tristate
rlabel metal3 s 0 2184 800 2304 6 flash_io3_oeb
port 21 nsew signal tristate
rlabel metal2 s 2594 0 2650 800 6 gpio_in_pad
port 22 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 gpio_inenb_pad
port 23 nsew signal tristate
rlabel metal2 s 13174 0 13230 800 6 gpio_mode0_pad
port 24 nsew signal tristate
rlabel metal2 s 18510 0 18566 800 6 gpio_mode1_pad
port 25 nsew signal tristate
rlabel metal2 s 23846 0 23902 800 6 gpio_out_pad
port 26 nsew signal tristate
rlabel metal2 s 29182 0 29238 800 6 gpio_outenb_pad
port 27 nsew signal tristate
rlabel metal2 s 103610 0 103666 800 6 hk_ack_i
port 28 nsew signal input
rlabel metal2 s 114282 0 114338 800 6 hk_dat_i[0]
port 29 nsew signal input
rlabel metal2 s 167458 0 167514 800 6 hk_dat_i[10]
port 30 nsew signal input
rlabel metal2 s 172794 0 172850 800 6 hk_dat_i[11]
port 31 nsew signal input
rlabel metal2 s 178130 0 178186 800 6 hk_dat_i[12]
port 32 nsew signal input
rlabel metal2 s 183466 0 183522 800 6 hk_dat_i[13]
port 33 nsew signal input
rlabel metal2 s 188802 0 188858 800 6 hk_dat_i[14]
port 34 nsew signal input
rlabel metal2 s 194138 0 194194 800 6 hk_dat_i[15]
port 35 nsew signal input
rlabel metal2 s 199382 0 199438 800 6 hk_dat_i[16]
port 36 nsew signal input
rlabel metal2 s 204718 0 204774 800 6 hk_dat_i[17]
port 37 nsew signal input
rlabel metal2 s 210054 0 210110 800 6 hk_dat_i[18]
port 38 nsew signal input
rlabel metal2 s 215390 0 215446 800 6 hk_dat_i[19]
port 39 nsew signal input
rlabel metal2 s 119618 0 119674 800 6 hk_dat_i[1]
port 40 nsew signal input
rlabel metal2 s 220726 0 220782 800 6 hk_dat_i[20]
port 41 nsew signal input
rlabel metal2 s 226062 0 226118 800 6 hk_dat_i[21]
port 42 nsew signal input
rlabel metal2 s 231306 0 231362 800 6 hk_dat_i[22]
port 43 nsew signal input
rlabel metal2 s 236642 0 236698 800 6 hk_dat_i[23]
port 44 nsew signal input
rlabel metal2 s 241978 0 242034 800 6 hk_dat_i[24]
port 45 nsew signal input
rlabel metal2 s 247314 0 247370 800 6 hk_dat_i[25]
port 46 nsew signal input
rlabel metal2 s 252650 0 252706 800 6 hk_dat_i[26]
port 47 nsew signal input
rlabel metal2 s 257986 0 258042 800 6 hk_dat_i[27]
port 48 nsew signal input
rlabel metal2 s 263230 0 263286 800 6 hk_dat_i[28]
port 49 nsew signal input
rlabel metal2 s 268566 0 268622 800 6 hk_dat_i[29]
port 50 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 hk_dat_i[2]
port 51 nsew signal input
rlabel metal2 s 273902 0 273958 800 6 hk_dat_i[30]
port 52 nsew signal input
rlabel metal2 s 279238 0 279294 800 6 hk_dat_i[31]
port 53 nsew signal input
rlabel metal2 s 130290 0 130346 800 6 hk_dat_i[3]
port 54 nsew signal input
rlabel metal2 s 135534 0 135590 800 6 hk_dat_i[4]
port 55 nsew signal input
rlabel metal2 s 140870 0 140926 800 6 hk_dat_i[5]
port 56 nsew signal input
rlabel metal2 s 146206 0 146262 800 6 hk_dat_i[6]
port 57 nsew signal input
rlabel metal2 s 151542 0 151598 800 6 hk_dat_i[7]
port 58 nsew signal input
rlabel metal2 s 156878 0 156934 800 6 hk_dat_i[8]
port 59 nsew signal input
rlabel metal2 s 162214 0 162270 800 6 hk_dat_i[9]
port 60 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 hk_stb_o
port 61 nsew signal tristate
rlabel metal2 s 574558 159200 574614 160000 6 irq[0]
port 62 nsew signal input
rlabel metal2 s 575570 159200 575626 160000 6 irq[1]
port 63 nsew signal input
rlabel metal2 s 576490 159200 576546 160000 6 irq[2]
port 64 nsew signal input
rlabel metal2 s 577502 159200 577558 160000 6 irq[3]
port 65 nsew signal input
rlabel metal2 s 578422 159200 578478 160000 6 irq[4]
port 66 nsew signal input
rlabel metal2 s 579434 159200 579490 160000 6 irq[5]
port 67 nsew signal input
rlabel metal2 s 2410 159200 2466 160000 6 la_iena[0]
port 68 nsew signal tristate
rlabel metal2 s 392306 159200 392362 160000 6 la_iena[100]
port 69 nsew signal tristate
rlabel metal2 s 396170 159200 396226 160000 6 la_iena[101]
port 70 nsew signal tristate
rlabel metal2 s 400034 159200 400090 160000 6 la_iena[102]
port 71 nsew signal tristate
rlabel metal2 s 403990 159200 404046 160000 6 la_iena[103]
port 72 nsew signal tristate
rlabel metal2 s 407854 159200 407910 160000 6 la_iena[104]
port 73 nsew signal tristate
rlabel metal2 s 411810 159200 411866 160000 6 la_iena[105]
port 74 nsew signal tristate
rlabel metal2 s 415674 159200 415730 160000 6 la_iena[106]
port 75 nsew signal tristate
rlabel metal2 s 419538 159200 419594 160000 6 la_iena[107]
port 76 nsew signal tristate
rlabel metal2 s 423494 159200 423550 160000 6 la_iena[108]
port 77 nsew signal tristate
rlabel metal2 s 427358 159200 427414 160000 6 la_iena[109]
port 78 nsew signal tristate
rlabel metal2 s 41326 159200 41382 160000 6 la_iena[10]
port 79 nsew signal tristate
rlabel metal2 s 431222 159200 431278 160000 6 la_iena[110]
port 80 nsew signal tristate
rlabel metal2 s 435178 159200 435234 160000 6 la_iena[111]
port 81 nsew signal tristate
rlabel metal2 s 439042 159200 439098 160000 6 la_iena[112]
port 82 nsew signal tristate
rlabel metal2 s 442998 159200 443054 160000 6 la_iena[113]
port 83 nsew signal tristate
rlabel metal2 s 446862 159200 446918 160000 6 la_iena[114]
port 84 nsew signal tristate
rlabel metal2 s 450726 159200 450782 160000 6 la_iena[115]
port 85 nsew signal tristate
rlabel metal2 s 454682 159200 454738 160000 6 la_iena[116]
port 86 nsew signal tristate
rlabel metal2 s 458546 159200 458602 160000 6 la_iena[117]
port 87 nsew signal tristate
rlabel metal2 s 462502 159200 462558 160000 6 la_iena[118]
port 88 nsew signal tristate
rlabel metal2 s 466366 159200 466422 160000 6 la_iena[119]
port 89 nsew signal tristate
rlabel metal2 s 45282 159200 45338 160000 6 la_iena[11]
port 90 nsew signal tristate
rlabel metal2 s 470230 159200 470286 160000 6 la_iena[120]
port 91 nsew signal tristate
rlabel metal2 s 474186 159200 474242 160000 6 la_iena[121]
port 92 nsew signal tristate
rlabel metal2 s 478050 159200 478106 160000 6 la_iena[122]
port 93 nsew signal tristate
rlabel metal2 s 481914 159200 481970 160000 6 la_iena[123]
port 94 nsew signal tristate
rlabel metal2 s 485870 159200 485926 160000 6 la_iena[124]
port 95 nsew signal tristate
rlabel metal2 s 489734 159200 489790 160000 6 la_iena[125]
port 96 nsew signal tristate
rlabel metal2 s 493690 159200 493746 160000 6 la_iena[126]
port 97 nsew signal tristate
rlabel metal2 s 497554 159200 497610 160000 6 la_iena[127]
port 98 nsew signal tristate
rlabel metal2 s 49146 159200 49202 160000 6 la_iena[12]
port 99 nsew signal tristate
rlabel metal2 s 53102 159200 53158 160000 6 la_iena[13]
port 100 nsew signal tristate
rlabel metal2 s 56966 159200 57022 160000 6 la_iena[14]
port 101 nsew signal tristate
rlabel metal2 s 60830 159200 60886 160000 6 la_iena[15]
port 102 nsew signal tristate
rlabel metal2 s 64786 159200 64842 160000 6 la_iena[16]
port 103 nsew signal tristate
rlabel metal2 s 68650 159200 68706 160000 6 la_iena[17]
port 104 nsew signal tristate
rlabel metal2 s 72606 159200 72662 160000 6 la_iena[18]
port 105 nsew signal tristate
rlabel metal2 s 76470 159200 76526 160000 6 la_iena[19]
port 106 nsew signal tristate
rlabel metal2 s 6274 159200 6330 160000 6 la_iena[1]
port 107 nsew signal tristate
rlabel metal2 s 80334 159200 80390 160000 6 la_iena[20]
port 108 nsew signal tristate
rlabel metal2 s 84290 159200 84346 160000 6 la_iena[21]
port 109 nsew signal tristate
rlabel metal2 s 88154 159200 88210 160000 6 la_iena[22]
port 110 nsew signal tristate
rlabel metal2 s 92018 159200 92074 160000 6 la_iena[23]
port 111 nsew signal tristate
rlabel metal2 s 95974 159200 96030 160000 6 la_iena[24]
port 112 nsew signal tristate
rlabel metal2 s 99838 159200 99894 160000 6 la_iena[25]
port 113 nsew signal tristate
rlabel metal2 s 103794 159200 103850 160000 6 la_iena[26]
port 114 nsew signal tristate
rlabel metal2 s 107658 159200 107714 160000 6 la_iena[27]
port 115 nsew signal tristate
rlabel metal2 s 111522 159200 111578 160000 6 la_iena[28]
port 116 nsew signal tristate
rlabel metal2 s 115478 159200 115534 160000 6 la_iena[29]
port 117 nsew signal tristate
rlabel metal2 s 10138 159200 10194 160000 6 la_iena[2]
port 118 nsew signal tristate
rlabel metal2 s 119342 159200 119398 160000 6 la_iena[30]
port 119 nsew signal tristate
rlabel metal2 s 123206 159200 123262 160000 6 la_iena[31]
port 120 nsew signal tristate
rlabel metal2 s 127162 159200 127218 160000 6 la_iena[32]
port 121 nsew signal tristate
rlabel metal2 s 131026 159200 131082 160000 6 la_iena[33]
port 122 nsew signal tristate
rlabel metal2 s 134982 159200 135038 160000 6 la_iena[34]
port 123 nsew signal tristate
rlabel metal2 s 138846 159200 138902 160000 6 la_iena[35]
port 124 nsew signal tristate
rlabel metal2 s 142710 159200 142766 160000 6 la_iena[36]
port 125 nsew signal tristate
rlabel metal2 s 146666 159200 146722 160000 6 la_iena[37]
port 126 nsew signal tristate
rlabel metal2 s 150530 159200 150586 160000 6 la_iena[38]
port 127 nsew signal tristate
rlabel metal2 s 154486 159200 154542 160000 6 la_iena[39]
port 128 nsew signal tristate
rlabel metal2 s 14094 159200 14150 160000 6 la_iena[3]
port 129 nsew signal tristate
rlabel metal2 s 158350 159200 158406 160000 6 la_iena[40]
port 130 nsew signal tristate
rlabel metal2 s 162214 159200 162270 160000 6 la_iena[41]
port 131 nsew signal tristate
rlabel metal2 s 166170 159200 166226 160000 6 la_iena[42]
port 132 nsew signal tristate
rlabel metal2 s 170034 159200 170090 160000 6 la_iena[43]
port 133 nsew signal tristate
rlabel metal2 s 173898 159200 173954 160000 6 la_iena[44]
port 134 nsew signal tristate
rlabel metal2 s 177854 159200 177910 160000 6 la_iena[45]
port 135 nsew signal tristate
rlabel metal2 s 181718 159200 181774 160000 6 la_iena[46]
port 136 nsew signal tristate
rlabel metal2 s 185674 159200 185730 160000 6 la_iena[47]
port 137 nsew signal tristate
rlabel metal2 s 189538 159200 189594 160000 6 la_iena[48]
port 138 nsew signal tristate
rlabel metal2 s 193402 159200 193458 160000 6 la_iena[49]
port 139 nsew signal tristate
rlabel metal2 s 17958 159200 18014 160000 6 la_iena[4]
port 140 nsew signal tristate
rlabel metal2 s 197358 159200 197414 160000 6 la_iena[50]
port 141 nsew signal tristate
rlabel metal2 s 201222 159200 201278 160000 6 la_iena[51]
port 142 nsew signal tristate
rlabel metal2 s 205086 159200 205142 160000 6 la_iena[52]
port 143 nsew signal tristate
rlabel metal2 s 209042 159200 209098 160000 6 la_iena[53]
port 144 nsew signal tristate
rlabel metal2 s 212906 159200 212962 160000 6 la_iena[54]
port 145 nsew signal tristate
rlabel metal2 s 216862 159200 216918 160000 6 la_iena[55]
port 146 nsew signal tristate
rlabel metal2 s 220726 159200 220782 160000 6 la_iena[56]
port 147 nsew signal tristate
rlabel metal2 s 224590 159200 224646 160000 6 la_iena[57]
port 148 nsew signal tristate
rlabel metal2 s 228546 159200 228602 160000 6 la_iena[58]
port 149 nsew signal tristate
rlabel metal2 s 232410 159200 232466 160000 6 la_iena[59]
port 150 nsew signal tristate
rlabel metal2 s 21914 159200 21970 160000 6 la_iena[5]
port 151 nsew signal tristate
rlabel metal2 s 236274 159200 236330 160000 6 la_iena[60]
port 152 nsew signal tristate
rlabel metal2 s 240230 159200 240286 160000 6 la_iena[61]
port 153 nsew signal tristate
rlabel metal2 s 244094 159200 244150 160000 6 la_iena[62]
port 154 nsew signal tristate
rlabel metal2 s 248050 159200 248106 160000 6 la_iena[63]
port 155 nsew signal tristate
rlabel metal2 s 251914 159200 251970 160000 6 la_iena[64]
port 156 nsew signal tristate
rlabel metal2 s 255778 159200 255834 160000 6 la_iena[65]
port 157 nsew signal tristate
rlabel metal2 s 259734 159200 259790 160000 6 la_iena[66]
port 158 nsew signal tristate
rlabel metal2 s 263598 159200 263654 160000 6 la_iena[67]
port 159 nsew signal tristate
rlabel metal2 s 267554 159200 267610 160000 6 la_iena[68]
port 160 nsew signal tristate
rlabel metal2 s 271418 159200 271474 160000 6 la_iena[69]
port 161 nsew signal tristate
rlabel metal2 s 25778 159200 25834 160000 6 la_iena[6]
port 162 nsew signal tristate
rlabel metal2 s 275282 159200 275338 160000 6 la_iena[70]
port 163 nsew signal tristate
rlabel metal2 s 279238 159200 279294 160000 6 la_iena[71]
port 164 nsew signal tristate
rlabel metal2 s 283102 159200 283158 160000 6 la_iena[72]
port 165 nsew signal tristate
rlabel metal2 s 286966 159200 287022 160000 6 la_iena[73]
port 166 nsew signal tristate
rlabel metal2 s 290922 159200 290978 160000 6 la_iena[74]
port 167 nsew signal tristate
rlabel metal2 s 294786 159200 294842 160000 6 la_iena[75]
port 168 nsew signal tristate
rlabel metal2 s 298742 159200 298798 160000 6 la_iena[76]
port 169 nsew signal tristate
rlabel metal2 s 302606 159200 302662 160000 6 la_iena[77]
port 170 nsew signal tristate
rlabel metal2 s 306470 159200 306526 160000 6 la_iena[78]
port 171 nsew signal tristate
rlabel metal2 s 310426 159200 310482 160000 6 la_iena[79]
port 172 nsew signal tristate
rlabel metal2 s 29642 159200 29698 160000 6 la_iena[7]
port 173 nsew signal tristate
rlabel metal2 s 314290 159200 314346 160000 6 la_iena[80]
port 174 nsew signal tristate
rlabel metal2 s 318154 159200 318210 160000 6 la_iena[81]
port 175 nsew signal tristate
rlabel metal2 s 322110 159200 322166 160000 6 la_iena[82]
port 176 nsew signal tristate
rlabel metal2 s 325974 159200 326030 160000 6 la_iena[83]
port 177 nsew signal tristate
rlabel metal2 s 329930 159200 329986 160000 6 la_iena[84]
port 178 nsew signal tristate
rlabel metal2 s 333794 159200 333850 160000 6 la_iena[85]
port 179 nsew signal tristate
rlabel metal2 s 337658 159200 337714 160000 6 la_iena[86]
port 180 nsew signal tristate
rlabel metal2 s 341614 159200 341670 160000 6 la_iena[87]
port 181 nsew signal tristate
rlabel metal2 s 345478 159200 345534 160000 6 la_iena[88]
port 182 nsew signal tristate
rlabel metal2 s 349342 159200 349398 160000 6 la_iena[89]
port 183 nsew signal tristate
rlabel metal2 s 33598 159200 33654 160000 6 la_iena[8]
port 184 nsew signal tristate
rlabel metal2 s 353298 159200 353354 160000 6 la_iena[90]
port 185 nsew signal tristate
rlabel metal2 s 357162 159200 357218 160000 6 la_iena[91]
port 186 nsew signal tristate
rlabel metal2 s 361118 159200 361174 160000 6 la_iena[92]
port 187 nsew signal tristate
rlabel metal2 s 364982 159200 365038 160000 6 la_iena[93]
port 188 nsew signal tristate
rlabel metal2 s 368846 159200 368902 160000 6 la_iena[94]
port 189 nsew signal tristate
rlabel metal2 s 372802 159200 372858 160000 6 la_iena[95]
port 190 nsew signal tristate
rlabel metal2 s 376666 159200 376722 160000 6 la_iena[96]
port 191 nsew signal tristate
rlabel metal2 s 380622 159200 380678 160000 6 la_iena[97]
port 192 nsew signal tristate
rlabel metal2 s 384486 159200 384542 160000 6 la_iena[98]
port 193 nsew signal tristate
rlabel metal2 s 388350 159200 388406 160000 6 la_iena[99]
port 194 nsew signal tristate
rlabel metal2 s 37462 159200 37518 160000 6 la_iena[9]
port 195 nsew signal tristate
rlabel metal2 s 3330 159200 3386 160000 6 la_input[0]
port 196 nsew signal input
rlabel metal2 s 393226 159200 393282 160000 6 la_input[100]
port 197 nsew signal input
rlabel metal2 s 397182 159200 397238 160000 6 la_input[101]
port 198 nsew signal input
rlabel metal2 s 401046 159200 401102 160000 6 la_input[102]
port 199 nsew signal input
rlabel metal2 s 404910 159200 404966 160000 6 la_input[103]
port 200 nsew signal input
rlabel metal2 s 408866 159200 408922 160000 6 la_input[104]
port 201 nsew signal input
rlabel metal2 s 412730 159200 412786 160000 6 la_input[105]
port 202 nsew signal input
rlabel metal2 s 416686 159200 416742 160000 6 la_input[106]
port 203 nsew signal input
rlabel metal2 s 420550 159200 420606 160000 6 la_input[107]
port 204 nsew signal input
rlabel metal2 s 424414 159200 424470 160000 6 la_input[108]
port 205 nsew signal input
rlabel metal2 s 428370 159200 428426 160000 6 la_input[109]
port 206 nsew signal input
rlabel metal2 s 42338 159200 42394 160000 6 la_input[10]
port 207 nsew signal input
rlabel metal2 s 432234 159200 432290 160000 6 la_input[110]
port 208 nsew signal input
rlabel metal2 s 436098 159200 436154 160000 6 la_input[111]
port 209 nsew signal input
rlabel metal2 s 440054 159200 440110 160000 6 la_input[112]
port 210 nsew signal input
rlabel metal2 s 443918 159200 443974 160000 6 la_input[113]
port 211 nsew signal input
rlabel metal2 s 447874 159200 447930 160000 6 la_input[114]
port 212 nsew signal input
rlabel metal2 s 451738 159200 451794 160000 6 la_input[115]
port 213 nsew signal input
rlabel metal2 s 455602 159200 455658 160000 6 la_input[116]
port 214 nsew signal input
rlabel metal2 s 459558 159200 459614 160000 6 la_input[117]
port 215 nsew signal input
rlabel metal2 s 463422 159200 463478 160000 6 la_input[118]
port 216 nsew signal input
rlabel metal2 s 467286 159200 467342 160000 6 la_input[119]
port 217 nsew signal input
rlabel metal2 s 46202 159200 46258 160000 6 la_input[11]
port 218 nsew signal input
rlabel metal2 s 471242 159200 471298 160000 6 la_input[120]
port 219 nsew signal input
rlabel metal2 s 475106 159200 475162 160000 6 la_input[121]
port 220 nsew signal input
rlabel metal2 s 479062 159200 479118 160000 6 la_input[122]
port 221 nsew signal input
rlabel metal2 s 482926 159200 482982 160000 6 la_input[123]
port 222 nsew signal input
rlabel metal2 s 486790 159200 486846 160000 6 la_input[124]
port 223 nsew signal input
rlabel metal2 s 490746 159200 490802 160000 6 la_input[125]
port 224 nsew signal input
rlabel metal2 s 494610 159200 494666 160000 6 la_input[126]
port 225 nsew signal input
rlabel metal2 s 498566 159200 498622 160000 6 la_input[127]
port 226 nsew signal input
rlabel metal2 s 50158 159200 50214 160000 6 la_input[12]
port 227 nsew signal input
rlabel metal2 s 54022 159200 54078 160000 6 la_input[13]
port 228 nsew signal input
rlabel metal2 s 57978 159200 58034 160000 6 la_input[14]
port 229 nsew signal input
rlabel metal2 s 61842 159200 61898 160000 6 la_input[15]
port 230 nsew signal input
rlabel metal2 s 65706 159200 65762 160000 6 la_input[16]
port 231 nsew signal input
rlabel metal2 s 69662 159200 69718 160000 6 la_input[17]
port 232 nsew signal input
rlabel metal2 s 73526 159200 73582 160000 6 la_input[18]
port 233 nsew signal input
rlabel metal2 s 77482 159200 77538 160000 6 la_input[19]
port 234 nsew signal input
rlabel metal2 s 7286 159200 7342 160000 6 la_input[1]
port 235 nsew signal input
rlabel metal2 s 81346 159200 81402 160000 6 la_input[20]
port 236 nsew signal input
rlabel metal2 s 85210 159200 85266 160000 6 la_input[21]
port 237 nsew signal input
rlabel metal2 s 89166 159200 89222 160000 6 la_input[22]
port 238 nsew signal input
rlabel metal2 s 93030 159200 93086 160000 6 la_input[23]
port 239 nsew signal input
rlabel metal2 s 96894 159200 96950 160000 6 la_input[24]
port 240 nsew signal input
rlabel metal2 s 100850 159200 100906 160000 6 la_input[25]
port 241 nsew signal input
rlabel metal2 s 104714 159200 104770 160000 6 la_input[26]
port 242 nsew signal input
rlabel metal2 s 108670 159200 108726 160000 6 la_input[27]
port 243 nsew signal input
rlabel metal2 s 112534 159200 112590 160000 6 la_input[28]
port 244 nsew signal input
rlabel metal2 s 116398 159200 116454 160000 6 la_input[29]
port 245 nsew signal input
rlabel metal2 s 11150 159200 11206 160000 6 la_input[2]
port 246 nsew signal input
rlabel metal2 s 120354 159200 120410 160000 6 la_input[30]
port 247 nsew signal input
rlabel metal2 s 124218 159200 124274 160000 6 la_input[31]
port 248 nsew signal input
rlabel metal2 s 128082 159200 128138 160000 6 la_input[32]
port 249 nsew signal input
rlabel metal2 s 132038 159200 132094 160000 6 la_input[33]
port 250 nsew signal input
rlabel metal2 s 135902 159200 135958 160000 6 la_input[34]
port 251 nsew signal input
rlabel metal2 s 139858 159200 139914 160000 6 la_input[35]
port 252 nsew signal input
rlabel metal2 s 143722 159200 143778 160000 6 la_input[36]
port 253 nsew signal input
rlabel metal2 s 147586 159200 147642 160000 6 la_input[37]
port 254 nsew signal input
rlabel metal2 s 151542 159200 151598 160000 6 la_input[38]
port 255 nsew signal input
rlabel metal2 s 155406 159200 155462 160000 6 la_input[39]
port 256 nsew signal input
rlabel metal2 s 15014 159200 15070 160000 6 la_input[3]
port 257 nsew signal input
rlabel metal2 s 159270 159200 159326 160000 6 la_input[40]
port 258 nsew signal input
rlabel metal2 s 163226 159200 163282 160000 6 la_input[41]
port 259 nsew signal input
rlabel metal2 s 167090 159200 167146 160000 6 la_input[42]
port 260 nsew signal input
rlabel metal2 s 171046 159200 171102 160000 6 la_input[43]
port 261 nsew signal input
rlabel metal2 s 174910 159200 174966 160000 6 la_input[44]
port 262 nsew signal input
rlabel metal2 s 178774 159200 178830 160000 6 la_input[45]
port 263 nsew signal input
rlabel metal2 s 182730 159200 182786 160000 6 la_input[46]
port 264 nsew signal input
rlabel metal2 s 186594 159200 186650 160000 6 la_input[47]
port 265 nsew signal input
rlabel metal2 s 190550 159200 190606 160000 6 la_input[48]
port 266 nsew signal input
rlabel metal2 s 194414 159200 194470 160000 6 la_input[49]
port 267 nsew signal input
rlabel metal2 s 18970 159200 19026 160000 6 la_input[4]
port 268 nsew signal input
rlabel metal2 s 198278 159200 198334 160000 6 la_input[50]
port 269 nsew signal input
rlabel metal2 s 202234 159200 202290 160000 6 la_input[51]
port 270 nsew signal input
rlabel metal2 s 206098 159200 206154 160000 6 la_input[52]
port 271 nsew signal input
rlabel metal2 s 209962 159200 210018 160000 6 la_input[53]
port 272 nsew signal input
rlabel metal2 s 213918 159200 213974 160000 6 la_input[54]
port 273 nsew signal input
rlabel metal2 s 217782 159200 217838 160000 6 la_input[55]
port 274 nsew signal input
rlabel metal2 s 221738 159200 221794 160000 6 la_input[56]
port 275 nsew signal input
rlabel metal2 s 225602 159200 225658 160000 6 la_input[57]
port 276 nsew signal input
rlabel metal2 s 229466 159200 229522 160000 6 la_input[58]
port 277 nsew signal input
rlabel metal2 s 233422 159200 233478 160000 6 la_input[59]
port 278 nsew signal input
rlabel metal2 s 22834 159200 22890 160000 6 la_input[5]
port 279 nsew signal input
rlabel metal2 s 237286 159200 237342 160000 6 la_input[60]
port 280 nsew signal input
rlabel metal2 s 241150 159200 241206 160000 6 la_input[61]
port 281 nsew signal input
rlabel metal2 s 245106 159200 245162 160000 6 la_input[62]
port 282 nsew signal input
rlabel metal2 s 248970 159200 249026 160000 6 la_input[63]
port 283 nsew signal input
rlabel metal2 s 252926 159200 252982 160000 6 la_input[64]
port 284 nsew signal input
rlabel metal2 s 256790 159200 256846 160000 6 la_input[65]
port 285 nsew signal input
rlabel metal2 s 260654 159200 260710 160000 6 la_input[66]
port 286 nsew signal input
rlabel metal2 s 264610 159200 264666 160000 6 la_input[67]
port 287 nsew signal input
rlabel metal2 s 268474 159200 268530 160000 6 la_input[68]
port 288 nsew signal input
rlabel metal2 s 272338 159200 272394 160000 6 la_input[69]
port 289 nsew signal input
rlabel metal2 s 26790 159200 26846 160000 6 la_input[6]
port 290 nsew signal input
rlabel metal2 s 276294 159200 276350 160000 6 la_input[70]
port 291 nsew signal input
rlabel metal2 s 280158 159200 280214 160000 6 la_input[71]
port 292 nsew signal input
rlabel metal2 s 284114 159200 284170 160000 6 la_input[72]
port 293 nsew signal input
rlabel metal2 s 287978 159200 288034 160000 6 la_input[73]
port 294 nsew signal input
rlabel metal2 s 291842 159200 291898 160000 6 la_input[74]
port 295 nsew signal input
rlabel metal2 s 295798 159200 295854 160000 6 la_input[75]
port 296 nsew signal input
rlabel metal2 s 299662 159200 299718 160000 6 la_input[76]
port 297 nsew signal input
rlabel metal2 s 303618 159200 303674 160000 6 la_input[77]
port 298 nsew signal input
rlabel metal2 s 307482 159200 307538 160000 6 la_input[78]
port 299 nsew signal input
rlabel metal2 s 311346 159200 311402 160000 6 la_input[79]
port 300 nsew signal input
rlabel metal2 s 30654 159200 30710 160000 6 la_input[7]
port 301 nsew signal input
rlabel metal2 s 315302 159200 315358 160000 6 la_input[80]
port 302 nsew signal input
rlabel metal2 s 319166 159200 319222 160000 6 la_input[81]
port 303 nsew signal input
rlabel metal2 s 323030 159200 323086 160000 6 la_input[82]
port 304 nsew signal input
rlabel metal2 s 326986 159200 327042 160000 6 la_input[83]
port 305 nsew signal input
rlabel metal2 s 330850 159200 330906 160000 6 la_input[84]
port 306 nsew signal input
rlabel metal2 s 334806 159200 334862 160000 6 la_input[85]
port 307 nsew signal input
rlabel metal2 s 338670 159200 338726 160000 6 la_input[86]
port 308 nsew signal input
rlabel metal2 s 342534 159200 342590 160000 6 la_input[87]
port 309 nsew signal input
rlabel metal2 s 346490 159200 346546 160000 6 la_input[88]
port 310 nsew signal input
rlabel metal2 s 350354 159200 350410 160000 6 la_input[89]
port 311 nsew signal input
rlabel metal2 s 34518 159200 34574 160000 6 la_input[8]
port 312 nsew signal input
rlabel metal2 s 354218 159200 354274 160000 6 la_input[90]
port 313 nsew signal input
rlabel metal2 s 358174 159200 358230 160000 6 la_input[91]
port 314 nsew signal input
rlabel metal2 s 362038 159200 362094 160000 6 la_input[92]
port 315 nsew signal input
rlabel metal2 s 365994 159200 366050 160000 6 la_input[93]
port 316 nsew signal input
rlabel metal2 s 369858 159200 369914 160000 6 la_input[94]
port 317 nsew signal input
rlabel metal2 s 373722 159200 373778 160000 6 la_input[95]
port 318 nsew signal input
rlabel metal2 s 377678 159200 377734 160000 6 la_input[96]
port 319 nsew signal input
rlabel metal2 s 381542 159200 381598 160000 6 la_input[97]
port 320 nsew signal input
rlabel metal2 s 385498 159200 385554 160000 6 la_input[98]
port 321 nsew signal input
rlabel metal2 s 389362 159200 389418 160000 6 la_input[99]
port 322 nsew signal input
rlabel metal2 s 38474 159200 38530 160000 6 la_input[9]
port 323 nsew signal input
rlabel metal2 s 4342 159200 4398 160000 6 la_oenb[0]
port 324 nsew signal tristate
rlabel metal2 s 394238 159200 394294 160000 6 la_oenb[100]
port 325 nsew signal tristate
rlabel metal2 s 398102 159200 398158 160000 6 la_oenb[101]
port 326 nsew signal tristate
rlabel metal2 s 402058 159200 402114 160000 6 la_oenb[102]
port 327 nsew signal tristate
rlabel metal2 s 405922 159200 405978 160000 6 la_oenb[103]
port 328 nsew signal tristate
rlabel metal2 s 409786 159200 409842 160000 6 la_oenb[104]
port 329 nsew signal tristate
rlabel metal2 s 413742 159200 413798 160000 6 la_oenb[105]
port 330 nsew signal tristate
rlabel metal2 s 417606 159200 417662 160000 6 la_oenb[106]
port 331 nsew signal tristate
rlabel metal2 s 421562 159200 421618 160000 6 la_oenb[107]
port 332 nsew signal tristate
rlabel metal2 s 425426 159200 425482 160000 6 la_oenb[108]
port 333 nsew signal tristate
rlabel metal2 s 429290 159200 429346 160000 6 la_oenb[109]
port 334 nsew signal tristate
rlabel metal2 s 43350 159200 43406 160000 6 la_oenb[10]
port 335 nsew signal tristate
rlabel metal2 s 433246 159200 433302 160000 6 la_oenb[110]
port 336 nsew signal tristate
rlabel metal2 s 437110 159200 437166 160000 6 la_oenb[111]
port 337 nsew signal tristate
rlabel metal2 s 440974 159200 441030 160000 6 la_oenb[112]
port 338 nsew signal tristate
rlabel metal2 s 444930 159200 444986 160000 6 la_oenb[113]
port 339 nsew signal tristate
rlabel metal2 s 448794 159200 448850 160000 6 la_oenb[114]
port 340 nsew signal tristate
rlabel metal2 s 452750 159200 452806 160000 6 la_oenb[115]
port 341 nsew signal tristate
rlabel metal2 s 456614 159200 456670 160000 6 la_oenb[116]
port 342 nsew signal tristate
rlabel metal2 s 460478 159200 460534 160000 6 la_oenb[117]
port 343 nsew signal tristate
rlabel metal2 s 464434 159200 464490 160000 6 la_oenb[118]
port 344 nsew signal tristate
rlabel metal2 s 468298 159200 468354 160000 6 la_oenb[119]
port 345 nsew signal tristate
rlabel metal2 s 47214 159200 47270 160000 6 la_oenb[11]
port 346 nsew signal tristate
rlabel metal2 s 472162 159200 472218 160000 6 la_oenb[120]
port 347 nsew signal tristate
rlabel metal2 s 476118 159200 476174 160000 6 la_oenb[121]
port 348 nsew signal tristate
rlabel metal2 s 479982 159200 480038 160000 6 la_oenb[122]
port 349 nsew signal tristate
rlabel metal2 s 483938 159200 483994 160000 6 la_oenb[123]
port 350 nsew signal tristate
rlabel metal2 s 487802 159200 487858 160000 6 la_oenb[124]
port 351 nsew signal tristate
rlabel metal2 s 491666 159200 491722 160000 6 la_oenb[125]
port 352 nsew signal tristate
rlabel metal2 s 495622 159200 495678 160000 6 la_oenb[126]
port 353 nsew signal tristate
rlabel metal2 s 499486 159200 499542 160000 6 la_oenb[127]
port 354 nsew signal tristate
rlabel metal2 s 51078 159200 51134 160000 6 la_oenb[12]
port 355 nsew signal tristate
rlabel metal2 s 55034 159200 55090 160000 6 la_oenb[13]
port 356 nsew signal tristate
rlabel metal2 s 58898 159200 58954 160000 6 la_oenb[14]
port 357 nsew signal tristate
rlabel metal2 s 62854 159200 62910 160000 6 la_oenb[15]
port 358 nsew signal tristate
rlabel metal2 s 66718 159200 66774 160000 6 la_oenb[16]
port 359 nsew signal tristate
rlabel metal2 s 70582 159200 70638 160000 6 la_oenb[17]
port 360 nsew signal tristate
rlabel metal2 s 74538 159200 74594 160000 6 la_oenb[18]
port 361 nsew signal tristate
rlabel metal2 s 78402 159200 78458 160000 6 la_oenb[19]
port 362 nsew signal tristate
rlabel metal2 s 8206 159200 8262 160000 6 la_oenb[1]
port 363 nsew signal tristate
rlabel metal2 s 82266 159200 82322 160000 6 la_oenb[20]
port 364 nsew signal tristate
rlabel metal2 s 86222 159200 86278 160000 6 la_oenb[21]
port 365 nsew signal tristate
rlabel metal2 s 90086 159200 90142 160000 6 la_oenb[22]
port 366 nsew signal tristate
rlabel metal2 s 94042 159200 94098 160000 6 la_oenb[23]
port 367 nsew signal tristate
rlabel metal2 s 97906 159200 97962 160000 6 la_oenb[24]
port 368 nsew signal tristate
rlabel metal2 s 101770 159200 101826 160000 6 la_oenb[25]
port 369 nsew signal tristate
rlabel metal2 s 105726 159200 105782 160000 6 la_oenb[26]
port 370 nsew signal tristate
rlabel metal2 s 109590 159200 109646 160000 6 la_oenb[27]
port 371 nsew signal tristate
rlabel metal2 s 113546 159200 113602 160000 6 la_oenb[28]
port 372 nsew signal tristate
rlabel metal2 s 117410 159200 117466 160000 6 la_oenb[29]
port 373 nsew signal tristate
rlabel metal2 s 12162 159200 12218 160000 6 la_oenb[2]
port 374 nsew signal tristate
rlabel metal2 s 121274 159200 121330 160000 6 la_oenb[30]
port 375 nsew signal tristate
rlabel metal2 s 125230 159200 125286 160000 6 la_oenb[31]
port 376 nsew signal tristate
rlabel metal2 s 129094 159200 129150 160000 6 la_oenb[32]
port 377 nsew signal tristate
rlabel metal2 s 132958 159200 133014 160000 6 la_oenb[33]
port 378 nsew signal tristate
rlabel metal2 s 136914 159200 136970 160000 6 la_oenb[34]
port 379 nsew signal tristate
rlabel metal2 s 140778 159200 140834 160000 6 la_oenb[35]
port 380 nsew signal tristate
rlabel metal2 s 144734 159200 144790 160000 6 la_oenb[36]
port 381 nsew signal tristate
rlabel metal2 s 148598 159200 148654 160000 6 la_oenb[37]
port 382 nsew signal tristate
rlabel metal2 s 152462 159200 152518 160000 6 la_oenb[38]
port 383 nsew signal tristate
rlabel metal2 s 156418 159200 156474 160000 6 la_oenb[39]
port 384 nsew signal tristate
rlabel metal2 s 16026 159200 16082 160000 6 la_oenb[3]
port 385 nsew signal tristate
rlabel metal2 s 160282 159200 160338 160000 6 la_oenb[40]
port 386 nsew signal tristate
rlabel metal2 s 164146 159200 164202 160000 6 la_oenb[41]
port 387 nsew signal tristate
rlabel metal2 s 168102 159200 168158 160000 6 la_oenb[42]
port 388 nsew signal tristate
rlabel metal2 s 171966 159200 172022 160000 6 la_oenb[43]
port 389 nsew signal tristate
rlabel metal2 s 175922 159200 175978 160000 6 la_oenb[44]
port 390 nsew signal tristate
rlabel metal2 s 179786 159200 179842 160000 6 la_oenb[45]
port 391 nsew signal tristate
rlabel metal2 s 183650 159200 183706 160000 6 la_oenb[46]
port 392 nsew signal tristate
rlabel metal2 s 187606 159200 187662 160000 6 la_oenb[47]
port 393 nsew signal tristate
rlabel metal2 s 191470 159200 191526 160000 6 la_oenb[48]
port 394 nsew signal tristate
rlabel metal2 s 195334 159200 195390 160000 6 la_oenb[49]
port 395 nsew signal tristate
rlabel metal2 s 19890 159200 19946 160000 6 la_oenb[4]
port 396 nsew signal tristate
rlabel metal2 s 199290 159200 199346 160000 6 la_oenb[50]
port 397 nsew signal tristate
rlabel metal2 s 203154 159200 203210 160000 6 la_oenb[51]
port 398 nsew signal tristate
rlabel metal2 s 207110 159200 207166 160000 6 la_oenb[52]
port 399 nsew signal tristate
rlabel metal2 s 210974 159200 211030 160000 6 la_oenb[53]
port 400 nsew signal tristate
rlabel metal2 s 214838 159200 214894 160000 6 la_oenb[54]
port 401 nsew signal tristate
rlabel metal2 s 218794 159200 218850 160000 6 la_oenb[55]
port 402 nsew signal tristate
rlabel metal2 s 222658 159200 222714 160000 6 la_oenb[56]
port 403 nsew signal tristate
rlabel metal2 s 226614 159200 226670 160000 6 la_oenb[57]
port 404 nsew signal tristate
rlabel metal2 s 230478 159200 230534 160000 6 la_oenb[58]
port 405 nsew signal tristate
rlabel metal2 s 234342 159200 234398 160000 6 la_oenb[59]
port 406 nsew signal tristate
rlabel metal2 s 23846 159200 23902 160000 6 la_oenb[5]
port 407 nsew signal tristate
rlabel metal2 s 238298 159200 238354 160000 6 la_oenb[60]
port 408 nsew signal tristate
rlabel metal2 s 242162 159200 242218 160000 6 la_oenb[61]
port 409 nsew signal tristate
rlabel metal2 s 246026 159200 246082 160000 6 la_oenb[62]
port 410 nsew signal tristate
rlabel metal2 s 249982 159200 250038 160000 6 la_oenb[63]
port 411 nsew signal tristate
rlabel metal2 s 253846 159200 253902 160000 6 la_oenb[64]
port 412 nsew signal tristate
rlabel metal2 s 257802 159200 257858 160000 6 la_oenb[65]
port 413 nsew signal tristate
rlabel metal2 s 261666 159200 261722 160000 6 la_oenb[66]
port 414 nsew signal tristate
rlabel metal2 s 265530 159200 265586 160000 6 la_oenb[67]
port 415 nsew signal tristate
rlabel metal2 s 269486 159200 269542 160000 6 la_oenb[68]
port 416 nsew signal tristate
rlabel metal2 s 273350 159200 273406 160000 6 la_oenb[69]
port 417 nsew signal tristate
rlabel metal2 s 27710 159200 27766 160000 6 la_oenb[6]
port 418 nsew signal tristate
rlabel metal2 s 277214 159200 277270 160000 6 la_oenb[70]
port 419 nsew signal tristate
rlabel metal2 s 281170 159200 281226 160000 6 la_oenb[71]
port 420 nsew signal tristate
rlabel metal2 s 285034 159200 285090 160000 6 la_oenb[72]
port 421 nsew signal tristate
rlabel metal2 s 288990 159200 289046 160000 6 la_oenb[73]
port 422 nsew signal tristate
rlabel metal2 s 292854 159200 292910 160000 6 la_oenb[74]
port 423 nsew signal tristate
rlabel metal2 s 296718 159200 296774 160000 6 la_oenb[75]
port 424 nsew signal tristate
rlabel metal2 s 300674 159200 300730 160000 6 la_oenb[76]
port 425 nsew signal tristate
rlabel metal2 s 304538 159200 304594 160000 6 la_oenb[77]
port 426 nsew signal tristate
rlabel metal2 s 308494 159200 308550 160000 6 la_oenb[78]
port 427 nsew signal tristate
rlabel metal2 s 312358 159200 312414 160000 6 la_oenb[79]
port 428 nsew signal tristate
rlabel metal2 s 31666 159200 31722 160000 6 la_oenb[7]
port 429 nsew signal tristate
rlabel metal2 s 316222 159200 316278 160000 6 la_oenb[80]
port 430 nsew signal tristate
rlabel metal2 s 320178 159200 320234 160000 6 la_oenb[81]
port 431 nsew signal tristate
rlabel metal2 s 324042 159200 324098 160000 6 la_oenb[82]
port 432 nsew signal tristate
rlabel metal2 s 327906 159200 327962 160000 6 la_oenb[83]
port 433 nsew signal tristate
rlabel metal2 s 331862 159200 331918 160000 6 la_oenb[84]
port 434 nsew signal tristate
rlabel metal2 s 335726 159200 335782 160000 6 la_oenb[85]
port 435 nsew signal tristate
rlabel metal2 s 339682 159200 339738 160000 6 la_oenb[86]
port 436 nsew signal tristate
rlabel metal2 s 343546 159200 343602 160000 6 la_oenb[87]
port 437 nsew signal tristate
rlabel metal2 s 347410 159200 347466 160000 6 la_oenb[88]
port 438 nsew signal tristate
rlabel metal2 s 351366 159200 351422 160000 6 la_oenb[89]
port 439 nsew signal tristate
rlabel metal2 s 35530 159200 35586 160000 6 la_oenb[8]
port 440 nsew signal tristate
rlabel metal2 s 355230 159200 355286 160000 6 la_oenb[90]
port 441 nsew signal tristate
rlabel metal2 s 359094 159200 359150 160000 6 la_oenb[91]
port 442 nsew signal tristate
rlabel metal2 s 363050 159200 363106 160000 6 la_oenb[92]
port 443 nsew signal tristate
rlabel metal2 s 366914 159200 366970 160000 6 la_oenb[93]
port 444 nsew signal tristate
rlabel metal2 s 370870 159200 370926 160000 6 la_oenb[94]
port 445 nsew signal tristate
rlabel metal2 s 374734 159200 374790 160000 6 la_oenb[95]
port 446 nsew signal tristate
rlabel metal2 s 378598 159200 378654 160000 6 la_oenb[96]
port 447 nsew signal tristate
rlabel metal2 s 382554 159200 382610 160000 6 la_oenb[97]
port 448 nsew signal tristate
rlabel metal2 s 386418 159200 386474 160000 6 la_oenb[98]
port 449 nsew signal tristate
rlabel metal2 s 390282 159200 390338 160000 6 la_oenb[99]
port 450 nsew signal tristate
rlabel metal2 s 39394 159200 39450 160000 6 la_oenb[9]
port 451 nsew signal tristate
rlabel metal2 s 5262 159200 5318 160000 6 la_output[0]
port 452 nsew signal tristate
rlabel metal2 s 395158 159200 395214 160000 6 la_output[100]
port 453 nsew signal tristate
rlabel metal2 s 399114 159200 399170 160000 6 la_output[101]
port 454 nsew signal tristate
rlabel metal2 s 402978 159200 403034 160000 6 la_output[102]
port 455 nsew signal tristate
rlabel metal2 s 406934 159200 406990 160000 6 la_output[103]
port 456 nsew signal tristate
rlabel metal2 s 410798 159200 410854 160000 6 la_output[104]
port 457 nsew signal tristate
rlabel metal2 s 414662 159200 414718 160000 6 la_output[105]
port 458 nsew signal tristate
rlabel metal2 s 418618 159200 418674 160000 6 la_output[106]
port 459 nsew signal tristate
rlabel metal2 s 422482 159200 422538 160000 6 la_output[107]
port 460 nsew signal tristate
rlabel metal2 s 426346 159200 426402 160000 6 la_output[108]
port 461 nsew signal tristate
rlabel metal2 s 430302 159200 430358 160000 6 la_output[109]
port 462 nsew signal tristate
rlabel metal2 s 44270 159200 44326 160000 6 la_output[10]
port 463 nsew signal tristate
rlabel metal2 s 434166 159200 434222 160000 6 la_output[110]
port 464 nsew signal tristate
rlabel metal2 s 438122 159200 438178 160000 6 la_output[111]
port 465 nsew signal tristate
rlabel metal2 s 441986 159200 442042 160000 6 la_output[112]
port 466 nsew signal tristate
rlabel metal2 s 445850 159200 445906 160000 6 la_output[113]
port 467 nsew signal tristate
rlabel metal2 s 449806 159200 449862 160000 6 la_output[114]
port 468 nsew signal tristate
rlabel metal2 s 453670 159200 453726 160000 6 la_output[115]
port 469 nsew signal tristate
rlabel metal2 s 457626 159200 457682 160000 6 la_output[116]
port 470 nsew signal tristate
rlabel metal2 s 461490 159200 461546 160000 6 la_output[117]
port 471 nsew signal tristate
rlabel metal2 s 465354 159200 465410 160000 6 la_output[118]
port 472 nsew signal tristate
rlabel metal2 s 469310 159200 469366 160000 6 la_output[119]
port 473 nsew signal tristate
rlabel metal2 s 48226 159200 48282 160000 6 la_output[11]
port 474 nsew signal tristate
rlabel metal2 s 473174 159200 473230 160000 6 la_output[120]
port 475 nsew signal tristate
rlabel metal2 s 477038 159200 477094 160000 6 la_output[121]
port 476 nsew signal tristate
rlabel metal2 s 480994 159200 481050 160000 6 la_output[122]
port 477 nsew signal tristate
rlabel metal2 s 484858 159200 484914 160000 6 la_output[123]
port 478 nsew signal tristate
rlabel metal2 s 488814 159200 488870 160000 6 la_output[124]
port 479 nsew signal tristate
rlabel metal2 s 492678 159200 492734 160000 6 la_output[125]
port 480 nsew signal tristate
rlabel metal2 s 496542 159200 496598 160000 6 la_output[126]
port 481 nsew signal tristate
rlabel metal2 s 500498 159200 500554 160000 6 la_output[127]
port 482 nsew signal tristate
rlabel metal2 s 52090 159200 52146 160000 6 la_output[12]
port 483 nsew signal tristate
rlabel metal2 s 55954 159200 56010 160000 6 la_output[13]
port 484 nsew signal tristate
rlabel metal2 s 59910 159200 59966 160000 6 la_output[14]
port 485 nsew signal tristate
rlabel metal2 s 63774 159200 63830 160000 6 la_output[15]
port 486 nsew signal tristate
rlabel metal2 s 67730 159200 67786 160000 6 la_output[16]
port 487 nsew signal tristate
rlabel metal2 s 71594 159200 71650 160000 6 la_output[17]
port 488 nsew signal tristate
rlabel metal2 s 75458 159200 75514 160000 6 la_output[18]
port 489 nsew signal tristate
rlabel metal2 s 79414 159200 79470 160000 6 la_output[19]
port 490 nsew signal tristate
rlabel metal2 s 9218 159200 9274 160000 6 la_output[1]
port 491 nsew signal tristate
rlabel metal2 s 83278 159200 83334 160000 6 la_output[20]
port 492 nsew signal tristate
rlabel metal2 s 87142 159200 87198 160000 6 la_output[21]
port 493 nsew signal tristate
rlabel metal2 s 91098 159200 91154 160000 6 la_output[22]
port 494 nsew signal tristate
rlabel metal2 s 94962 159200 95018 160000 6 la_output[23]
port 495 nsew signal tristate
rlabel metal2 s 98918 159200 98974 160000 6 la_output[24]
port 496 nsew signal tristate
rlabel metal2 s 102782 159200 102838 160000 6 la_output[25]
port 497 nsew signal tristate
rlabel metal2 s 106646 159200 106702 160000 6 la_output[26]
port 498 nsew signal tristate
rlabel metal2 s 110602 159200 110658 160000 6 la_output[27]
port 499 nsew signal tristate
rlabel metal2 s 114466 159200 114522 160000 6 la_output[28]
port 500 nsew signal tristate
rlabel metal2 s 118330 159200 118386 160000 6 la_output[29]
port 501 nsew signal tristate
rlabel metal2 s 13082 159200 13138 160000 6 la_output[2]
port 502 nsew signal tristate
rlabel metal2 s 122286 159200 122342 160000 6 la_output[30]
port 503 nsew signal tristate
rlabel metal2 s 126150 159200 126206 160000 6 la_output[31]
port 504 nsew signal tristate
rlabel metal2 s 130106 159200 130162 160000 6 la_output[32]
port 505 nsew signal tristate
rlabel metal2 s 133970 159200 134026 160000 6 la_output[33]
port 506 nsew signal tristate
rlabel metal2 s 137834 159200 137890 160000 6 la_output[34]
port 507 nsew signal tristate
rlabel metal2 s 141790 159200 141846 160000 6 la_output[35]
port 508 nsew signal tristate
rlabel metal2 s 145654 159200 145710 160000 6 la_output[36]
port 509 nsew signal tristate
rlabel metal2 s 149610 159200 149666 160000 6 la_output[37]
port 510 nsew signal tristate
rlabel metal2 s 153474 159200 153530 160000 6 la_output[38]
port 511 nsew signal tristate
rlabel metal2 s 157338 159200 157394 160000 6 la_output[39]
port 512 nsew signal tristate
rlabel metal2 s 17038 159200 17094 160000 6 la_output[3]
port 513 nsew signal tristate
rlabel metal2 s 161294 159200 161350 160000 6 la_output[40]
port 514 nsew signal tristate
rlabel metal2 s 165158 159200 165214 160000 6 la_output[41]
port 515 nsew signal tristate
rlabel metal2 s 169022 159200 169078 160000 6 la_output[42]
port 516 nsew signal tristate
rlabel metal2 s 172978 159200 173034 160000 6 la_output[43]
port 517 nsew signal tristate
rlabel metal2 s 176842 159200 176898 160000 6 la_output[44]
port 518 nsew signal tristate
rlabel metal2 s 180798 159200 180854 160000 6 la_output[45]
port 519 nsew signal tristate
rlabel metal2 s 184662 159200 184718 160000 6 la_output[46]
port 520 nsew signal tristate
rlabel metal2 s 188526 159200 188582 160000 6 la_output[47]
port 521 nsew signal tristate
rlabel metal2 s 192482 159200 192538 160000 6 la_output[48]
port 522 nsew signal tristate
rlabel metal2 s 196346 159200 196402 160000 6 la_output[49]
port 523 nsew signal tristate
rlabel metal2 s 20902 159200 20958 160000 6 la_output[4]
port 524 nsew signal tristate
rlabel metal2 s 200210 159200 200266 160000 6 la_output[50]
port 525 nsew signal tristate
rlabel metal2 s 204166 159200 204222 160000 6 la_output[51]
port 526 nsew signal tristate
rlabel metal2 s 208030 159200 208086 160000 6 la_output[52]
port 527 nsew signal tristate
rlabel metal2 s 211986 159200 212042 160000 6 la_output[53]
port 528 nsew signal tristate
rlabel metal2 s 215850 159200 215906 160000 6 la_output[54]
port 529 nsew signal tristate
rlabel metal2 s 219714 159200 219770 160000 6 la_output[55]
port 530 nsew signal tristate
rlabel metal2 s 223670 159200 223726 160000 6 la_output[56]
port 531 nsew signal tristate
rlabel metal2 s 227534 159200 227590 160000 6 la_output[57]
port 532 nsew signal tristate
rlabel metal2 s 231490 159200 231546 160000 6 la_output[58]
port 533 nsew signal tristate
rlabel metal2 s 235354 159200 235410 160000 6 la_output[59]
port 534 nsew signal tristate
rlabel metal2 s 24766 159200 24822 160000 6 la_output[5]
port 535 nsew signal tristate
rlabel metal2 s 239218 159200 239274 160000 6 la_output[60]
port 536 nsew signal tristate
rlabel metal2 s 243174 159200 243230 160000 6 la_output[61]
port 537 nsew signal tristate
rlabel metal2 s 247038 159200 247094 160000 6 la_output[62]
port 538 nsew signal tristate
rlabel metal2 s 250902 159200 250958 160000 6 la_output[63]
port 539 nsew signal tristate
rlabel metal2 s 254858 159200 254914 160000 6 la_output[64]
port 540 nsew signal tristate
rlabel metal2 s 258722 159200 258778 160000 6 la_output[65]
port 541 nsew signal tristate
rlabel metal2 s 262678 159200 262734 160000 6 la_output[66]
port 542 nsew signal tristate
rlabel metal2 s 266542 159200 266598 160000 6 la_output[67]
port 543 nsew signal tristate
rlabel metal2 s 270406 159200 270462 160000 6 la_output[68]
port 544 nsew signal tristate
rlabel metal2 s 274362 159200 274418 160000 6 la_output[69]
port 545 nsew signal tristate
rlabel metal2 s 28722 159200 28778 160000 6 la_output[6]
port 546 nsew signal tristate
rlabel metal2 s 278226 159200 278282 160000 6 la_output[70]
port 547 nsew signal tristate
rlabel metal2 s 282090 159200 282146 160000 6 la_output[71]
port 548 nsew signal tristate
rlabel metal2 s 286046 159200 286102 160000 6 la_output[72]
port 549 nsew signal tristate
rlabel metal2 s 289910 159200 289966 160000 6 la_output[73]
port 550 nsew signal tristate
rlabel metal2 s 293866 159200 293922 160000 6 la_output[74]
port 551 nsew signal tristate
rlabel metal2 s 297730 159200 297786 160000 6 la_output[75]
port 552 nsew signal tristate
rlabel metal2 s 301594 159200 301650 160000 6 la_output[76]
port 553 nsew signal tristate
rlabel metal2 s 305550 159200 305606 160000 6 la_output[77]
port 554 nsew signal tristate
rlabel metal2 s 309414 159200 309470 160000 6 la_output[78]
port 555 nsew signal tristate
rlabel metal2 s 313278 159200 313334 160000 6 la_output[79]
port 556 nsew signal tristate
rlabel metal2 s 32586 159200 32642 160000 6 la_output[7]
port 557 nsew signal tristate
rlabel metal2 s 317234 159200 317290 160000 6 la_output[80]
port 558 nsew signal tristate
rlabel metal2 s 321098 159200 321154 160000 6 la_output[81]
port 559 nsew signal tristate
rlabel metal2 s 325054 159200 325110 160000 6 la_output[82]
port 560 nsew signal tristate
rlabel metal2 s 328918 159200 328974 160000 6 la_output[83]
port 561 nsew signal tristate
rlabel metal2 s 332782 159200 332838 160000 6 la_output[84]
port 562 nsew signal tristate
rlabel metal2 s 336738 159200 336794 160000 6 la_output[85]
port 563 nsew signal tristate
rlabel metal2 s 340602 159200 340658 160000 6 la_output[86]
port 564 nsew signal tristate
rlabel metal2 s 344558 159200 344614 160000 6 la_output[87]
port 565 nsew signal tristate
rlabel metal2 s 348422 159200 348478 160000 6 la_output[88]
port 566 nsew signal tristate
rlabel metal2 s 352286 159200 352342 160000 6 la_output[89]
port 567 nsew signal tristate
rlabel metal2 s 36542 159200 36598 160000 6 la_output[8]
port 568 nsew signal tristate
rlabel metal2 s 356242 159200 356298 160000 6 la_output[90]
port 569 nsew signal tristate
rlabel metal2 s 360106 159200 360162 160000 6 la_output[91]
port 570 nsew signal tristate
rlabel metal2 s 363970 159200 364026 160000 6 la_output[92]
port 571 nsew signal tristate
rlabel metal2 s 367926 159200 367982 160000 6 la_output[93]
port 572 nsew signal tristate
rlabel metal2 s 371790 159200 371846 160000 6 la_output[94]
port 573 nsew signal tristate
rlabel metal2 s 375746 159200 375802 160000 6 la_output[95]
port 574 nsew signal tristate
rlabel metal2 s 379610 159200 379666 160000 6 la_output[96]
port 575 nsew signal tristate
rlabel metal2 s 383474 159200 383530 160000 6 la_output[97]
port 576 nsew signal tristate
rlabel metal2 s 387430 159200 387486 160000 6 la_output[98]
port 577 nsew signal tristate
rlabel metal2 s 391294 159200 391350 160000 6 la_output[99]
port 578 nsew signal tristate
rlabel metal2 s 40406 159200 40462 160000 6 la_output[9]
port 579 nsew signal tristate
rlabel metal3 s 0 157496 800 157616 6 mprj_ack_i
port 580 nsew signal input
rlabel metal2 s 504362 159200 504418 160000 6 mprj_adr_o[0]
port 581 nsew signal tristate
rlabel metal2 s 527730 159200 527786 160000 6 mprj_adr_o[10]
port 582 nsew signal tristate
rlabel metal2 s 529754 159200 529810 160000 6 mprj_adr_o[11]
port 583 nsew signal tristate
rlabel metal2 s 531686 159200 531742 160000 6 mprj_adr_o[12]
port 584 nsew signal tristate
rlabel metal2 s 533618 159200 533674 160000 6 mprj_adr_o[13]
port 585 nsew signal tristate
rlabel metal2 s 535550 159200 535606 160000 6 mprj_adr_o[14]
port 586 nsew signal tristate
rlabel metal2 s 537482 159200 537538 160000 6 mprj_adr_o[15]
port 587 nsew signal tristate
rlabel metal2 s 539506 159200 539562 160000 6 mprj_adr_o[16]
port 588 nsew signal tristate
rlabel metal2 s 541438 159200 541494 160000 6 mprj_adr_o[17]
port 589 nsew signal tristate
rlabel metal2 s 543370 159200 543426 160000 6 mprj_adr_o[18]
port 590 nsew signal tristate
rlabel metal2 s 545302 159200 545358 160000 6 mprj_adr_o[19]
port 591 nsew signal tristate
rlabel metal2 s 507306 159200 507362 160000 6 mprj_adr_o[1]
port 592 nsew signal tristate
rlabel metal2 s 547234 159200 547290 160000 6 mprj_adr_o[20]
port 593 nsew signal tristate
rlabel metal2 s 549166 159200 549222 160000 6 mprj_adr_o[21]
port 594 nsew signal tristate
rlabel metal2 s 551190 159200 551246 160000 6 mprj_adr_o[22]
port 595 nsew signal tristate
rlabel metal2 s 553122 159200 553178 160000 6 mprj_adr_o[23]
port 596 nsew signal tristate
rlabel metal2 s 555054 159200 555110 160000 6 mprj_adr_o[24]
port 597 nsew signal tristate
rlabel metal2 s 556986 159200 557042 160000 6 mprj_adr_o[25]
port 598 nsew signal tristate
rlabel metal2 s 558918 159200 558974 160000 6 mprj_adr_o[26]
port 599 nsew signal tristate
rlabel metal2 s 560942 159200 560998 160000 6 mprj_adr_o[27]
port 600 nsew signal tristate
rlabel metal2 s 562874 159200 562930 160000 6 mprj_adr_o[28]
port 601 nsew signal tristate
rlabel metal2 s 564806 159200 564862 160000 6 mprj_adr_o[29]
port 602 nsew signal tristate
rlabel metal2 s 510250 159200 510306 160000 6 mprj_adr_o[2]
port 603 nsew signal tristate
rlabel metal2 s 566738 159200 566794 160000 6 mprj_adr_o[30]
port 604 nsew signal tristate
rlabel metal2 s 568670 159200 568726 160000 6 mprj_adr_o[31]
port 605 nsew signal tristate
rlabel metal2 s 513102 159200 513158 160000 6 mprj_adr_o[3]
port 606 nsew signal tristate
rlabel metal2 s 516046 159200 516102 160000 6 mprj_adr_o[4]
port 607 nsew signal tristate
rlabel metal2 s 517978 159200 518034 160000 6 mprj_adr_o[5]
port 608 nsew signal tristate
rlabel metal2 s 520002 159200 520058 160000 6 mprj_adr_o[6]
port 609 nsew signal tristate
rlabel metal2 s 521934 159200 521990 160000 6 mprj_adr_o[7]
port 610 nsew signal tristate
rlabel metal2 s 523866 159200 523922 160000 6 mprj_adr_o[8]
port 611 nsew signal tristate
rlabel metal2 s 525798 159200 525854 160000 6 mprj_adr_o[9]
port 612 nsew signal tristate
rlabel metal2 s 501418 159200 501474 160000 6 mprj_cyc_o
port 613 nsew signal tristate
rlabel metal3 s 0 11296 800 11416 6 mprj_dat_i[0]
port 614 nsew signal input
rlabel metal3 s 0 56992 800 57112 6 mprj_dat_i[10]
port 615 nsew signal input
rlabel metal3 s 0 61480 800 61600 6 mprj_dat_i[11]
port 616 nsew signal input
rlabel metal3 s 0 66104 800 66224 6 mprj_dat_i[12]
port 617 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 mprj_dat_i[13]
port 618 nsew signal input
rlabel metal3 s 0 75216 800 75336 6 mprj_dat_i[14]
port 619 nsew signal input
rlabel metal3 s 0 79840 800 79960 6 mprj_dat_i[15]
port 620 nsew signal input
rlabel metal3 s 0 84328 800 84448 6 mprj_dat_i[16]
port 621 nsew signal input
rlabel metal3 s 0 88952 800 89072 6 mprj_dat_i[17]
port 622 nsew signal input
rlabel metal3 s 0 93576 800 93696 6 mprj_dat_i[18]
port 623 nsew signal input
rlabel metal3 s 0 98064 800 98184 6 mprj_dat_i[19]
port 624 nsew signal input
rlabel metal3 s 0 15784 800 15904 6 mprj_dat_i[1]
port 625 nsew signal input
rlabel metal3 s 0 102688 800 102808 6 mprj_dat_i[20]
port 626 nsew signal input
rlabel metal3 s 0 107176 800 107296 6 mprj_dat_i[21]
port 627 nsew signal input
rlabel metal3 s 0 111800 800 111920 6 mprj_dat_i[22]
port 628 nsew signal input
rlabel metal3 s 0 116424 800 116544 6 mprj_dat_i[23]
port 629 nsew signal input
rlabel metal3 s 0 120912 800 121032 6 mprj_dat_i[24]
port 630 nsew signal input
rlabel metal3 s 0 125536 800 125656 6 mprj_dat_i[25]
port 631 nsew signal input
rlabel metal3 s 0 130024 800 130144 6 mprj_dat_i[26]
port 632 nsew signal input
rlabel metal3 s 0 134648 800 134768 6 mprj_dat_i[27]
port 633 nsew signal input
rlabel metal3 s 0 139272 800 139392 6 mprj_dat_i[28]
port 634 nsew signal input
rlabel metal3 s 0 143760 800 143880 6 mprj_dat_i[29]
port 635 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 mprj_dat_i[2]
port 636 nsew signal input
rlabel metal3 s 0 148384 800 148504 6 mprj_dat_i[30]
port 637 nsew signal input
rlabel metal3 s 0 152872 800 152992 6 mprj_dat_i[31]
port 638 nsew signal input
rlabel metal3 s 0 25032 800 25152 6 mprj_dat_i[3]
port 639 nsew signal input
rlabel metal3 s 0 29520 800 29640 6 mprj_dat_i[4]
port 640 nsew signal input
rlabel metal3 s 0 34144 800 34264 6 mprj_dat_i[5]
port 641 nsew signal input
rlabel metal3 s 0 38632 800 38752 6 mprj_dat_i[6]
port 642 nsew signal input
rlabel metal3 s 0 43256 800 43376 6 mprj_dat_i[7]
port 643 nsew signal input
rlabel metal3 s 0 47880 800 48000 6 mprj_dat_i[8]
port 644 nsew signal input
rlabel metal3 s 0 52368 800 52488 6 mprj_dat_i[9]
port 645 nsew signal input
rlabel metal2 s 505374 159200 505430 160000 6 mprj_dat_o[0]
port 646 nsew signal tristate
rlabel metal2 s 528742 159200 528798 160000 6 mprj_dat_o[10]
port 647 nsew signal tristate
rlabel metal2 s 530674 159200 530730 160000 6 mprj_dat_o[11]
port 648 nsew signal tristate
rlabel metal2 s 532606 159200 532662 160000 6 mprj_dat_o[12]
port 649 nsew signal tristate
rlabel metal2 s 534630 159200 534686 160000 6 mprj_dat_o[13]
port 650 nsew signal tristate
rlabel metal2 s 536562 159200 536618 160000 6 mprj_dat_o[14]
port 651 nsew signal tristate
rlabel metal2 s 538494 159200 538550 160000 6 mprj_dat_o[15]
port 652 nsew signal tristate
rlabel metal2 s 540426 159200 540482 160000 6 mprj_dat_o[16]
port 653 nsew signal tristate
rlabel metal2 s 542358 159200 542414 160000 6 mprj_dat_o[17]
port 654 nsew signal tristate
rlabel metal2 s 544290 159200 544346 160000 6 mprj_dat_o[18]
port 655 nsew signal tristate
rlabel metal2 s 546314 159200 546370 160000 6 mprj_dat_o[19]
port 656 nsew signal tristate
rlabel metal2 s 508226 159200 508282 160000 6 mprj_dat_o[1]
port 657 nsew signal tristate
rlabel metal2 s 548246 159200 548302 160000 6 mprj_dat_o[20]
port 658 nsew signal tristate
rlabel metal2 s 550178 159200 550234 160000 6 mprj_dat_o[21]
port 659 nsew signal tristate
rlabel metal2 s 552110 159200 552166 160000 6 mprj_dat_o[22]
port 660 nsew signal tristate
rlabel metal2 s 554042 159200 554098 160000 6 mprj_dat_o[23]
port 661 nsew signal tristate
rlabel metal2 s 556066 159200 556122 160000 6 mprj_dat_o[24]
port 662 nsew signal tristate
rlabel metal2 s 557998 159200 558054 160000 6 mprj_dat_o[25]
port 663 nsew signal tristate
rlabel metal2 s 559930 159200 559986 160000 6 mprj_dat_o[26]
port 664 nsew signal tristate
rlabel metal2 s 561862 159200 561918 160000 6 mprj_dat_o[27]
port 665 nsew signal tristate
rlabel metal2 s 563794 159200 563850 160000 6 mprj_dat_o[28]
port 666 nsew signal tristate
rlabel metal2 s 565818 159200 565874 160000 6 mprj_dat_o[29]
port 667 nsew signal tristate
rlabel metal2 s 511170 159200 511226 160000 6 mprj_dat_o[2]
port 668 nsew signal tristate
rlabel metal2 s 567750 159200 567806 160000 6 mprj_dat_o[30]
port 669 nsew signal tristate
rlabel metal2 s 569682 159200 569738 160000 6 mprj_dat_o[31]
port 670 nsew signal tristate
rlabel metal2 s 514114 159200 514170 160000 6 mprj_dat_o[3]
port 671 nsew signal tristate
rlabel metal2 s 517058 159200 517114 160000 6 mprj_dat_o[4]
port 672 nsew signal tristate
rlabel metal2 s 518990 159200 519046 160000 6 mprj_dat_o[5]
port 673 nsew signal tristate
rlabel metal2 s 520922 159200 520978 160000 6 mprj_dat_o[6]
port 674 nsew signal tristate
rlabel metal2 s 522854 159200 522910 160000 6 mprj_dat_o[7]
port 675 nsew signal tristate
rlabel metal2 s 524878 159200 524934 160000 6 mprj_dat_o[8]
port 676 nsew signal tristate
rlabel metal2 s 526810 159200 526866 160000 6 mprj_dat_o[9]
port 677 nsew signal tristate
rlabel metal2 s 506294 159200 506350 160000 6 mprj_sel_o[0]
port 678 nsew signal tristate
rlabel metal2 s 509238 159200 509294 160000 6 mprj_sel_o[1]
port 679 nsew signal tristate
rlabel metal2 s 512182 159200 512238 160000 6 mprj_sel_o[2]
port 680 nsew signal tristate
rlabel metal2 s 515126 159200 515182 160000 6 mprj_sel_o[3]
port 681 nsew signal tristate
rlabel metal2 s 502430 159200 502486 160000 6 mprj_stb_o
port 682 nsew signal tristate
rlabel metal2 s 570694 159200 570750 160000 6 mprj_wb_iena
port 683 nsew signal tristate
rlabel metal2 s 503350 159200 503406 160000 6 mprj_we_o
port 684 nsew signal tristate
rlabel metal2 s 98366 0 98422 800 6 qspi_enabled
port 685 nsew signal tristate
rlabel metal2 s 577226 0 577282 800 6 ser_rx
port 686 nsew signal input
rlabel metal2 s 566554 0 566610 800 6 ser_tx
port 687 nsew signal tristate
rlabel metal2 s 529294 0 529350 800 6 spi_csb
port 688 nsew signal tristate
rlabel metal2 s 534630 0 534686 800 6 spi_enabled
port 689 nsew signal tristate
rlabel metal2 s 539966 0 540022 800 6 spi_sck
port 690 nsew signal tristate
rlabel metal2 s 545302 0 545358 800 6 spi_sdi
port 691 nsew signal input
rlabel metal2 s 550546 0 550602 800 6 spi_sdo
port 692 nsew signal tristate
rlabel metal2 s 555882 0 555938 800 6 spi_sdoenb
port 693 nsew signal tristate
rlabel metal2 s 295154 0 295210 800 6 sram_ro_addr[0]
port 694 nsew signal input
rlabel metal2 s 300490 0 300546 800 6 sram_ro_addr[1]
port 695 nsew signal input
rlabel metal2 s 305826 0 305882 800 6 sram_ro_addr[2]
port 696 nsew signal input
rlabel metal2 s 311162 0 311218 800 6 sram_ro_addr[3]
port 697 nsew signal input
rlabel metal2 s 316498 0 316554 800 6 sram_ro_addr[4]
port 698 nsew signal input
rlabel metal2 s 321834 0 321890 800 6 sram_ro_addr[5]
port 699 nsew signal input
rlabel metal2 s 327078 0 327134 800 6 sram_ro_addr[6]
port 700 nsew signal input
rlabel metal2 s 332414 0 332470 800 6 sram_ro_addr[7]
port 701 nsew signal input
rlabel metal2 s 284574 0 284630 800 6 sram_ro_clk
port 702 nsew signal input
rlabel metal2 s 289910 0 289966 800 6 sram_ro_csb
port 703 nsew signal input
rlabel metal2 s 337750 0 337806 800 6 sram_ro_data[0]
port 704 nsew signal tristate
rlabel metal2 s 390926 0 390982 800 6 sram_ro_data[10]
port 705 nsew signal tristate
rlabel metal2 s 396262 0 396318 800 6 sram_ro_data[11]
port 706 nsew signal tristate
rlabel metal2 s 401598 0 401654 800 6 sram_ro_data[12]
port 707 nsew signal tristate
rlabel metal2 s 406934 0 406990 800 6 sram_ro_data[13]
port 708 nsew signal tristate
rlabel metal2 s 412270 0 412326 800 6 sram_ro_data[14]
port 709 nsew signal tristate
rlabel metal2 s 417606 0 417662 800 6 sram_ro_data[15]
port 710 nsew signal tristate
rlabel metal2 s 422850 0 422906 800 6 sram_ro_data[16]
port 711 nsew signal tristate
rlabel metal2 s 428186 0 428242 800 6 sram_ro_data[17]
port 712 nsew signal tristate
rlabel metal2 s 433522 0 433578 800 6 sram_ro_data[18]
port 713 nsew signal tristate
rlabel metal2 s 438858 0 438914 800 6 sram_ro_data[19]
port 714 nsew signal tristate
rlabel metal2 s 343086 0 343142 800 6 sram_ro_data[1]
port 715 nsew signal tristate
rlabel metal2 s 444194 0 444250 800 6 sram_ro_data[20]
port 716 nsew signal tristate
rlabel metal2 s 449530 0 449586 800 6 sram_ro_data[21]
port 717 nsew signal tristate
rlabel metal2 s 454774 0 454830 800 6 sram_ro_data[22]
port 718 nsew signal tristate
rlabel metal2 s 460110 0 460166 800 6 sram_ro_data[23]
port 719 nsew signal tristate
rlabel metal2 s 465446 0 465502 800 6 sram_ro_data[24]
port 720 nsew signal tristate
rlabel metal2 s 470782 0 470838 800 6 sram_ro_data[25]
port 721 nsew signal tristate
rlabel metal2 s 476118 0 476174 800 6 sram_ro_data[26]
port 722 nsew signal tristate
rlabel metal2 s 481454 0 481510 800 6 sram_ro_data[27]
port 723 nsew signal tristate
rlabel metal2 s 486698 0 486754 800 6 sram_ro_data[28]
port 724 nsew signal tristate
rlabel metal2 s 492034 0 492090 800 6 sram_ro_data[29]
port 725 nsew signal tristate
rlabel metal2 s 348422 0 348478 800 6 sram_ro_data[2]
port 726 nsew signal tristate
rlabel metal2 s 497370 0 497426 800 6 sram_ro_data[30]
port 727 nsew signal tristate
rlabel metal2 s 502706 0 502762 800 6 sram_ro_data[31]
port 728 nsew signal tristate
rlabel metal2 s 353758 0 353814 800 6 sram_ro_data[3]
port 729 nsew signal tristate
rlabel metal2 s 359002 0 359058 800 6 sram_ro_data[4]
port 730 nsew signal tristate
rlabel metal2 s 364338 0 364394 800 6 sram_ro_data[5]
port 731 nsew signal tristate
rlabel metal2 s 369674 0 369730 800 6 sram_ro_data[6]
port 732 nsew signal tristate
rlabel metal2 s 375010 0 375066 800 6 sram_ro_data[7]
port 733 nsew signal tristate
rlabel metal2 s 380346 0 380402 800 6 sram_ro_data[8]
port 734 nsew signal tristate
rlabel metal2 s 385682 0 385738 800 6 sram_ro_data[9]
port 735 nsew signal tristate
rlabel metal2 s 561218 0 561274 800 6 trap
port 736 nsew signal tristate
rlabel metal2 s 571890 0 571946 800 6 uart_enabled
port 737 nsew signal tristate
rlabel metal2 s 571614 159200 571670 160000 6 user_irq_ena[0]
port 738 nsew signal tristate
rlabel metal2 s 572626 159200 572682 160000 6 user_irq_ena[1]
port 739 nsew signal tristate
rlabel metal2 s 573546 159200 573602 160000 6 user_irq_ena[2]
port 740 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 580000 160000
<< end >>
