magic
tech sky130A
magscale 1 2
timestamp 1667926533
<< nwell >>
rect 882 106885 159106 107451
rect 882 105797 159106 106363
rect 882 105265 74088 105275
rect 882 104719 159106 105265
rect 882 104709 48131 104719
rect 882 104177 25223 104187
rect 882 103631 159106 104177
rect 882 103621 18428 103631
rect 882 103089 7191 103099
rect 882 102543 159106 103089
rect 882 102533 26695 102543
rect 882 102001 15287 102011
rect 882 101455 159106 102001
rect 882 101445 7559 101455
rect 882 100913 22371 100923
rect 882 100367 159106 100913
rect 882 100357 51088 100367
rect 882 99825 6823 99835
rect 882 99279 159106 99825
rect 882 99269 18428 99279
rect 882 98737 38011 98747
rect 882 98191 159106 98737
rect 882 98181 27707 98191
rect 882 97649 17232 97659
rect 882 97103 159106 97649
rect 882 97093 60459 97103
rect 882 96561 7467 96571
rect 882 96015 159106 96561
rect 882 96005 6836 96015
rect 882 95473 20163 95483
rect 882 94927 159106 95473
rect 882 94917 39851 94927
rect 882 94385 15852 94395
rect 882 93839 159106 94385
rect 882 93829 28075 93839
rect 882 93297 6928 93307
rect 882 92751 159106 93297
rect 882 92741 7848 92751
rect 882 92209 48236 92219
rect 882 91663 159106 92209
rect 882 91653 11804 91663
rect 882 91121 15484 91131
rect 882 90575 159106 91121
rect 882 90565 10792 90575
rect 882 90033 10332 90043
rect 882 89487 159106 90033
rect 882 89477 24395 89487
rect 882 88945 87415 88955
rect 882 88399 159106 88945
rect 882 88389 7296 88399
rect 882 87857 54019 87867
rect 882 87311 159106 87857
rect 882 87301 28167 87311
rect 882 86769 11515 86779
rect 882 86223 159106 86769
rect 882 86213 24671 86223
rect 882 85681 49235 85691
rect 882 85125 159106 85681
rect 882 84593 19716 84603
rect 882 84047 159106 84593
rect 882 84037 39851 84047
rect 882 83505 8847 83515
rect 882 82959 159106 83505
rect 882 82949 17863 82959
rect 882 82417 8400 82427
rect 882 81871 159106 82417
rect 882 81861 68568 81871
rect 882 81329 27799 81339
rect 882 80783 159106 81329
rect 882 80773 122283 80783
rect 882 80241 12080 80251
rect 882 79695 159106 80241
rect 882 79685 8939 79695
rect 882 79153 16667 79163
rect 882 78607 159106 79153
rect 882 78597 8124 78607
rect 882 78065 18231 78075
rect 882 77519 159106 78065
rect 882 77509 16575 77519
rect 882 76977 12080 76987
rect 882 76431 159106 76977
rect 882 76421 29547 76431
rect 882 75889 20439 75899
rect 882 75343 159106 75889
rect 882 75333 53112 75343
rect 882 74801 64796 74811
rect 882 74255 159106 74801
rect 882 74245 97259 74255
rect 882 73713 58448 73723
rect 882 73167 159106 73713
rect 882 73157 120259 73167
rect 882 72625 49892 72635
rect 882 72079 159106 72625
rect 882 72069 59644 72079
rect 882 71537 72524 71547
rect 882 70991 159106 71537
rect 882 70981 25499 70991
rect 882 70449 19243 70459
rect 882 69903 159106 70449
rect 882 69893 21727 69903
rect 882 69361 136451 69371
rect 882 68815 159106 69361
rect 882 68805 5719 68815
rect 882 68273 13723 68283
rect 882 67727 159106 68273
rect 882 67717 37643 67727
rect 882 67185 15287 67195
rect 882 66639 159106 67185
rect 882 66629 23028 66639
rect 882 66097 4996 66107
rect 882 65551 159106 66097
rect 882 65541 55872 65551
rect 882 65009 40127 65019
rect 882 64463 159106 65009
rect 882 64453 14656 64463
rect 882 63921 5088 63931
rect 882 63375 159106 63921
rect 882 63365 48775 63375
rect 882 62833 7651 62843
rect 882 62287 159106 62833
rect 882 62277 18428 62287
rect 882 61745 41047 61755
rect 882 61199 159106 61745
rect 882 61189 4523 61199
rect 882 60657 12895 60667
rect 882 60111 159106 60657
rect 882 60101 23212 60111
rect 882 59569 10700 59579
rect 882 59023 159106 59569
rect 882 59013 4615 59023
rect 882 58481 49879 58491
rect 882 57935 159106 58481
rect 882 57925 64796 57935
rect 882 57393 17232 57403
rect 882 56847 159106 57393
rect 882 56837 5364 56847
rect 882 56305 10424 56315
rect 882 55759 159106 56305
rect 882 55749 14091 55759
rect 882 55217 52731 55227
rect 882 54671 159106 55217
rect 882 54661 5167 54671
rect 882 54129 22923 54139
rect 882 53583 159106 54129
rect 882 53573 35803 53583
rect 882 53041 8019 53051
rect 882 52495 159106 53041
rect 882 52485 5351 52495
rect 882 51953 4260 51963
rect 882 51407 159106 51953
rect 882 51397 9123 51407
rect 882 50865 25591 50875
rect 882 50309 159106 50865
rect 882 49777 37275 49787
rect 882 49231 159106 49777
rect 882 49221 34699 49231
rect 882 48689 4996 48699
rect 882 48143 159106 48689
rect 882 48133 51811 48143
rect 882 47601 42427 47611
rect 882 47055 159106 47601
rect 882 47045 138304 47055
rect 882 46513 8216 46523
rect 882 45967 159106 46513
rect 882 45957 14656 45967
rect 882 45425 115396 45435
rect 882 44879 159106 45425
rect 882 44869 4628 44879
rect 882 44337 44911 44347
rect 882 43791 159106 44337
rect 882 43781 10976 43791
rect 882 43249 121560 43259
rect 882 42703 159106 43249
rect 882 42693 50615 42703
rect 882 41615 159106 42171
rect 882 41605 16496 41615
rect 882 41073 9675 41083
rect 882 40527 159106 41073
rect 882 40517 43347 40527
rect 882 39985 4615 39995
rect 882 39439 159106 39985
rect 882 39429 4996 39439
rect 882 38897 23567 38907
rect 882 38351 159106 38897
rect 882 38341 14091 38351
rect 882 37809 7743 37819
rect 882 37263 159106 37809
rect 882 37253 15103 37263
rect 882 36721 5364 36731
rect 882 36175 159106 36721
rect 882 36165 27155 36175
rect 882 35633 82828 35643
rect 882 35087 159106 35633
rect 882 35077 78872 35087
rect 882 34545 59999 34555
rect 882 33999 159106 34545
rect 882 33989 57791 33999
rect 882 33457 51456 33467
rect 882 32911 159106 33457
rect 882 32901 106827 32911
rect 882 32369 8952 32379
rect 882 31823 159106 32369
rect 882 31813 19611 31823
rect 882 31281 4904 31291
rect 882 30735 159106 31281
rect 882 30725 8939 30735
rect 882 30193 8400 30203
rect 882 29647 159106 30193
rect 882 29637 11975 29647
rect 882 29105 38287 29115
rect 882 28559 159106 29105
rect 882 28549 37564 28559
rect 882 28017 18796 28027
rect 882 27471 159106 28017
rect 882 27461 8939 27471
rect 882 26929 5364 26939
rect 882 26383 159106 26929
rect 882 26373 33884 26383
rect 882 25841 105171 25851
rect 882 25295 159106 25841
rect 882 25285 20255 25295
rect 882 24753 4799 24763
rect 882 24207 159106 24753
rect 882 24197 28167 24207
rect 882 23665 39207 23675
rect 882 23119 159106 23665
rect 882 23109 35264 23119
rect 882 22577 21819 22587
rect 882 22031 159106 22577
rect 882 22021 4904 22031
rect 882 21489 9320 21499
rect 882 20943 159106 21489
rect 882 20933 8032 20943
rect 882 20401 12159 20411
rect 882 19855 159106 20401
rect 882 19845 11804 19855
rect 882 19313 4812 19323
rect 882 18767 159106 19313
rect 882 18757 47684 18767
rect 882 17679 159106 18235
rect 882 17669 7664 17679
rect 882 17137 8019 17147
rect 882 16591 159106 17137
rect 882 16581 31479 16591
rect 882 16049 20452 16059
rect 882 15503 159106 16049
rect 882 15493 4891 15503
rect 882 14961 12343 14971
rect 882 14415 159106 14961
rect 882 14405 7559 14415
rect 882 13873 53296 13883
rect 882 13327 159106 13873
rect 882 13317 12067 13327
rect 882 12785 5364 12795
rect 882 12239 159106 12785
rect 882 12229 17863 12239
rect 882 11697 36460 11707
rect 882 11151 159106 11697
rect 882 11141 4707 11151
rect 882 10609 8663 10619
rect 882 10063 159106 10609
rect 882 10053 11975 10063
rect 882 9521 17035 9531
rect 882 8975 159106 9521
rect 882 8965 7664 8975
rect 882 8433 27983 8443
rect 882 7887 159106 8433
rect 882 7877 22371 7887
rect 882 7345 90451 7355
rect 882 6799 159106 7345
rect 882 6789 95708 6799
rect 882 6257 151723 6267
rect 882 5711 159106 6257
rect 882 5701 72235 5711
rect 882 5169 115015 5179
rect 882 4613 159106 5169
rect 882 3525 159106 4091
rect 882 2437 159106 3003
<< obsli1 >>
rect 920 2159 159068 107729
<< obsm1 >>
rect 920 2128 159068 107840
<< metal2 >>
rect 2962 109200 3018 110000
rect 7930 109200 7986 110000
rect 12898 109200 12954 110000
rect 17866 109200 17922 110000
rect 22834 109200 22890 110000
rect 27802 109200 27858 110000
rect 32770 109200 32826 110000
rect 37738 109200 37794 110000
rect 42706 109200 42762 110000
rect 47674 109200 47730 110000
rect 52642 109200 52698 110000
rect 57610 109200 57666 110000
rect 62578 109200 62634 110000
rect 67546 109200 67602 110000
rect 72514 109200 72570 110000
rect 77482 109200 77538 110000
rect 82450 109200 82506 110000
rect 87418 109200 87474 110000
rect 92386 109200 92442 110000
rect 97354 109200 97410 110000
rect 102322 109200 102378 110000
rect 107290 109200 107346 110000
rect 112258 109200 112314 110000
rect 117226 109200 117282 110000
rect 122194 109200 122250 110000
rect 127162 109200 127218 110000
rect 132130 109200 132186 110000
rect 137098 109200 137154 110000
rect 142066 109200 142122 110000
rect 147034 109200 147090 110000
rect 152002 109200 152058 110000
rect 156970 109200 157026 110000
<< obsm2 >>
rect 1400 109144 2906 109290
rect 3074 109144 7874 109290
rect 8042 109144 12842 109290
rect 13010 109144 17810 109290
rect 17978 109144 22778 109290
rect 22946 109144 27746 109290
rect 27914 109144 32714 109290
rect 32882 109144 37682 109290
rect 37850 109144 42650 109290
rect 42818 109144 47618 109290
rect 47786 109144 52586 109290
rect 52754 109144 57554 109290
rect 57722 109144 62522 109290
rect 62690 109144 67490 109290
rect 67658 109144 72458 109290
rect 72626 109144 77426 109290
rect 77594 109144 82394 109290
rect 82562 109144 87362 109290
rect 87530 109144 92330 109290
rect 92498 109144 97298 109290
rect 97466 109144 102266 109290
rect 102434 109144 107234 109290
rect 107402 109144 112202 109290
rect 112370 109144 117170 109290
rect 117338 109144 122138 109290
rect 122306 109144 127106 109290
rect 127274 109144 132074 109290
rect 132242 109144 137042 109290
rect 137210 109144 142010 109290
rect 142178 109144 146978 109290
rect 147146 109144 151946 109290
rect 152114 109144 156914 109290
rect 157082 109144 158772 109290
rect 1400 2139 158772 109144
<< metal3 >>
rect 159200 106904 160000 107024
rect 159200 104592 160000 104712
rect 159200 102280 160000 102400
rect 159200 99968 160000 100088
rect 159200 97656 160000 97776
rect 159200 95344 160000 95464
rect 159200 93032 160000 93152
rect 159200 90720 160000 90840
rect 159200 88408 160000 88528
rect 159200 86096 160000 86216
rect 159200 83784 160000 83904
rect 159200 81472 160000 81592
rect 159200 79160 160000 79280
rect 159200 76848 160000 76968
rect 159200 74536 160000 74656
rect 159200 72224 160000 72344
rect 159200 69912 160000 70032
rect 159200 67600 160000 67720
rect 159200 65288 160000 65408
rect 159200 62976 160000 63096
rect 159200 60664 160000 60784
rect 159200 58352 160000 58472
rect 159200 56040 160000 56160
rect 159200 53728 160000 53848
rect 159200 51416 160000 51536
rect 159200 49104 160000 49224
rect 159200 46792 160000 46912
rect 159200 44480 160000 44600
rect 159200 42168 160000 42288
rect 159200 39856 160000 39976
rect 159200 37544 160000 37664
rect 159200 35232 160000 35352
rect 159200 32920 160000 33040
rect 159200 30608 160000 30728
rect 159200 28296 160000 28416
rect 159200 25984 160000 26104
rect 159200 23672 160000 23792
rect 159200 21360 160000 21480
rect 159200 19048 160000 19168
rect 159200 16736 160000 16856
rect 159200 14424 160000 14544
rect 159200 12112 160000 12232
rect 159200 9800 160000 9920
rect 159200 7488 160000 7608
rect 159200 5176 160000 5296
rect 159200 2864 160000 2984
<< obsm3 >>
rect 2865 107104 159282 107745
rect 2865 106824 159120 107104
rect 2865 104792 159282 106824
rect 2865 104512 159120 104792
rect 2865 102480 159282 104512
rect 2865 102200 159120 102480
rect 2865 100168 159282 102200
rect 2865 99888 159120 100168
rect 2865 97856 159282 99888
rect 2865 97576 159120 97856
rect 2865 95544 159282 97576
rect 2865 95264 159120 95544
rect 2865 93232 159282 95264
rect 2865 92952 159120 93232
rect 2865 90920 159282 92952
rect 2865 90640 159120 90920
rect 2865 88608 159282 90640
rect 2865 88328 159120 88608
rect 2865 86296 159282 88328
rect 2865 86016 159120 86296
rect 2865 83984 159282 86016
rect 2865 83704 159120 83984
rect 2865 81672 159282 83704
rect 2865 81392 159120 81672
rect 2865 79360 159282 81392
rect 2865 79080 159120 79360
rect 2865 77048 159282 79080
rect 2865 76768 159120 77048
rect 2865 74736 159282 76768
rect 2865 74456 159120 74736
rect 2865 72424 159282 74456
rect 2865 72144 159120 72424
rect 2865 70112 159282 72144
rect 2865 69832 159120 70112
rect 2865 67800 159282 69832
rect 2865 67520 159120 67800
rect 2865 65488 159282 67520
rect 2865 65208 159120 65488
rect 2865 63176 159282 65208
rect 2865 62896 159120 63176
rect 2865 60864 159282 62896
rect 2865 60584 159120 60864
rect 2865 58552 159282 60584
rect 2865 58272 159120 58552
rect 2865 56240 159282 58272
rect 2865 55960 159120 56240
rect 2865 53928 159282 55960
rect 2865 53648 159120 53928
rect 2865 51616 159282 53648
rect 2865 51336 159120 51616
rect 2865 49304 159282 51336
rect 2865 49024 159120 49304
rect 2865 46992 159282 49024
rect 2865 46712 159120 46992
rect 2865 44680 159282 46712
rect 2865 44400 159120 44680
rect 2865 42368 159282 44400
rect 2865 42088 159120 42368
rect 2865 40056 159282 42088
rect 2865 39776 159120 40056
rect 2865 37744 159282 39776
rect 2865 37464 159120 37744
rect 2865 35432 159282 37464
rect 2865 35152 159120 35432
rect 2865 33120 159282 35152
rect 2865 32840 159120 33120
rect 2865 30808 159282 32840
rect 2865 30528 159120 30808
rect 2865 28496 159282 30528
rect 2865 28216 159120 28496
rect 2865 26184 159282 28216
rect 2865 25904 159120 26184
rect 2865 23872 159282 25904
rect 2865 23592 159120 23872
rect 2865 21560 159282 23592
rect 2865 21280 159120 21560
rect 2865 19248 159282 21280
rect 2865 18968 159120 19248
rect 2865 16936 159282 18968
rect 2865 16656 159120 16936
rect 2865 14624 159282 16656
rect 2865 14344 159120 14624
rect 2865 12312 159282 14344
rect 2865 12032 159120 12312
rect 2865 10000 159282 12032
rect 2865 9720 159120 10000
rect 2865 7688 159282 9720
rect 2865 7408 159120 7688
rect 2865 5376 159282 7408
rect 2865 5096 159120 5376
rect 2865 3064 159282 5096
rect 2865 2784 159120 3064
rect 2865 2143 159282 2784
<< metal4 >>
rect 4024 2128 4344 107760
rect 19384 2128 19704 107760
rect 34744 2128 35064 107760
rect 50104 2128 50424 107760
rect 65464 2128 65784 107760
rect 80824 2128 81144 107760
rect 96184 2128 96504 107760
rect 111544 2128 111864 107760
rect 126904 2128 127224 107760
rect 142264 2128 142584 107760
rect 157624 2128 157944 107760
<< obsm4 >>
rect 4659 6427 19304 104957
rect 19784 6427 34664 104957
rect 35144 6427 50024 104957
rect 50504 6427 65384 104957
rect 65864 6427 80744 104957
rect 81224 6427 96104 104957
rect 96584 6427 111464 104957
rect 111944 6427 126824 104957
rect 127304 6427 141805 104957
<< labels >>
rlabel metal3 s 159200 2864 160000 2984 6 A0[0]
port 1 nsew signal input
rlabel metal3 s 159200 5176 160000 5296 6 A0[1]
port 2 nsew signal input
rlabel metal3 s 159200 7488 160000 7608 6 A0[2]
port 3 nsew signal input
rlabel metal3 s 159200 9800 160000 9920 6 A0[3]
port 4 nsew signal input
rlabel metal3 s 159200 12112 160000 12232 6 A0[4]
port 5 nsew signal input
rlabel metal3 s 159200 14424 160000 14544 6 A0[5]
port 6 nsew signal input
rlabel metal3 s 159200 16736 160000 16856 6 A0[6]
port 7 nsew signal input
rlabel metal3 s 159200 19048 160000 19168 6 A0[7]
port 8 nsew signal input
rlabel metal3 s 159200 69912 160000 70032 6 CLK
port 9 nsew signal input
rlabel metal3 s 159200 32920 160000 33040 6 Di0[0]
port 10 nsew signal input
rlabel metal3 s 159200 56040 160000 56160 6 Di0[10]
port 11 nsew signal input
rlabel metal3 s 159200 58352 160000 58472 6 Di0[11]
port 12 nsew signal input
rlabel metal3 s 159200 60664 160000 60784 6 Di0[12]
port 13 nsew signal input
rlabel metal3 s 159200 62976 160000 63096 6 Di0[13]
port 14 nsew signal input
rlabel metal3 s 159200 65288 160000 65408 6 Di0[14]
port 15 nsew signal input
rlabel metal3 s 159200 67600 160000 67720 6 Di0[15]
port 16 nsew signal input
rlabel metal3 s 159200 72224 160000 72344 6 Di0[16]
port 17 nsew signal input
rlabel metal3 s 159200 74536 160000 74656 6 Di0[17]
port 18 nsew signal input
rlabel metal3 s 159200 76848 160000 76968 6 Di0[18]
port 19 nsew signal input
rlabel metal3 s 159200 79160 160000 79280 6 Di0[19]
port 20 nsew signal input
rlabel metal3 s 159200 35232 160000 35352 6 Di0[1]
port 21 nsew signal input
rlabel metal3 s 159200 81472 160000 81592 6 Di0[20]
port 22 nsew signal input
rlabel metal3 s 159200 83784 160000 83904 6 Di0[21]
port 23 nsew signal input
rlabel metal3 s 159200 86096 160000 86216 6 Di0[22]
port 24 nsew signal input
rlabel metal3 s 159200 88408 160000 88528 6 Di0[23]
port 25 nsew signal input
rlabel metal3 s 159200 90720 160000 90840 6 Di0[24]
port 26 nsew signal input
rlabel metal3 s 159200 93032 160000 93152 6 Di0[25]
port 27 nsew signal input
rlabel metal3 s 159200 95344 160000 95464 6 Di0[26]
port 28 nsew signal input
rlabel metal3 s 159200 97656 160000 97776 6 Di0[27]
port 29 nsew signal input
rlabel metal3 s 159200 99968 160000 100088 6 Di0[28]
port 30 nsew signal input
rlabel metal3 s 159200 102280 160000 102400 6 Di0[29]
port 31 nsew signal input
rlabel metal3 s 159200 37544 160000 37664 6 Di0[2]
port 32 nsew signal input
rlabel metal3 s 159200 104592 160000 104712 6 Di0[30]
port 33 nsew signal input
rlabel metal3 s 159200 106904 160000 107024 6 Di0[31]
port 34 nsew signal input
rlabel metal3 s 159200 39856 160000 39976 6 Di0[3]
port 35 nsew signal input
rlabel metal3 s 159200 42168 160000 42288 6 Di0[4]
port 36 nsew signal input
rlabel metal3 s 159200 44480 160000 44600 6 Di0[5]
port 37 nsew signal input
rlabel metal3 s 159200 46792 160000 46912 6 Di0[6]
port 38 nsew signal input
rlabel metal3 s 159200 49104 160000 49224 6 Di0[7]
port 39 nsew signal input
rlabel metal3 s 159200 51416 160000 51536 6 Di0[8]
port 40 nsew signal input
rlabel metal3 s 159200 53728 160000 53848 6 Di0[9]
port 41 nsew signal input
rlabel metal2 s 2962 109200 3018 110000 6 Do0[0]
port 42 nsew signal output
rlabel metal2 s 52642 109200 52698 110000 6 Do0[10]
port 43 nsew signal output
rlabel metal2 s 57610 109200 57666 110000 6 Do0[11]
port 44 nsew signal output
rlabel metal2 s 62578 109200 62634 110000 6 Do0[12]
port 45 nsew signal output
rlabel metal2 s 67546 109200 67602 110000 6 Do0[13]
port 46 nsew signal output
rlabel metal2 s 72514 109200 72570 110000 6 Do0[14]
port 47 nsew signal output
rlabel metal2 s 77482 109200 77538 110000 6 Do0[15]
port 48 nsew signal output
rlabel metal2 s 82450 109200 82506 110000 6 Do0[16]
port 49 nsew signal output
rlabel metal2 s 87418 109200 87474 110000 6 Do0[17]
port 50 nsew signal output
rlabel metal2 s 92386 109200 92442 110000 6 Do0[18]
port 51 nsew signal output
rlabel metal2 s 97354 109200 97410 110000 6 Do0[19]
port 52 nsew signal output
rlabel metal2 s 7930 109200 7986 110000 6 Do0[1]
port 53 nsew signal output
rlabel metal2 s 102322 109200 102378 110000 6 Do0[20]
port 54 nsew signal output
rlabel metal2 s 107290 109200 107346 110000 6 Do0[21]
port 55 nsew signal output
rlabel metal2 s 112258 109200 112314 110000 6 Do0[22]
port 56 nsew signal output
rlabel metal2 s 117226 109200 117282 110000 6 Do0[23]
port 57 nsew signal output
rlabel metal2 s 122194 109200 122250 110000 6 Do0[24]
port 58 nsew signal output
rlabel metal2 s 127162 109200 127218 110000 6 Do0[25]
port 59 nsew signal output
rlabel metal2 s 132130 109200 132186 110000 6 Do0[26]
port 60 nsew signal output
rlabel metal2 s 137098 109200 137154 110000 6 Do0[27]
port 61 nsew signal output
rlabel metal2 s 142066 109200 142122 110000 6 Do0[28]
port 62 nsew signal output
rlabel metal2 s 147034 109200 147090 110000 6 Do0[29]
port 63 nsew signal output
rlabel metal2 s 12898 109200 12954 110000 6 Do0[2]
port 64 nsew signal output
rlabel metal2 s 152002 109200 152058 110000 6 Do0[30]
port 65 nsew signal output
rlabel metal2 s 156970 109200 157026 110000 6 Do0[31]
port 66 nsew signal output
rlabel metal2 s 17866 109200 17922 110000 6 Do0[3]
port 67 nsew signal output
rlabel metal2 s 22834 109200 22890 110000 6 Do0[4]
port 68 nsew signal output
rlabel metal2 s 27802 109200 27858 110000 6 Do0[5]
port 69 nsew signal output
rlabel metal2 s 32770 109200 32826 110000 6 Do0[6]
port 70 nsew signal output
rlabel metal2 s 37738 109200 37794 110000 6 Do0[7]
port 71 nsew signal output
rlabel metal2 s 42706 109200 42762 110000 6 Do0[8]
port 72 nsew signal output
rlabel metal2 s 47674 109200 47730 110000 6 Do0[9]
port 73 nsew signal output
rlabel metal3 s 159200 30608 160000 30728 6 EN0
port 74 nsew signal input
rlabel metal4 s 19384 2128 19704 107760 6 VGND
port 75 nsew ground bidirectional
rlabel metal4 s 50104 2128 50424 107760 6 VGND
port 75 nsew ground bidirectional
rlabel metal4 s 80824 2128 81144 107760 6 VGND
port 75 nsew ground bidirectional
rlabel metal4 s 111544 2128 111864 107760 6 VGND
port 75 nsew ground bidirectional
rlabel metal4 s 142264 2128 142584 107760 6 VGND
port 75 nsew ground bidirectional
rlabel metal4 s 4024 2128 4344 107760 6 VPWR
port 76 nsew power bidirectional
rlabel metal4 s 34744 2128 35064 107760 6 VPWR
port 76 nsew power bidirectional
rlabel metal4 s 65464 2128 65784 107760 6 VPWR
port 76 nsew power bidirectional
rlabel metal4 s 96184 2128 96504 107760 6 VPWR
port 76 nsew power bidirectional
rlabel metal4 s 126904 2128 127224 107760 6 VPWR
port 76 nsew power bidirectional
rlabel metal4 s 157624 2128 157944 107760 6 VPWR
port 76 nsew power bidirectional
rlabel metal3 s 159200 21360 160000 21480 6 WE0[0]
port 77 nsew signal input
rlabel metal3 s 159200 23672 160000 23792 6 WE0[1]
port 78 nsew signal input
rlabel metal3 s 159200 25984 160000 26104 6 WE0[2]
port 79 nsew signal input
rlabel metal3 s 159200 28296 160000 28416 6 WE0[3]
port 80 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 160000 110000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 61522492
string GDS_FILE /home/hosni/caravel_mgmt_soc_litex/openlane/RAM256/runs/RUN_2022.11.08_16.25.03/results/signoff/RAM256.magic.gds
string GDS_START 184572
<< end >>

