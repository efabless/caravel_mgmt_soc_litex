magic
tech sky130A
magscale 1 2
timestamp 1665156864
<< obsli1 >>
rect 920 2159 98992 137649
<< obsm1 >>
rect 920 1368 99438 138168
<< metal2 >>
rect 2870 139200 2926 140000
rect 5906 139200 5962 140000
rect 8942 139200 8998 140000
rect 11978 139200 12034 140000
rect 15014 139200 15070 140000
rect 18050 139200 18106 140000
rect 21086 139200 21142 140000
rect 24122 139200 24178 140000
rect 27158 139200 27214 140000
rect 30194 139200 30250 140000
rect 33230 139200 33286 140000
rect 36266 139200 36322 140000
rect 39302 139200 39358 140000
rect 42338 139200 42394 140000
rect 45374 139200 45430 140000
rect 48410 139200 48466 140000
rect 51446 139200 51502 140000
rect 54482 139200 54538 140000
rect 57518 139200 57574 140000
rect 60554 139200 60610 140000
rect 63590 139200 63646 140000
rect 66626 139200 66682 140000
rect 69662 139200 69718 140000
rect 72698 139200 72754 140000
rect 75734 139200 75790 140000
rect 78770 139200 78826 140000
rect 81806 139200 81862 140000
rect 84842 139200 84898 140000
rect 87878 139200 87934 140000
rect 90914 139200 90970 140000
rect 93950 139200 94006 140000
rect 96986 139200 97042 140000
<< obsm2 >>
rect 1214 139144 2814 139346
rect 2982 139144 5850 139346
rect 6018 139144 8886 139346
rect 9054 139144 11922 139346
rect 12090 139144 14958 139346
rect 15126 139144 17994 139346
rect 18162 139144 21030 139346
rect 21198 139144 24066 139346
rect 24234 139144 27102 139346
rect 27270 139144 30138 139346
rect 30306 139144 33174 139346
rect 33342 139144 36210 139346
rect 36378 139144 39246 139346
rect 39414 139144 42282 139346
rect 42450 139144 45318 139346
rect 45486 139144 48354 139346
rect 48522 139144 51390 139346
rect 51558 139144 54426 139346
rect 54594 139144 57462 139346
rect 57630 139144 60498 139346
rect 60666 139144 63534 139346
rect 63702 139144 66570 139346
rect 66738 139144 69606 139346
rect 69774 139144 72642 139346
rect 72810 139144 75678 139346
rect 75846 139144 78714 139346
rect 78882 139144 81750 139346
rect 81918 139144 84786 139346
rect 84954 139144 87822 139346
rect 87990 139144 90858 139346
rect 91026 139144 93894 139346
rect 94062 139144 96930 139346
rect 97098 139144 99432 139346
rect 1214 1362 99432 139144
<< metal3 >>
rect 99200 137232 100000 137352
rect 99200 134240 100000 134360
rect 99200 131248 100000 131368
rect 99200 128256 100000 128376
rect 99200 125264 100000 125384
rect 99200 122272 100000 122392
rect 99200 119280 100000 119400
rect 99200 116288 100000 116408
rect 99200 113296 100000 113416
rect 99200 110304 100000 110424
rect 99200 107312 100000 107432
rect 99200 104320 100000 104440
rect 99200 101328 100000 101448
rect 99200 98336 100000 98456
rect 99200 95344 100000 95464
rect 99200 92352 100000 92472
rect 99200 89360 100000 89480
rect 99200 86368 100000 86488
rect 99200 83376 100000 83496
rect 99200 80384 100000 80504
rect 99200 77392 100000 77512
rect 99200 74400 100000 74520
rect 99200 71408 100000 71528
rect 99200 68416 100000 68536
rect 99200 65424 100000 65544
rect 99200 62432 100000 62552
rect 99200 59440 100000 59560
rect 99200 56448 100000 56568
rect 99200 53456 100000 53576
rect 99200 50464 100000 50584
rect 99200 47472 100000 47592
rect 99200 44480 100000 44600
rect 99200 41488 100000 41608
rect 99200 38496 100000 38616
rect 99200 35504 100000 35624
rect 99200 32512 100000 32632
rect 99200 29520 100000 29640
rect 99200 26528 100000 26648
rect 99200 23536 100000 23656
rect 99200 20544 100000 20664
rect 99200 17552 100000 17672
rect 99200 14560 100000 14680
rect 99200 11568 100000 11688
rect 99200 8576 100000 8696
rect 99200 5584 100000 5704
rect 99200 2592 100000 2712
<< obsm3 >>
rect 1209 137432 99200 137733
rect 1209 137152 99120 137432
rect 1209 134440 99200 137152
rect 1209 134160 99120 134440
rect 1209 131448 99200 134160
rect 1209 131168 99120 131448
rect 1209 128456 99200 131168
rect 1209 128176 99120 128456
rect 1209 125464 99200 128176
rect 1209 125184 99120 125464
rect 1209 122472 99200 125184
rect 1209 122192 99120 122472
rect 1209 119480 99200 122192
rect 1209 119200 99120 119480
rect 1209 116488 99200 119200
rect 1209 116208 99120 116488
rect 1209 113496 99200 116208
rect 1209 113216 99120 113496
rect 1209 110504 99200 113216
rect 1209 110224 99120 110504
rect 1209 107512 99200 110224
rect 1209 107232 99120 107512
rect 1209 104520 99200 107232
rect 1209 104240 99120 104520
rect 1209 101528 99200 104240
rect 1209 101248 99120 101528
rect 1209 98536 99200 101248
rect 1209 98256 99120 98536
rect 1209 95544 99200 98256
rect 1209 95264 99120 95544
rect 1209 92552 99200 95264
rect 1209 92272 99120 92552
rect 1209 89560 99200 92272
rect 1209 89280 99120 89560
rect 1209 86568 99200 89280
rect 1209 86288 99120 86568
rect 1209 83576 99200 86288
rect 1209 83296 99120 83576
rect 1209 80584 99200 83296
rect 1209 80304 99120 80584
rect 1209 77592 99200 80304
rect 1209 77312 99120 77592
rect 1209 74600 99200 77312
rect 1209 74320 99120 74600
rect 1209 71608 99200 74320
rect 1209 71328 99120 71608
rect 1209 68616 99200 71328
rect 1209 68336 99120 68616
rect 1209 65624 99200 68336
rect 1209 65344 99120 65624
rect 1209 62632 99200 65344
rect 1209 62352 99120 62632
rect 1209 59640 99200 62352
rect 1209 59360 99120 59640
rect 1209 56648 99200 59360
rect 1209 56368 99120 56648
rect 1209 53656 99200 56368
rect 1209 53376 99120 53656
rect 1209 50664 99200 53376
rect 1209 50384 99120 50664
rect 1209 47672 99200 50384
rect 1209 47392 99120 47672
rect 1209 44680 99200 47392
rect 1209 44400 99120 44680
rect 1209 41688 99200 44400
rect 1209 41408 99120 41688
rect 1209 38696 99200 41408
rect 1209 38416 99120 38696
rect 1209 35704 99200 38416
rect 1209 35424 99120 35704
rect 1209 32712 99200 35424
rect 1209 32432 99120 32712
rect 1209 29720 99200 32432
rect 1209 29440 99120 29720
rect 1209 26728 99200 29440
rect 1209 26448 99120 26728
rect 1209 23736 99200 26448
rect 1209 23456 99120 23736
rect 1209 20744 99200 23456
rect 1209 20464 99120 20744
rect 1209 17752 99200 20464
rect 1209 17472 99120 17752
rect 1209 14760 99200 17472
rect 1209 14480 99120 14760
rect 1209 11768 99200 14480
rect 1209 11488 99120 11768
rect 1209 8776 99200 11488
rect 1209 8496 99120 8776
rect 1209 5784 99200 8496
rect 1209 5504 99120 5784
rect 1209 2792 99200 5504
rect 1209 2512 99120 2792
rect 1209 2143 99200 2512
<< metal4 >>
rect -1260 -4 -940 139812
rect -600 656 -280 139152
rect 4024 -4 4344 139812
rect 19384 -4 19704 139812
rect 34744 -4 35064 139812
rect 50104 -4 50424 139812
rect 65464 -4 65784 139812
rect 80824 -4 81144 139812
rect 96184 -4 96504 139812
rect 100192 656 100512 139152
rect 100852 -4 101172 139812
<< obsm4 >>
rect 4475 3979 19304 137189
rect 19784 3979 34664 137189
rect 35144 3979 50024 137189
rect 50504 3979 65384 137189
rect 65864 3979 80744 137189
rect 81224 3979 96104 137189
rect 96584 3979 97829 137189
<< metal5 >>
rect -1260 139492 101172 139812
rect -600 138832 100512 139152
rect -1260 135346 101172 135666
rect -1260 122346 101172 122666
rect -1260 109346 101172 109666
rect -1260 96346 101172 96666
rect -1260 83346 101172 83666
rect -1260 70346 101172 70666
rect -1260 57346 101172 57666
rect -1260 44346 101172 44666
rect -1260 31346 101172 31666
rect -1260 18346 101172 18666
rect -1260 5346 101172 5666
rect -600 656 100512 976
rect -1260 -4 101172 316
<< labels >>
rlabel metal3 s 99200 2592 100000 2712 6 A[0]
port 1 nsew signal input
rlabel metal3 s 99200 5584 100000 5704 6 A[1]
port 2 nsew signal input
rlabel metal3 s 99200 8576 100000 8696 6 A[2]
port 3 nsew signal input
rlabel metal3 s 99200 11568 100000 11688 6 A[3]
port 4 nsew signal input
rlabel metal3 s 99200 14560 100000 14680 6 A[4]
port 5 nsew signal input
rlabel metal3 s 99200 17552 100000 17672 6 A[5]
port 6 nsew signal input
rlabel metal3 s 99200 20544 100000 20664 6 A[6]
port 7 nsew signal input
rlabel metal3 s 99200 23536 100000 23656 6 A[7]
port 8 nsew signal input
rlabel metal3 s 99200 89360 100000 89480 6 CLK
port 9 nsew signal input
rlabel metal3 s 99200 41488 100000 41608 6 Di[0]
port 10 nsew signal input
rlabel metal3 s 99200 71408 100000 71528 6 Di[10]
port 11 nsew signal input
rlabel metal3 s 99200 74400 100000 74520 6 Di[11]
port 12 nsew signal input
rlabel metal3 s 99200 77392 100000 77512 6 Di[12]
port 13 nsew signal input
rlabel metal3 s 99200 80384 100000 80504 6 Di[13]
port 14 nsew signal input
rlabel metal3 s 99200 83376 100000 83496 6 Di[14]
port 15 nsew signal input
rlabel metal3 s 99200 86368 100000 86488 6 Di[15]
port 16 nsew signal input
rlabel metal3 s 99200 92352 100000 92472 6 Di[16]
port 17 nsew signal input
rlabel metal3 s 99200 95344 100000 95464 6 Di[17]
port 18 nsew signal input
rlabel metal3 s 99200 98336 100000 98456 6 Di[18]
port 19 nsew signal input
rlabel metal3 s 99200 101328 100000 101448 6 Di[19]
port 20 nsew signal input
rlabel metal3 s 99200 44480 100000 44600 6 Di[1]
port 21 nsew signal input
rlabel metal3 s 99200 104320 100000 104440 6 Di[20]
port 22 nsew signal input
rlabel metal3 s 99200 107312 100000 107432 6 Di[21]
port 23 nsew signal input
rlabel metal3 s 99200 110304 100000 110424 6 Di[22]
port 24 nsew signal input
rlabel metal3 s 99200 113296 100000 113416 6 Di[23]
port 25 nsew signal input
rlabel metal3 s 99200 116288 100000 116408 6 Di[24]
port 26 nsew signal input
rlabel metal3 s 99200 119280 100000 119400 6 Di[25]
port 27 nsew signal input
rlabel metal3 s 99200 122272 100000 122392 6 Di[26]
port 28 nsew signal input
rlabel metal3 s 99200 125264 100000 125384 6 Di[27]
port 29 nsew signal input
rlabel metal3 s 99200 128256 100000 128376 6 Di[28]
port 30 nsew signal input
rlabel metal3 s 99200 131248 100000 131368 6 Di[29]
port 31 nsew signal input
rlabel metal3 s 99200 47472 100000 47592 6 Di[2]
port 32 nsew signal input
rlabel metal3 s 99200 134240 100000 134360 6 Di[30]
port 33 nsew signal input
rlabel metal3 s 99200 137232 100000 137352 6 Di[31]
port 34 nsew signal input
rlabel metal3 s 99200 50464 100000 50584 6 Di[3]
port 35 nsew signal input
rlabel metal3 s 99200 53456 100000 53576 6 Di[4]
port 36 nsew signal input
rlabel metal3 s 99200 56448 100000 56568 6 Di[5]
port 37 nsew signal input
rlabel metal3 s 99200 59440 100000 59560 6 Di[6]
port 38 nsew signal input
rlabel metal3 s 99200 62432 100000 62552 6 Di[7]
port 39 nsew signal input
rlabel metal3 s 99200 65424 100000 65544 6 Di[8]
port 40 nsew signal input
rlabel metal3 s 99200 68416 100000 68536 6 Di[9]
port 41 nsew signal input
rlabel metal2 s 2870 139200 2926 140000 6 Do[0]
port 42 nsew signal output
rlabel metal2 s 33230 139200 33286 140000 6 Do[10]
port 43 nsew signal output
rlabel metal2 s 36266 139200 36322 140000 6 Do[11]
port 44 nsew signal output
rlabel metal2 s 39302 139200 39358 140000 6 Do[12]
port 45 nsew signal output
rlabel metal2 s 42338 139200 42394 140000 6 Do[13]
port 46 nsew signal output
rlabel metal2 s 45374 139200 45430 140000 6 Do[14]
port 47 nsew signal output
rlabel metal2 s 48410 139200 48466 140000 6 Do[15]
port 48 nsew signal output
rlabel metal2 s 51446 139200 51502 140000 6 Do[16]
port 49 nsew signal output
rlabel metal2 s 54482 139200 54538 140000 6 Do[17]
port 50 nsew signal output
rlabel metal2 s 57518 139200 57574 140000 6 Do[18]
port 51 nsew signal output
rlabel metal2 s 60554 139200 60610 140000 6 Do[19]
port 52 nsew signal output
rlabel metal2 s 5906 139200 5962 140000 6 Do[1]
port 53 nsew signal output
rlabel metal2 s 63590 139200 63646 140000 6 Do[20]
port 54 nsew signal output
rlabel metal2 s 66626 139200 66682 140000 6 Do[21]
port 55 nsew signal output
rlabel metal2 s 69662 139200 69718 140000 6 Do[22]
port 56 nsew signal output
rlabel metal2 s 72698 139200 72754 140000 6 Do[23]
port 57 nsew signal output
rlabel metal2 s 75734 139200 75790 140000 6 Do[24]
port 58 nsew signal output
rlabel metal2 s 78770 139200 78826 140000 6 Do[25]
port 59 nsew signal output
rlabel metal2 s 81806 139200 81862 140000 6 Do[26]
port 60 nsew signal output
rlabel metal2 s 84842 139200 84898 140000 6 Do[27]
port 61 nsew signal output
rlabel metal2 s 87878 139200 87934 140000 6 Do[28]
port 62 nsew signal output
rlabel metal2 s 90914 139200 90970 140000 6 Do[29]
port 63 nsew signal output
rlabel metal2 s 8942 139200 8998 140000 6 Do[2]
port 64 nsew signal output
rlabel metal2 s 93950 139200 94006 140000 6 Do[30]
port 65 nsew signal output
rlabel metal2 s 96986 139200 97042 140000 6 Do[31]
port 66 nsew signal output
rlabel metal2 s 11978 139200 12034 140000 6 Do[3]
port 67 nsew signal output
rlabel metal2 s 15014 139200 15070 140000 6 Do[4]
port 68 nsew signal output
rlabel metal2 s 18050 139200 18106 140000 6 Do[5]
port 69 nsew signal output
rlabel metal2 s 21086 139200 21142 140000 6 Do[6]
port 70 nsew signal output
rlabel metal2 s 24122 139200 24178 140000 6 Do[7]
port 71 nsew signal output
rlabel metal2 s 27158 139200 27214 140000 6 Do[8]
port 72 nsew signal output
rlabel metal2 s 30194 139200 30250 140000 6 Do[9]
port 73 nsew signal output
rlabel metal3 s 99200 38496 100000 38616 6 EN
port 74 nsew signal input
rlabel metal4 s -1260 -4 -940 139812 4 VGND
port 75 nsew ground bidirectional
rlabel metal5 s -1260 -4 101172 316 6 VGND
port 75 nsew ground bidirectional
rlabel metal5 s -1260 139492 101172 139812 6 VGND
port 75 nsew ground bidirectional
rlabel metal4 s 100852 -4 101172 139812 6 VGND
port 75 nsew ground bidirectional
rlabel metal4 s 19384 -4 19704 139812 6 VGND
port 75 nsew ground bidirectional
rlabel metal4 s 50104 -4 50424 139812 6 VGND
port 75 nsew ground bidirectional
rlabel metal4 s 80824 -4 81144 139812 6 VGND
port 75 nsew ground bidirectional
rlabel metal5 s -1260 18346 101172 18666 6 VGND
port 75 nsew ground bidirectional
rlabel metal5 s -1260 44346 101172 44666 6 VGND
port 75 nsew ground bidirectional
rlabel metal5 s -1260 70346 101172 70666 6 VGND
port 75 nsew ground bidirectional
rlabel metal5 s -1260 96346 101172 96666 6 VGND
port 75 nsew ground bidirectional
rlabel metal5 s -1260 122346 101172 122666 6 VGND
port 75 nsew ground bidirectional
rlabel metal4 s -600 656 -280 139152 4 VPWR
port 76 nsew power bidirectional
rlabel metal5 s -600 656 100512 976 6 VPWR
port 76 nsew power bidirectional
rlabel metal5 s -600 138832 100512 139152 6 VPWR
port 76 nsew power bidirectional
rlabel metal4 s 100192 656 100512 139152 6 VPWR
port 76 nsew power bidirectional
rlabel metal4 s 4024 -4 4344 139812 6 VPWR
port 76 nsew power bidirectional
rlabel metal4 s 34744 -4 35064 139812 6 VPWR
port 76 nsew power bidirectional
rlabel metal4 s 65464 -4 65784 139812 6 VPWR
port 76 nsew power bidirectional
rlabel metal4 s 96184 -4 96504 139812 6 VPWR
port 76 nsew power bidirectional
rlabel metal5 s -1260 5346 101172 5666 6 VPWR
port 76 nsew power bidirectional
rlabel metal5 s -1260 31346 101172 31666 6 VPWR
port 76 nsew power bidirectional
rlabel metal5 s -1260 57346 101172 57666 6 VPWR
port 76 nsew power bidirectional
rlabel metal5 s -1260 83346 101172 83666 6 VPWR
port 76 nsew power bidirectional
rlabel metal5 s -1260 109346 101172 109666 6 VPWR
port 76 nsew power bidirectional
rlabel metal5 s -1260 135346 101172 135666 6 VPWR
port 76 nsew power bidirectional
rlabel metal3 s 99200 26528 100000 26648 6 WE[0]
port 77 nsew signal input
rlabel metal3 s 99200 29520 100000 29640 6 WE[1]
port 78 nsew signal input
rlabel metal3 s 99200 32512 100000 32632 6 WE[2]
port 79 nsew signal input
rlabel metal3 s 99200 35504 100000 35624 6 WE[3]
port 80 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 100000 140000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 56317716
string GDS_FILE /home/kareem_farid/caravel_mgmt_soc_litex/openlane/DFFRAM/runs/22_10_07_08_04/results/signoff/DFFRAM.magic.gds
string GDS_START 184572
<< end >>

