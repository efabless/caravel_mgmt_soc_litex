VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mgmt_core_wrapper
  CLASS BLOCK ;
  FOREIGN mgmt_core_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2520.000 BY 740.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -5.380 -0.020 -3.780 739.860 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 -0.020 2525.260 1.580 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 738.260 2525.260 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2523.660 -0.020 2525.260 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 32.640 -0.020 34.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 82.640 -0.020 84.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 132.640 -0.020 134.240 52.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 132.640 585.510 134.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 182.640 -0.020 184.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 232.640 -0.020 234.240 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 232.640 554.875 234.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 282.640 -0.020 284.240 52.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 282.640 585.510 284.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 332.640 -0.020 334.240 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 332.640 554.875 334.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 382.640 -0.020 384.240 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 382.640 554.875 384.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 432.640 -0.020 434.240 52.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 432.640 585.510 434.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 482.640 -0.020 484.240 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 482.640 554.875 484.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 532.640 -0.020 534.240 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 532.640 554.875 534.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 582.640 -0.020 584.240 52.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 582.640 585.510 584.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.640 -0.020 634.240 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.640 554.875 634.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 682.640 -0.020 684.240 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 682.640 554.875 684.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 732.640 -0.020 734.240 52.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 732.640 585.510 734.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 782.640 -0.020 784.240 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 782.640 554.875 784.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 832.640 -0.020 834.240 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 832.640 554.875 834.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 882.640 -0.020 884.240 52.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 882.640 585.510 884.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 932.640 -0.020 934.240 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 932.640 554.875 934.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 982.640 -0.020 984.240 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 982.640 554.875 984.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1032.640 -0.020 1034.240 52.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 1032.640 585.510 1034.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1082.640 -0.020 1084.240 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 1082.640 554.875 1084.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1132.640 -0.020 1134.240 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 1132.640 554.875 1134.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1182.640 -0.020 1184.240 52.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 1182.640 585.510 1184.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1232.640 -0.020 1234.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1282.640 -0.020 1284.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1332.640 -0.020 1334.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1382.640 -0.020 1384.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1432.640 -0.020 1434.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1482.640 -0.020 1484.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1532.640 -0.020 1534.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1582.640 -0.020 1584.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1632.640 -0.020 1634.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1682.640 -0.020 1684.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1732.640 -0.020 1734.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1782.640 -0.020 1784.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1832.640 -0.020 1834.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1882.640 -0.020 1884.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1932.640 -0.020 1934.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1982.640 -0.020 1984.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2032.640 -0.020 2034.240 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2032.640 581.160 2034.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2082.640 -0.020 2084.240 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2082.640 581.160 2084.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2132.640 -0.020 2134.240 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2132.640 581.160 2134.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2182.640 -0.020 2184.240 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2182.640 581.160 2184.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2232.640 -0.020 2234.240 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2232.640 581.160 2234.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2282.640 -0.020 2284.240 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2282.640 581.160 2284.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2332.640 -0.020 2334.240 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2332.640 581.160 2334.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2382.640 -0.020 2384.240 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2382.640 581.160 2384.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2432.640 -0.020 2434.240 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2432.640 581.160 2434.240 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2482.640 -0.020 2484.240 739.860 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 38.330 2525.260 39.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 88.330 2525.260 89.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 138.330 2525.260 139.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 188.330 2525.260 189.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 238.330 2525.260 239.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 288.330 2525.260 289.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 338.330 2525.260 339.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 388.330 2525.260 389.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 438.330 2525.260 439.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 488.330 2525.260 489.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 538.330 2525.260 539.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 588.330 2525.260 589.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 638.330 2525.260 639.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 688.330 2525.260 689.930 ;
    END
    PORT
      LAYER met4 ;
        RECT 2505.740 35.120 2507.340 625.840 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -2.080 3.280 -0.480 736.560 ;
    END
    PORT
      LAYER met5 ;
        RECT -2.080 3.280 2521.960 4.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -2.080 734.960 2521.960 736.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 2520.360 3.280 2521.960 736.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.040 -0.020 22.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.040 -0.020 72.640 52.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.040 585.510 72.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 121.040 -0.020 122.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.040 -0.020 172.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 221.040 -0.020 222.640 52.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 221.040 585.510 222.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 271.040 -0.020 272.640 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 271.040 554.875 272.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 -0.020 322.640 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 554.875 322.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 371.040 -0.020 372.640 52.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 371.040 585.510 372.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 421.040 -0.020 422.640 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 421.040 554.875 422.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 471.040 -0.020 472.640 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 471.040 554.875 472.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 521.040 -0.020 522.640 52.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 521.040 585.510 522.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 571.040 -0.020 572.640 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 571.040 554.875 572.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 621.040 -0.020 622.640 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 621.040 554.875 622.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.040 -0.020 672.640 52.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.040 585.510 672.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 721.040 -0.020 722.640 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 721.040 554.875 722.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 771.040 -0.020 772.640 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 771.040 554.875 772.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 821.040 -0.020 822.640 52.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 821.040 585.510 822.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 871.040 -0.020 872.640 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 871.040 554.875 872.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.040 -0.020 922.640 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.040 554.875 922.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 971.040 -0.020 972.640 52.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 971.040 585.510 972.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.040 -0.020 1022.640 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.040 554.875 1022.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1071.040 -0.020 1072.640 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 1071.040 554.875 1072.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1121.040 -0.020 1122.640 52.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 1121.040 585.510 1122.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1171.040 -0.020 1172.640 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 1171.040 554.875 1172.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1221.040 -0.020 1222.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1271.040 -0.020 1272.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1321.040 -0.020 1322.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1371.040 -0.020 1372.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1421.040 -0.020 1422.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1471.040 -0.020 1472.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1521.040 -0.020 1522.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1571.040 -0.020 1572.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1621.040 -0.020 1622.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1671.040 -0.020 1672.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1721.040 -0.020 1722.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1771.040 -0.020 1772.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1821.040 -0.020 1822.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1871.040 -0.020 1872.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1921.040 -0.020 1922.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 1971.040 -0.020 1972.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2021.040 -0.020 2022.640 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2021.040 581.160 2022.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2071.040 -0.020 2072.640 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2071.040 581.160 2072.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2121.040 -0.020 2122.640 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2121.040 581.160 2122.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.040 -0.020 2172.640 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.040 581.160 2172.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2221.040 -0.020 2222.640 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2221.040 581.160 2222.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2271.040 -0.020 2272.640 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2271.040 581.160 2272.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2321.040 -0.020 2322.640 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2321.040 581.160 2322.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2371.040 -0.020 2372.640 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2371.040 581.160 2372.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2421.040 -0.020 2422.640 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2421.040 581.160 2422.640 739.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 2471.040 -0.020 2472.640 739.860 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 26.730 2525.260 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 76.730 2525.260 78.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 126.730 2525.260 128.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 176.730 2525.260 178.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 226.730 2525.260 228.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 276.730 2525.260 278.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 326.730 2525.260 328.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 376.730 2525.260 378.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 426.730 2525.260 428.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 476.730 2525.260 478.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 526.730 2525.260 528.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 576.730 2525.260 578.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 626.730 2525.260 628.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 676.730 2525.260 678.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 726.730 2525.260 728.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 2493.780 35.120 2495.380 625.840 ;
    END
  END VPWR
  PIN core_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1385.150 0.000 1385.430 4.000 ;
    END
  END core_clk
  PIN core_rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1468.870 0.000 1469.150 4.000 ;
    END
  END core_rstn
  PIN debug_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 9.560 2520.000 10.160 ;
    END
  END debug_in
  PIN debug_mode
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 20.440 2520.000 21.040 ;
    END
  END debug_mode
  PIN debug_oeb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 31.320 2520.000 31.920 ;
    END
  END debug_oeb
  PIN debug_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 42.200 2520.000 42.800 ;
    END
  END debug_out
  PIN flash_clk
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 597.080 2520.000 597.680 ;
    END
  END flash_clk
  PIN flash_csb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 586.200 2520.000 586.800 ;
    END
  END flash_csb
  PIN flash_io0_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 607.960 2520.000 608.560 ;
    END
  END flash_io0_di
  PIN flash_io0_do
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 618.840 2520.000 619.440 ;
    END
  END flash_io0_do
  PIN flash_io0_oeb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 629.720 2520.000 630.320 ;
    END
  END flash_io0_oeb
  PIN flash_io1_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 640.600 2520.000 641.200 ;
    END
  END flash_io1_di
  PIN flash_io1_do
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 651.480 2520.000 652.080 ;
    END
  END flash_io1_do
  PIN flash_io1_oeb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2516.000 662.360 2520.000 662.960 ;
    END
  END flash_io1_oeb
  PIN flash_io2_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 673.240 2520.000 673.840 ;
    END
  END flash_io2_di
  PIN flash_io2_do
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 684.120 2520.000 684.720 ;
    END
  END flash_io2_do
  PIN flash_io2_oeb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 695.000 2520.000 695.600 ;
    END
  END flash_io2_oeb
  PIN flash_io3_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 705.880 2520.000 706.480 ;
    END
  END flash_io3_di
  PIN flash_io3_do
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 716.760 2520.000 717.360 ;
    END
  END flash_io3_do
  PIN flash_io3_oeb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 727.640 2520.000 728.240 ;
    END
  END flash_io3_oeb
  PIN gpio_in_pad
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1887.470 0.000 1887.750 4.000 ;
    END
  END gpio_in_pad
  PIN gpio_inenb_pad
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1971.190 0.000 1971.470 4.000 ;
    END
  END gpio_inenb_pad
  PIN gpio_mode0_pad
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2054.910 0.000 2055.190 4.000 ;
    END
  END gpio_mode0_pad
  PIN gpio_mode1_pad
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2138.630 0.000 2138.910 4.000 ;
    END
  END gpio_mode1_pad
  PIN gpio_out_pad
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2222.350 0.000 2222.630 4.000 ;
    END
  END gpio_out_pad
  PIN gpio_outenb_pad
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2306.070 0.000 2306.350 4.000 ;
    END
  END gpio_outenb_pad
  PIN hk_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 205.400 2520.000 206.000 ;
    END
  END hk_ack_i
  PIN hk_cyc_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 227.160 2520.000 227.760 ;
    END
  END hk_cyc_o
  PIN hk_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 238.040 2520.000 238.640 ;
    END
  END hk_dat_i[0]
  PIN hk_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 346.840 2520.000 347.440 ;
    END
  END hk_dat_i[10]
  PIN hk_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 357.720 2520.000 358.320 ;
    END
  END hk_dat_i[11]
  PIN hk_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 368.600 2520.000 369.200 ;
    END
  END hk_dat_i[12]
  PIN hk_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 379.480 2520.000 380.080 ;
    END
  END hk_dat_i[13]
  PIN hk_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 390.360 2520.000 390.960 ;
    END
  END hk_dat_i[14]
  PIN hk_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 401.240 2520.000 401.840 ;
    END
  END hk_dat_i[15]
  PIN hk_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 412.120 2520.000 412.720 ;
    END
  END hk_dat_i[16]
  PIN hk_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 423.000 2520.000 423.600 ;
    END
  END hk_dat_i[17]
  PIN hk_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 433.880 2520.000 434.480 ;
    END
  END hk_dat_i[18]
  PIN hk_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 444.760 2520.000 445.360 ;
    END
  END hk_dat_i[19]
  PIN hk_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 248.920 2520.000 249.520 ;
    END
  END hk_dat_i[1]
  PIN hk_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 455.640 2520.000 456.240 ;
    END
  END hk_dat_i[20]
  PIN hk_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 466.520 2520.000 467.120 ;
    END
  END hk_dat_i[21]
  PIN hk_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 477.400 2520.000 478.000 ;
    END
  END hk_dat_i[22]
  PIN hk_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 488.280 2520.000 488.880 ;
    END
  END hk_dat_i[23]
  PIN hk_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 499.160 2520.000 499.760 ;
    END
  END hk_dat_i[24]
  PIN hk_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 510.040 2520.000 510.640 ;
    END
  END hk_dat_i[25]
  PIN hk_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 520.920 2520.000 521.520 ;
    END
  END hk_dat_i[26]
  PIN hk_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 531.800 2520.000 532.400 ;
    END
  END hk_dat_i[27]
  PIN hk_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 542.680 2520.000 543.280 ;
    END
  END hk_dat_i[28]
  PIN hk_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 553.560 2520.000 554.160 ;
    END
  END hk_dat_i[29]
  PIN hk_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 259.800 2520.000 260.400 ;
    END
  END hk_dat_i[2]
  PIN hk_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 564.440 2520.000 565.040 ;
    END
  END hk_dat_i[30]
  PIN hk_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 575.320 2520.000 575.920 ;
    END
  END hk_dat_i[31]
  PIN hk_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 270.680 2520.000 271.280 ;
    END
  END hk_dat_i[3]
  PIN hk_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 281.560 2520.000 282.160 ;
    END
  END hk_dat_i[4]
  PIN hk_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 292.440 2520.000 293.040 ;
    END
  END hk_dat_i[5]
  PIN hk_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 303.320 2520.000 303.920 ;
    END
  END hk_dat_i[6]
  PIN hk_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 314.200 2520.000 314.800 ;
    END
  END hk_dat_i[7]
  PIN hk_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 325.080 2520.000 325.680 ;
    END
  END hk_dat_i[8]
  PIN hk_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 335.960 2520.000 336.560 ;
    END
  END hk_dat_i[9]
  PIN hk_stb_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 216.280 2520.000 216.880 ;
    END
  END hk_stb_o
  PIN irq[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2396.690 736.000 2396.970 740.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2400.370 736.000 2400.650 740.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2404.050 736.000 2404.330 740.000 ;
    END
  END irq[2]
  PIN irq[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 85.720 2520.000 86.320 ;
    END
  END irq[3]
  PIN irq[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 74.840 2520.000 75.440 ;
    END
  END irq[4]
  PIN irq[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 63.960 2520.000 64.560 ;
    END
  END irq[5]
  PIN la_iena[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 115.090 736.000 115.370 740.000 ;
    END
  END la_iena[0]
  PIN la_iena[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1587.090 736.000 1587.370 740.000 ;
    END
  END la_iena[100]
  PIN la_iena[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1601.810 736.000 1602.090 740.000 ;
    END
  END la_iena[101]
  PIN la_iena[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1616.530 736.000 1616.810 740.000 ;
    END
  END la_iena[102]
  PIN la_iena[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1631.250 736.000 1631.530 740.000 ;
    END
  END la_iena[103]
  PIN la_iena[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1645.970 736.000 1646.250 740.000 ;
    END
  END la_iena[104]
  PIN la_iena[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1660.690 736.000 1660.970 740.000 ;
    END
  END la_iena[105]
  PIN la_iena[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1675.410 736.000 1675.690 740.000 ;
    END
  END la_iena[106]
  PIN la_iena[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1690.130 736.000 1690.410 740.000 ;
    END
  END la_iena[107]
  PIN la_iena[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1704.850 736.000 1705.130 740.000 ;
    END
  END la_iena[108]
  PIN la_iena[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1719.570 736.000 1719.850 740.000 ;
    END
  END la_iena[109]
  PIN la_iena[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 262.290 736.000 262.570 740.000 ;
    END
  END la_iena[10]
  PIN la_iena[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1734.290 736.000 1734.570 740.000 ;
    END
  END la_iena[110]
  PIN la_iena[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1749.010 736.000 1749.290 740.000 ;
    END
  END la_iena[111]
  PIN la_iena[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1763.730 736.000 1764.010 740.000 ;
    END
  END la_iena[112]
  PIN la_iena[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1778.450 736.000 1778.730 740.000 ;
    END
  END la_iena[113]
  PIN la_iena[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1793.170 736.000 1793.450 740.000 ;
    END
  END la_iena[114]
  PIN la_iena[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1807.890 736.000 1808.170 740.000 ;
    END
  END la_iena[115]
  PIN la_iena[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1822.610 736.000 1822.890 740.000 ;
    END
  END la_iena[116]
  PIN la_iena[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1837.330 736.000 1837.610 740.000 ;
    END
  END la_iena[117]
  PIN la_iena[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1852.050 736.000 1852.330 740.000 ;
    END
  END la_iena[118]
  PIN la_iena[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1866.770 736.000 1867.050 740.000 ;
    END
  END la_iena[119]
  PIN la_iena[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 277.010 736.000 277.290 740.000 ;
    END
  END la_iena[11]
  PIN la_iena[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1881.490 736.000 1881.770 740.000 ;
    END
  END la_iena[120]
  PIN la_iena[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1896.210 736.000 1896.490 740.000 ;
    END
  END la_iena[121]
  PIN la_iena[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1910.930 736.000 1911.210 740.000 ;
    END
  END la_iena[122]
  PIN la_iena[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1925.650 736.000 1925.930 740.000 ;
    END
  END la_iena[123]
  PIN la_iena[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1940.370 736.000 1940.650 740.000 ;
    END
  END la_iena[124]
  PIN la_iena[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1955.090 736.000 1955.370 740.000 ;
    END
  END la_iena[125]
  PIN la_iena[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1969.810 736.000 1970.090 740.000 ;
    END
  END la_iena[126]
  PIN la_iena[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1984.530 736.000 1984.810 740.000 ;
    END
  END la_iena[127]
  PIN la_iena[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 291.730 736.000 292.010 740.000 ;
    END
  END la_iena[12]
  PIN la_iena[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 306.450 736.000 306.730 740.000 ;
    END
  END la_iena[13]
  PIN la_iena[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 321.170 736.000 321.450 740.000 ;
    END
  END la_iena[14]
  PIN la_iena[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 335.890 736.000 336.170 740.000 ;
    END
  END la_iena[15]
  PIN la_iena[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 350.610 736.000 350.890 740.000 ;
    END
  END la_iena[16]
  PIN la_iena[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 365.330 736.000 365.610 740.000 ;
    END
  END la_iena[17]
  PIN la_iena[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 380.050 736.000 380.330 740.000 ;
    END
  END la_iena[18]
  PIN la_iena[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 394.770 736.000 395.050 740.000 ;
    END
  END la_iena[19]
  PIN la_iena[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 129.810 736.000 130.090 740.000 ;
    END
  END la_iena[1]
  PIN la_iena[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 409.490 736.000 409.770 740.000 ;
    END
  END la_iena[20]
  PIN la_iena[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 424.210 736.000 424.490 740.000 ;
    END
  END la_iena[21]
  PIN la_iena[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 438.930 736.000 439.210 740.000 ;
    END
  END la_iena[22]
  PIN la_iena[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 453.650 736.000 453.930 740.000 ;
    END
  END la_iena[23]
  PIN la_iena[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 468.370 736.000 468.650 740.000 ;
    END
  END la_iena[24]
  PIN la_iena[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 483.090 736.000 483.370 740.000 ;
    END
  END la_iena[25]
  PIN la_iena[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 497.810 736.000 498.090 740.000 ;
    END
  END la_iena[26]
  PIN la_iena[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 512.530 736.000 512.810 740.000 ;
    END
  END la_iena[27]
  PIN la_iena[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 527.250 736.000 527.530 740.000 ;
    END
  END la_iena[28]
  PIN la_iena[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 541.970 736.000 542.250 740.000 ;
    END
  END la_iena[29]
  PIN la_iena[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 144.530 736.000 144.810 740.000 ;
    END
  END la_iena[2]
  PIN la_iena[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 556.690 736.000 556.970 740.000 ;
    END
  END la_iena[30]
  PIN la_iena[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 571.410 736.000 571.690 740.000 ;
    END
  END la_iena[31]
  PIN la_iena[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 586.130 736.000 586.410 740.000 ;
    END
  END la_iena[32]
  PIN la_iena[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 600.850 736.000 601.130 740.000 ;
    END
  END la_iena[33]
  PIN la_iena[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 615.570 736.000 615.850 740.000 ;
    END
  END la_iena[34]
  PIN la_iena[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 630.290 736.000 630.570 740.000 ;
    END
  END la_iena[35]
  PIN la_iena[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 645.010 736.000 645.290 740.000 ;
    END
  END la_iena[36]
  PIN la_iena[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 659.730 736.000 660.010 740.000 ;
    END
  END la_iena[37]
  PIN la_iena[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 674.450 736.000 674.730 740.000 ;
    END
  END la_iena[38]
  PIN la_iena[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 689.170 736.000 689.450 740.000 ;
    END
  END la_iena[39]
  PIN la_iena[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 159.250 736.000 159.530 740.000 ;
    END
  END la_iena[3]
  PIN la_iena[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 703.890 736.000 704.170 740.000 ;
    END
  END la_iena[40]
  PIN la_iena[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 718.610 736.000 718.890 740.000 ;
    END
  END la_iena[41]
  PIN la_iena[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 733.330 736.000 733.610 740.000 ;
    END
  END la_iena[42]
  PIN la_iena[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 748.050 736.000 748.330 740.000 ;
    END
  END la_iena[43]
  PIN la_iena[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 762.770 736.000 763.050 740.000 ;
    END
  END la_iena[44]
  PIN la_iena[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 777.490 736.000 777.770 740.000 ;
    END
  END la_iena[45]
  PIN la_iena[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 792.210 736.000 792.490 740.000 ;
    END
  END la_iena[46]
  PIN la_iena[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 806.930 736.000 807.210 740.000 ;
    END
  END la_iena[47]
  PIN la_iena[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 821.650 736.000 821.930 740.000 ;
    END
  END la_iena[48]
  PIN la_iena[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 836.370 736.000 836.650 740.000 ;
    END
  END la_iena[49]
  PIN la_iena[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 173.970 736.000 174.250 740.000 ;
    END
  END la_iena[4]
  PIN la_iena[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 851.090 736.000 851.370 740.000 ;
    END
  END la_iena[50]
  PIN la_iena[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 865.810 736.000 866.090 740.000 ;
    END
  END la_iena[51]
  PIN la_iena[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 880.530 736.000 880.810 740.000 ;
    END
  END la_iena[52]
  PIN la_iena[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 895.250 736.000 895.530 740.000 ;
    END
  END la_iena[53]
  PIN la_iena[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 909.970 736.000 910.250 740.000 ;
    END
  END la_iena[54]
  PIN la_iena[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 924.690 736.000 924.970 740.000 ;
    END
  END la_iena[55]
  PIN la_iena[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 939.410 736.000 939.690 740.000 ;
    END
  END la_iena[56]
  PIN la_iena[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 954.130 736.000 954.410 740.000 ;
    END
  END la_iena[57]
  PIN la_iena[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 968.850 736.000 969.130 740.000 ;
    END
  END la_iena[58]
  PIN la_iena[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 983.570 736.000 983.850 740.000 ;
    END
  END la_iena[59]
  PIN la_iena[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 188.690 736.000 188.970 740.000 ;
    END
  END la_iena[5]
  PIN la_iena[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 998.290 736.000 998.570 740.000 ;
    END
  END la_iena[60]
  PIN la_iena[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1013.010 736.000 1013.290 740.000 ;
    END
  END la_iena[61]
  PIN la_iena[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1027.730 736.000 1028.010 740.000 ;
    END
  END la_iena[62]
  PIN la_iena[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1042.450 736.000 1042.730 740.000 ;
    END
  END la_iena[63]
  PIN la_iena[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1057.170 736.000 1057.450 740.000 ;
    END
  END la_iena[64]
  PIN la_iena[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1071.890 736.000 1072.170 740.000 ;
    END
  END la_iena[65]
  PIN la_iena[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1086.610 736.000 1086.890 740.000 ;
    END
  END la_iena[66]
  PIN la_iena[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1101.330 736.000 1101.610 740.000 ;
    END
  END la_iena[67]
  PIN la_iena[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1116.050 736.000 1116.330 740.000 ;
    END
  END la_iena[68]
  PIN la_iena[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1130.770 736.000 1131.050 740.000 ;
    END
  END la_iena[69]
  PIN la_iena[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 203.410 736.000 203.690 740.000 ;
    END
  END la_iena[6]
  PIN la_iena[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1145.490 736.000 1145.770 740.000 ;
    END
  END la_iena[70]
  PIN la_iena[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1160.210 736.000 1160.490 740.000 ;
    END
  END la_iena[71]
  PIN la_iena[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1174.930 736.000 1175.210 740.000 ;
    END
  END la_iena[72]
  PIN la_iena[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1189.650 736.000 1189.930 740.000 ;
    END
  END la_iena[73]
  PIN la_iena[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1204.370 736.000 1204.650 740.000 ;
    END
  END la_iena[74]
  PIN la_iena[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1219.090 736.000 1219.370 740.000 ;
    END
  END la_iena[75]
  PIN la_iena[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1233.810 736.000 1234.090 740.000 ;
    END
  END la_iena[76]
  PIN la_iena[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1248.530 736.000 1248.810 740.000 ;
    END
  END la_iena[77]
  PIN la_iena[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1263.250 736.000 1263.530 740.000 ;
    END
  END la_iena[78]
  PIN la_iena[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1277.970 736.000 1278.250 740.000 ;
    END
  END la_iena[79]
  PIN la_iena[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 218.130 736.000 218.410 740.000 ;
    END
  END la_iena[7]
  PIN la_iena[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1292.690 736.000 1292.970 740.000 ;
    END
  END la_iena[80]
  PIN la_iena[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1307.410 736.000 1307.690 740.000 ;
    END
  END la_iena[81]
  PIN la_iena[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1322.130 736.000 1322.410 740.000 ;
    END
  END la_iena[82]
  PIN la_iena[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1336.850 736.000 1337.130 740.000 ;
    END
  END la_iena[83]
  PIN la_iena[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1351.570 736.000 1351.850 740.000 ;
    END
  END la_iena[84]
  PIN la_iena[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1366.290 736.000 1366.570 740.000 ;
    END
  END la_iena[85]
  PIN la_iena[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1381.010 736.000 1381.290 740.000 ;
    END
  END la_iena[86]
  PIN la_iena[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1395.730 736.000 1396.010 740.000 ;
    END
  END la_iena[87]
  PIN la_iena[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1410.450 736.000 1410.730 740.000 ;
    END
  END la_iena[88]
  PIN la_iena[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1425.170 736.000 1425.450 740.000 ;
    END
  END la_iena[89]
  PIN la_iena[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 232.850 736.000 233.130 740.000 ;
    END
  END la_iena[8]
  PIN la_iena[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1439.890 736.000 1440.170 740.000 ;
    END
  END la_iena[90]
  PIN la_iena[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1454.610 736.000 1454.890 740.000 ;
    END
  END la_iena[91]
  PIN la_iena[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1469.330 736.000 1469.610 740.000 ;
    END
  END la_iena[92]
  PIN la_iena[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1484.050 736.000 1484.330 740.000 ;
    END
  END la_iena[93]
  PIN la_iena[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1498.770 736.000 1499.050 740.000 ;
    END
  END la_iena[94]
  PIN la_iena[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1513.490 736.000 1513.770 740.000 ;
    END
  END la_iena[95]
  PIN la_iena[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1528.210 736.000 1528.490 740.000 ;
    END
  END la_iena[96]
  PIN la_iena[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1542.930 736.000 1543.210 740.000 ;
    END
  END la_iena[97]
  PIN la_iena[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1557.650 736.000 1557.930 740.000 ;
    END
  END la_iena[98]
  PIN la_iena[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1572.370 736.000 1572.650 740.000 ;
    END
  END la_iena[99]
  PIN la_iena[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 247.570 736.000 247.850 740.000 ;
    END
  END la_iena[9]
  PIN la_input[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 118.770 736.000 119.050 740.000 ;
    END
  END la_input[0]
  PIN la_input[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1590.770 736.000 1591.050 740.000 ;
    END
  END la_input[100]
  PIN la_input[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1605.490 736.000 1605.770 740.000 ;
    END
  END la_input[101]
  PIN la_input[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1620.210 736.000 1620.490 740.000 ;
    END
  END la_input[102]
  PIN la_input[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1634.930 736.000 1635.210 740.000 ;
    END
  END la_input[103]
  PIN la_input[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1649.650 736.000 1649.930 740.000 ;
    END
  END la_input[104]
  PIN la_input[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1664.370 736.000 1664.650 740.000 ;
    END
  END la_input[105]
  PIN la_input[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1679.090 736.000 1679.370 740.000 ;
    END
  END la_input[106]
  PIN la_input[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1693.810 736.000 1694.090 740.000 ;
    END
  END la_input[107]
  PIN la_input[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1708.530 736.000 1708.810 740.000 ;
    END
  END la_input[108]
  PIN la_input[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1723.250 736.000 1723.530 740.000 ;
    END
  END la_input[109]
  PIN la_input[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 265.970 736.000 266.250 740.000 ;
    END
  END la_input[10]
  PIN la_input[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1737.970 736.000 1738.250 740.000 ;
    END
  END la_input[110]
  PIN la_input[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1752.690 736.000 1752.970 740.000 ;
    END
  END la_input[111]
  PIN la_input[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1767.410 736.000 1767.690 740.000 ;
    END
  END la_input[112]
  PIN la_input[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1782.130 736.000 1782.410 740.000 ;
    END
  END la_input[113]
  PIN la_input[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1796.850 736.000 1797.130 740.000 ;
    END
  END la_input[114]
  PIN la_input[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1811.570 736.000 1811.850 740.000 ;
    END
  END la_input[115]
  PIN la_input[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1826.290 736.000 1826.570 740.000 ;
    END
  END la_input[116]
  PIN la_input[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1841.010 736.000 1841.290 740.000 ;
    END
  END la_input[117]
  PIN la_input[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1855.730 736.000 1856.010 740.000 ;
    END
  END la_input[118]
  PIN la_input[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1870.450 736.000 1870.730 740.000 ;
    END
  END la_input[119]
  PIN la_input[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 280.690 736.000 280.970 740.000 ;
    END
  END la_input[11]
  PIN la_input[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1885.170 736.000 1885.450 740.000 ;
    END
  END la_input[120]
  PIN la_input[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1899.890 736.000 1900.170 740.000 ;
    END
  END la_input[121]
  PIN la_input[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1914.610 736.000 1914.890 740.000 ;
    END
  END la_input[122]
  PIN la_input[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1929.330 736.000 1929.610 740.000 ;
    END
  END la_input[123]
  PIN la_input[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1944.050 736.000 1944.330 740.000 ;
    END
  END la_input[124]
  PIN la_input[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1958.770 736.000 1959.050 740.000 ;
    END
  END la_input[125]
  PIN la_input[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1973.490 736.000 1973.770 740.000 ;
    END
  END la_input[126]
  PIN la_input[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1988.210 736.000 1988.490 740.000 ;
    END
  END la_input[127]
  PIN la_input[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 295.410 736.000 295.690 740.000 ;
    END
  END la_input[12]
  PIN la_input[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 310.130 736.000 310.410 740.000 ;
    END
  END la_input[13]
  PIN la_input[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 324.850 736.000 325.130 740.000 ;
    END
  END la_input[14]
  PIN la_input[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 339.570 736.000 339.850 740.000 ;
    END
  END la_input[15]
  PIN la_input[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 354.290 736.000 354.570 740.000 ;
    END
  END la_input[16]
  PIN la_input[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 369.010 736.000 369.290 740.000 ;
    END
  END la_input[17]
  PIN la_input[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 383.730 736.000 384.010 740.000 ;
    END
  END la_input[18]
  PIN la_input[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 398.450 736.000 398.730 740.000 ;
    END
  END la_input[19]
  PIN la_input[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 133.490 736.000 133.770 740.000 ;
    END
  END la_input[1]
  PIN la_input[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 413.170 736.000 413.450 740.000 ;
    END
  END la_input[20]
  PIN la_input[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 427.890 736.000 428.170 740.000 ;
    END
  END la_input[21]
  PIN la_input[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 442.610 736.000 442.890 740.000 ;
    END
  END la_input[22]
  PIN la_input[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 457.330 736.000 457.610 740.000 ;
    END
  END la_input[23]
  PIN la_input[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 472.050 736.000 472.330 740.000 ;
    END
  END la_input[24]
  PIN la_input[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 486.770 736.000 487.050 740.000 ;
    END
  END la_input[25]
  PIN la_input[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 501.490 736.000 501.770 740.000 ;
    END
  END la_input[26]
  PIN la_input[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 516.210 736.000 516.490 740.000 ;
    END
  END la_input[27]
  PIN la_input[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 530.930 736.000 531.210 740.000 ;
    END
  END la_input[28]
  PIN la_input[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 545.650 736.000 545.930 740.000 ;
    END
  END la_input[29]
  PIN la_input[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 148.210 736.000 148.490 740.000 ;
    END
  END la_input[2]
  PIN la_input[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 560.370 736.000 560.650 740.000 ;
    END
  END la_input[30]
  PIN la_input[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 575.090 736.000 575.370 740.000 ;
    END
  END la_input[31]
  PIN la_input[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 589.810 736.000 590.090 740.000 ;
    END
  END la_input[32]
  PIN la_input[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 604.530 736.000 604.810 740.000 ;
    END
  END la_input[33]
  PIN la_input[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 619.250 736.000 619.530 740.000 ;
    END
  END la_input[34]
  PIN la_input[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 633.970 736.000 634.250 740.000 ;
    END
  END la_input[35]
  PIN la_input[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 648.690 736.000 648.970 740.000 ;
    END
  END la_input[36]
  PIN la_input[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 663.410 736.000 663.690 740.000 ;
    END
  END la_input[37]
  PIN la_input[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 678.130 736.000 678.410 740.000 ;
    END
  END la_input[38]
  PIN la_input[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 692.850 736.000 693.130 740.000 ;
    END
  END la_input[39]
  PIN la_input[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 162.930 736.000 163.210 740.000 ;
    END
  END la_input[3]
  PIN la_input[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 707.570 736.000 707.850 740.000 ;
    END
  END la_input[40]
  PIN la_input[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 722.290 736.000 722.570 740.000 ;
    END
  END la_input[41]
  PIN la_input[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 737.010 736.000 737.290 740.000 ;
    END
  END la_input[42]
  PIN la_input[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 751.730 736.000 752.010 740.000 ;
    END
  END la_input[43]
  PIN la_input[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 766.450 736.000 766.730 740.000 ;
    END
  END la_input[44]
  PIN la_input[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 781.170 736.000 781.450 740.000 ;
    END
  END la_input[45]
  PIN la_input[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 795.890 736.000 796.170 740.000 ;
    END
  END la_input[46]
  PIN la_input[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 810.610 736.000 810.890 740.000 ;
    END
  END la_input[47]
  PIN la_input[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 825.330 736.000 825.610 740.000 ;
    END
  END la_input[48]
  PIN la_input[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 840.050 736.000 840.330 740.000 ;
    END
  END la_input[49]
  PIN la_input[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 177.650 736.000 177.930 740.000 ;
    END
  END la_input[4]
  PIN la_input[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 854.770 736.000 855.050 740.000 ;
    END
  END la_input[50]
  PIN la_input[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 869.490 736.000 869.770 740.000 ;
    END
  END la_input[51]
  PIN la_input[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 884.210 736.000 884.490 740.000 ;
    END
  END la_input[52]
  PIN la_input[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 898.930 736.000 899.210 740.000 ;
    END
  END la_input[53]
  PIN la_input[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 913.650 736.000 913.930 740.000 ;
    END
  END la_input[54]
  PIN la_input[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 928.370 736.000 928.650 740.000 ;
    END
  END la_input[55]
  PIN la_input[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 943.090 736.000 943.370 740.000 ;
    END
  END la_input[56]
  PIN la_input[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 957.810 736.000 958.090 740.000 ;
    END
  END la_input[57]
  PIN la_input[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 972.530 736.000 972.810 740.000 ;
    END
  END la_input[58]
  PIN la_input[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 987.250 736.000 987.530 740.000 ;
    END
  END la_input[59]
  PIN la_input[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 192.370 736.000 192.650 740.000 ;
    END
  END la_input[5]
  PIN la_input[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1001.970 736.000 1002.250 740.000 ;
    END
  END la_input[60]
  PIN la_input[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1016.690 736.000 1016.970 740.000 ;
    END
  END la_input[61]
  PIN la_input[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1031.410 736.000 1031.690 740.000 ;
    END
  END la_input[62]
  PIN la_input[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1046.130 736.000 1046.410 740.000 ;
    END
  END la_input[63]
  PIN la_input[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1060.850 736.000 1061.130 740.000 ;
    END
  END la_input[64]
  PIN la_input[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1075.570 736.000 1075.850 740.000 ;
    END
  END la_input[65]
  PIN la_input[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1090.290 736.000 1090.570 740.000 ;
    END
  END la_input[66]
  PIN la_input[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1105.010 736.000 1105.290 740.000 ;
    END
  END la_input[67]
  PIN la_input[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1119.730 736.000 1120.010 740.000 ;
    END
  END la_input[68]
  PIN la_input[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1134.450 736.000 1134.730 740.000 ;
    END
  END la_input[69]
  PIN la_input[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 207.090 736.000 207.370 740.000 ;
    END
  END la_input[6]
  PIN la_input[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1149.170 736.000 1149.450 740.000 ;
    END
  END la_input[70]
  PIN la_input[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1163.890 736.000 1164.170 740.000 ;
    END
  END la_input[71]
  PIN la_input[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1178.610 736.000 1178.890 740.000 ;
    END
  END la_input[72]
  PIN la_input[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1193.330 736.000 1193.610 740.000 ;
    END
  END la_input[73]
  PIN la_input[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1208.050 736.000 1208.330 740.000 ;
    END
  END la_input[74]
  PIN la_input[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1222.770 736.000 1223.050 740.000 ;
    END
  END la_input[75]
  PIN la_input[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1237.490 736.000 1237.770 740.000 ;
    END
  END la_input[76]
  PIN la_input[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1252.210 736.000 1252.490 740.000 ;
    END
  END la_input[77]
  PIN la_input[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1266.930 736.000 1267.210 740.000 ;
    END
  END la_input[78]
  PIN la_input[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1281.650 736.000 1281.930 740.000 ;
    END
  END la_input[79]
  PIN la_input[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 221.810 736.000 222.090 740.000 ;
    END
  END la_input[7]
  PIN la_input[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1296.370 736.000 1296.650 740.000 ;
    END
  END la_input[80]
  PIN la_input[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1311.090 736.000 1311.370 740.000 ;
    END
  END la_input[81]
  PIN la_input[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1325.810 736.000 1326.090 740.000 ;
    END
  END la_input[82]
  PIN la_input[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1340.530 736.000 1340.810 740.000 ;
    END
  END la_input[83]
  PIN la_input[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1355.250 736.000 1355.530 740.000 ;
    END
  END la_input[84]
  PIN la_input[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1369.970 736.000 1370.250 740.000 ;
    END
  END la_input[85]
  PIN la_input[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1384.690 736.000 1384.970 740.000 ;
    END
  END la_input[86]
  PIN la_input[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1399.410 736.000 1399.690 740.000 ;
    END
  END la_input[87]
  PIN la_input[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1414.130 736.000 1414.410 740.000 ;
    END
  END la_input[88]
  PIN la_input[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1428.850 736.000 1429.130 740.000 ;
    END
  END la_input[89]
  PIN la_input[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 236.530 736.000 236.810 740.000 ;
    END
  END la_input[8]
  PIN la_input[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1443.570 736.000 1443.850 740.000 ;
    END
  END la_input[90]
  PIN la_input[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1458.290 736.000 1458.570 740.000 ;
    END
  END la_input[91]
  PIN la_input[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1473.010 736.000 1473.290 740.000 ;
    END
  END la_input[92]
  PIN la_input[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1487.730 736.000 1488.010 740.000 ;
    END
  END la_input[93]
  PIN la_input[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1502.450 736.000 1502.730 740.000 ;
    END
  END la_input[94]
  PIN la_input[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1517.170 736.000 1517.450 740.000 ;
    END
  END la_input[95]
  PIN la_input[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1531.890 736.000 1532.170 740.000 ;
    END
  END la_input[96]
  PIN la_input[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1546.610 736.000 1546.890 740.000 ;
    END
  END la_input[97]
  PIN la_input[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1561.330 736.000 1561.610 740.000 ;
    END
  END la_input[98]
  PIN la_input[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1576.050 736.000 1576.330 740.000 ;
    END
  END la_input[99]
  PIN la_input[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 251.250 736.000 251.530 740.000 ;
    END
  END la_input[9]
  PIN la_oenb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 122.450 736.000 122.730 740.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1594.450 736.000 1594.730 740.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1609.170 736.000 1609.450 740.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1623.890 736.000 1624.170 740.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1638.610 736.000 1638.890 740.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1653.330 736.000 1653.610 740.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1668.050 736.000 1668.330 740.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1682.770 736.000 1683.050 740.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1697.490 736.000 1697.770 740.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1712.210 736.000 1712.490 740.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1726.930 736.000 1727.210 740.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 269.650 736.000 269.930 740.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1741.650 736.000 1741.930 740.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1756.370 736.000 1756.650 740.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1771.090 736.000 1771.370 740.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1785.810 736.000 1786.090 740.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1800.530 736.000 1800.810 740.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1815.250 736.000 1815.530 740.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1829.970 736.000 1830.250 740.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1844.690 736.000 1844.970 740.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1859.410 736.000 1859.690 740.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1874.130 736.000 1874.410 740.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 284.370 736.000 284.650 740.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1888.850 736.000 1889.130 740.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1903.570 736.000 1903.850 740.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1918.290 736.000 1918.570 740.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1933.010 736.000 1933.290 740.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1947.730 736.000 1948.010 740.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1962.450 736.000 1962.730 740.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1977.170 736.000 1977.450 740.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1991.890 736.000 1992.170 740.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 299.090 736.000 299.370 740.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 313.810 736.000 314.090 740.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 328.530 736.000 328.810 740.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 343.250 736.000 343.530 740.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 357.970 736.000 358.250 740.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 372.690 736.000 372.970 740.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 387.410 736.000 387.690 740.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 402.130 736.000 402.410 740.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 137.170 736.000 137.450 740.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 416.850 736.000 417.130 740.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 431.570 736.000 431.850 740.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 446.290 736.000 446.570 740.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 461.010 736.000 461.290 740.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 475.730 736.000 476.010 740.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 490.450 736.000 490.730 740.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 505.170 736.000 505.450 740.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 519.890 736.000 520.170 740.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 534.610 736.000 534.890 740.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 549.330 736.000 549.610 740.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 151.890 736.000 152.170 740.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 564.050 736.000 564.330 740.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 578.770 736.000 579.050 740.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 593.490 736.000 593.770 740.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 608.210 736.000 608.490 740.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 622.930 736.000 623.210 740.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 637.650 736.000 637.930 740.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 652.370 736.000 652.650 740.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 667.090 736.000 667.370 740.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 681.810 736.000 682.090 740.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 696.530 736.000 696.810 740.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 166.610 736.000 166.890 740.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 711.250 736.000 711.530 740.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 725.970 736.000 726.250 740.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 740.690 736.000 740.970 740.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 755.410 736.000 755.690 740.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 770.130 736.000 770.410 740.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 784.850 736.000 785.130 740.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 799.570 736.000 799.850 740.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 814.290 736.000 814.570 740.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 829.010 736.000 829.290 740.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 843.730 736.000 844.010 740.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 181.330 736.000 181.610 740.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 858.450 736.000 858.730 740.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 873.170 736.000 873.450 740.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 887.890 736.000 888.170 740.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 902.610 736.000 902.890 740.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 917.330 736.000 917.610 740.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 932.050 736.000 932.330 740.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 946.770 736.000 947.050 740.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 961.490 736.000 961.770 740.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 976.210 736.000 976.490 740.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 990.930 736.000 991.210 740.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 196.050 736.000 196.330 740.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1005.650 736.000 1005.930 740.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1020.370 736.000 1020.650 740.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1035.090 736.000 1035.370 740.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1049.810 736.000 1050.090 740.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1064.530 736.000 1064.810 740.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1079.250 736.000 1079.530 740.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1093.970 736.000 1094.250 740.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1108.690 736.000 1108.970 740.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1123.410 736.000 1123.690 740.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1138.130 736.000 1138.410 740.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 210.770 736.000 211.050 740.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1152.850 736.000 1153.130 740.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1167.570 736.000 1167.850 740.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1182.290 736.000 1182.570 740.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1197.010 736.000 1197.290 740.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1211.730 736.000 1212.010 740.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1226.450 736.000 1226.730 740.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1241.170 736.000 1241.450 740.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1255.890 736.000 1256.170 740.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1270.610 736.000 1270.890 740.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1285.330 736.000 1285.610 740.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 225.490 736.000 225.770 740.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1300.050 736.000 1300.330 740.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1314.770 736.000 1315.050 740.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1329.490 736.000 1329.770 740.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1344.210 736.000 1344.490 740.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1358.930 736.000 1359.210 740.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1373.650 736.000 1373.930 740.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1388.370 736.000 1388.650 740.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1403.090 736.000 1403.370 740.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1417.810 736.000 1418.090 740.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1432.530 736.000 1432.810 740.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 240.210 736.000 240.490 740.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1447.250 736.000 1447.530 740.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1461.970 736.000 1462.250 740.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1476.690 736.000 1476.970 740.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1491.410 736.000 1491.690 740.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1506.130 736.000 1506.410 740.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1520.850 736.000 1521.130 740.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1535.570 736.000 1535.850 740.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1550.290 736.000 1550.570 740.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1565.010 736.000 1565.290 740.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1579.730 736.000 1580.010 740.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 254.930 736.000 255.210 740.000 ;
    END
  END la_oenb[9]
  PIN la_output[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 126.130 736.000 126.410 740.000 ;
    END
  END la_output[0]
  PIN la_output[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1598.130 736.000 1598.410 740.000 ;
    END
  END la_output[100]
  PIN la_output[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1612.850 736.000 1613.130 740.000 ;
    END
  END la_output[101]
  PIN la_output[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1627.570 736.000 1627.850 740.000 ;
    END
  END la_output[102]
  PIN la_output[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1642.290 736.000 1642.570 740.000 ;
    END
  END la_output[103]
  PIN la_output[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1657.010 736.000 1657.290 740.000 ;
    END
  END la_output[104]
  PIN la_output[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1671.730 736.000 1672.010 740.000 ;
    END
  END la_output[105]
  PIN la_output[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1686.450 736.000 1686.730 740.000 ;
    END
  END la_output[106]
  PIN la_output[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1701.170 736.000 1701.450 740.000 ;
    END
  END la_output[107]
  PIN la_output[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1715.890 736.000 1716.170 740.000 ;
    END
  END la_output[108]
  PIN la_output[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1730.610 736.000 1730.890 740.000 ;
    END
  END la_output[109]
  PIN la_output[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 273.330 736.000 273.610 740.000 ;
    END
  END la_output[10]
  PIN la_output[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1745.330 736.000 1745.610 740.000 ;
    END
  END la_output[110]
  PIN la_output[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1760.050 736.000 1760.330 740.000 ;
    END
  END la_output[111]
  PIN la_output[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1774.770 736.000 1775.050 740.000 ;
    END
  END la_output[112]
  PIN la_output[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1789.490 736.000 1789.770 740.000 ;
    END
  END la_output[113]
  PIN la_output[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1804.210 736.000 1804.490 740.000 ;
    END
  END la_output[114]
  PIN la_output[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1818.930 736.000 1819.210 740.000 ;
    END
  END la_output[115]
  PIN la_output[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1833.650 736.000 1833.930 740.000 ;
    END
  END la_output[116]
  PIN la_output[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1848.370 736.000 1848.650 740.000 ;
    END
  END la_output[117]
  PIN la_output[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1863.090 736.000 1863.370 740.000 ;
    END
  END la_output[118]
  PIN la_output[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1877.810 736.000 1878.090 740.000 ;
    END
  END la_output[119]
  PIN la_output[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 288.050 736.000 288.330 740.000 ;
    END
  END la_output[11]
  PIN la_output[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1892.530 736.000 1892.810 740.000 ;
    END
  END la_output[120]
  PIN la_output[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1907.250 736.000 1907.530 740.000 ;
    END
  END la_output[121]
  PIN la_output[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1921.970 736.000 1922.250 740.000 ;
    END
  END la_output[122]
  PIN la_output[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1936.690 736.000 1936.970 740.000 ;
    END
  END la_output[123]
  PIN la_output[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1951.410 736.000 1951.690 740.000 ;
    END
  END la_output[124]
  PIN la_output[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1966.130 736.000 1966.410 740.000 ;
    END
  END la_output[125]
  PIN la_output[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1980.850 736.000 1981.130 740.000 ;
    END
  END la_output[126]
  PIN la_output[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1995.570 736.000 1995.850 740.000 ;
    END
  END la_output[127]
  PIN la_output[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 302.770 736.000 303.050 740.000 ;
    END
  END la_output[12]
  PIN la_output[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 317.490 736.000 317.770 740.000 ;
    END
  END la_output[13]
  PIN la_output[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 332.210 736.000 332.490 740.000 ;
    END
  END la_output[14]
  PIN la_output[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 346.930 736.000 347.210 740.000 ;
    END
  END la_output[15]
  PIN la_output[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 361.650 736.000 361.930 740.000 ;
    END
  END la_output[16]
  PIN la_output[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 376.370 736.000 376.650 740.000 ;
    END
  END la_output[17]
  PIN la_output[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 391.090 736.000 391.370 740.000 ;
    END
  END la_output[18]
  PIN la_output[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 405.810 736.000 406.090 740.000 ;
    END
  END la_output[19]
  PIN la_output[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 140.850 736.000 141.130 740.000 ;
    END
  END la_output[1]
  PIN la_output[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 420.530 736.000 420.810 740.000 ;
    END
  END la_output[20]
  PIN la_output[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 435.250 736.000 435.530 740.000 ;
    END
  END la_output[21]
  PIN la_output[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 449.970 736.000 450.250 740.000 ;
    END
  END la_output[22]
  PIN la_output[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 464.690 736.000 464.970 740.000 ;
    END
  END la_output[23]
  PIN la_output[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 479.410 736.000 479.690 740.000 ;
    END
  END la_output[24]
  PIN la_output[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 494.130 736.000 494.410 740.000 ;
    END
  END la_output[25]
  PIN la_output[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 508.850 736.000 509.130 740.000 ;
    END
  END la_output[26]
  PIN la_output[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 523.570 736.000 523.850 740.000 ;
    END
  END la_output[27]
  PIN la_output[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 538.290 736.000 538.570 740.000 ;
    END
  END la_output[28]
  PIN la_output[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 553.010 736.000 553.290 740.000 ;
    END
  END la_output[29]
  PIN la_output[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 155.570 736.000 155.850 740.000 ;
    END
  END la_output[2]
  PIN la_output[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 567.730 736.000 568.010 740.000 ;
    END
  END la_output[30]
  PIN la_output[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 582.450 736.000 582.730 740.000 ;
    END
  END la_output[31]
  PIN la_output[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 597.170 736.000 597.450 740.000 ;
    END
  END la_output[32]
  PIN la_output[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 611.890 736.000 612.170 740.000 ;
    END
  END la_output[33]
  PIN la_output[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 626.610 736.000 626.890 740.000 ;
    END
  END la_output[34]
  PIN la_output[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 641.330 736.000 641.610 740.000 ;
    END
  END la_output[35]
  PIN la_output[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 656.050 736.000 656.330 740.000 ;
    END
  END la_output[36]
  PIN la_output[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 670.770 736.000 671.050 740.000 ;
    END
  END la_output[37]
  PIN la_output[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 685.490 736.000 685.770 740.000 ;
    END
  END la_output[38]
  PIN la_output[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 700.210 736.000 700.490 740.000 ;
    END
  END la_output[39]
  PIN la_output[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 170.290 736.000 170.570 740.000 ;
    END
  END la_output[3]
  PIN la_output[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 714.930 736.000 715.210 740.000 ;
    END
  END la_output[40]
  PIN la_output[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 729.650 736.000 729.930 740.000 ;
    END
  END la_output[41]
  PIN la_output[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 744.370 736.000 744.650 740.000 ;
    END
  END la_output[42]
  PIN la_output[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 759.090 736.000 759.370 740.000 ;
    END
  END la_output[43]
  PIN la_output[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 773.810 736.000 774.090 740.000 ;
    END
  END la_output[44]
  PIN la_output[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 788.530 736.000 788.810 740.000 ;
    END
  END la_output[45]
  PIN la_output[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 803.250 736.000 803.530 740.000 ;
    END
  END la_output[46]
  PIN la_output[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 817.970 736.000 818.250 740.000 ;
    END
  END la_output[47]
  PIN la_output[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 832.690 736.000 832.970 740.000 ;
    END
  END la_output[48]
  PIN la_output[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 847.410 736.000 847.690 740.000 ;
    END
  END la_output[49]
  PIN la_output[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 185.010 736.000 185.290 740.000 ;
    END
  END la_output[4]
  PIN la_output[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 862.130 736.000 862.410 740.000 ;
    END
  END la_output[50]
  PIN la_output[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 876.850 736.000 877.130 740.000 ;
    END
  END la_output[51]
  PIN la_output[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 891.570 736.000 891.850 740.000 ;
    END
  END la_output[52]
  PIN la_output[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 906.290 736.000 906.570 740.000 ;
    END
  END la_output[53]
  PIN la_output[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 921.010 736.000 921.290 740.000 ;
    END
  END la_output[54]
  PIN la_output[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 935.730 736.000 936.010 740.000 ;
    END
  END la_output[55]
  PIN la_output[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 950.450 736.000 950.730 740.000 ;
    END
  END la_output[56]
  PIN la_output[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 965.170 736.000 965.450 740.000 ;
    END
  END la_output[57]
  PIN la_output[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 979.890 736.000 980.170 740.000 ;
    END
  END la_output[58]
  PIN la_output[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 994.610 736.000 994.890 740.000 ;
    END
  END la_output[59]
  PIN la_output[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 199.730 736.000 200.010 740.000 ;
    END
  END la_output[5]
  PIN la_output[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1009.330 736.000 1009.610 740.000 ;
    END
  END la_output[60]
  PIN la_output[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1024.050 736.000 1024.330 740.000 ;
    END
  END la_output[61]
  PIN la_output[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1038.770 736.000 1039.050 740.000 ;
    END
  END la_output[62]
  PIN la_output[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1053.490 736.000 1053.770 740.000 ;
    END
  END la_output[63]
  PIN la_output[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1068.210 736.000 1068.490 740.000 ;
    END
  END la_output[64]
  PIN la_output[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1082.930 736.000 1083.210 740.000 ;
    END
  END la_output[65]
  PIN la_output[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1097.650 736.000 1097.930 740.000 ;
    END
  END la_output[66]
  PIN la_output[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1112.370 736.000 1112.650 740.000 ;
    END
  END la_output[67]
  PIN la_output[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1127.090 736.000 1127.370 740.000 ;
    END
  END la_output[68]
  PIN la_output[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1141.810 736.000 1142.090 740.000 ;
    END
  END la_output[69]
  PIN la_output[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 214.450 736.000 214.730 740.000 ;
    END
  END la_output[6]
  PIN la_output[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1156.530 736.000 1156.810 740.000 ;
    END
  END la_output[70]
  PIN la_output[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1171.250 736.000 1171.530 740.000 ;
    END
  END la_output[71]
  PIN la_output[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1185.970 736.000 1186.250 740.000 ;
    END
  END la_output[72]
  PIN la_output[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1200.690 736.000 1200.970 740.000 ;
    END
  END la_output[73]
  PIN la_output[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1215.410 736.000 1215.690 740.000 ;
    END
  END la_output[74]
  PIN la_output[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1230.130 736.000 1230.410 740.000 ;
    END
  END la_output[75]
  PIN la_output[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1244.850 736.000 1245.130 740.000 ;
    END
  END la_output[76]
  PIN la_output[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1259.570 736.000 1259.850 740.000 ;
    END
  END la_output[77]
  PIN la_output[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1274.290 736.000 1274.570 740.000 ;
    END
  END la_output[78]
  PIN la_output[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1289.010 736.000 1289.290 740.000 ;
    END
  END la_output[79]
  PIN la_output[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 229.170 736.000 229.450 740.000 ;
    END
  END la_output[7]
  PIN la_output[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1303.730 736.000 1304.010 740.000 ;
    END
  END la_output[80]
  PIN la_output[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1318.450 736.000 1318.730 740.000 ;
    END
  END la_output[81]
  PIN la_output[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1333.170 736.000 1333.450 740.000 ;
    END
  END la_output[82]
  PIN la_output[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1347.890 736.000 1348.170 740.000 ;
    END
  END la_output[83]
  PIN la_output[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1362.610 736.000 1362.890 740.000 ;
    END
  END la_output[84]
  PIN la_output[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1377.330 736.000 1377.610 740.000 ;
    END
  END la_output[85]
  PIN la_output[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1392.050 736.000 1392.330 740.000 ;
    END
  END la_output[86]
  PIN la_output[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1406.770 736.000 1407.050 740.000 ;
    END
  END la_output[87]
  PIN la_output[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1421.490 736.000 1421.770 740.000 ;
    END
  END la_output[88]
  PIN la_output[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1436.210 736.000 1436.490 740.000 ;
    END
  END la_output[89]
  PIN la_output[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 243.890 736.000 244.170 740.000 ;
    END
  END la_output[8]
  PIN la_output[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1450.930 736.000 1451.210 740.000 ;
    END
  END la_output[90]
  PIN la_output[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1465.650 736.000 1465.930 740.000 ;
    END
  END la_output[91]
  PIN la_output[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1480.370 736.000 1480.650 740.000 ;
    END
  END la_output[92]
  PIN la_output[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1495.090 736.000 1495.370 740.000 ;
    END
  END la_output[93]
  PIN la_output[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1509.810 736.000 1510.090 740.000 ;
    END
  END la_output[94]
  PIN la_output[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1524.530 736.000 1524.810 740.000 ;
    END
  END la_output[95]
  PIN la_output[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1539.250 736.000 1539.530 740.000 ;
    END
  END la_output[96]
  PIN la_output[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1553.970 736.000 1554.250 740.000 ;
    END
  END la_output[97]
  PIN la_output[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1568.690 736.000 1568.970 740.000 ;
    END
  END la_output[98]
  PIN la_output[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1583.410 736.000 1583.690 740.000 ;
    END
  END la_output[99]
  PIN la_output[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 258.610 736.000 258.890 740.000 ;
    END
  END la_output[9]
  PIN mprj_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1999.250 736.000 1999.530 740.000 ;
    END
  END mprj_ack_i
  PIN mprj_adr_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 2017.650 736.000 2017.930 740.000 ;
    END
  END mprj_adr_o[0]
  PIN mprj_adr_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2142.770 736.000 2143.050 740.000 ;
    END
  END mprj_adr_o[10]
  PIN mprj_adr_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2153.810 736.000 2154.090 740.000 ;
    END
  END mprj_adr_o[11]
  PIN mprj_adr_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2164.850 736.000 2165.130 740.000 ;
    END
  END mprj_adr_o[12]
  PIN mprj_adr_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2175.890 736.000 2176.170 740.000 ;
    END
  END mprj_adr_o[13]
  PIN mprj_adr_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2186.930 736.000 2187.210 740.000 ;
    END
  END mprj_adr_o[14]
  PIN mprj_adr_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2197.970 736.000 2198.250 740.000 ;
    END
  END mprj_adr_o[15]
  PIN mprj_adr_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2209.010 736.000 2209.290 740.000 ;
    END
  END mprj_adr_o[16]
  PIN mprj_adr_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2220.050 736.000 2220.330 740.000 ;
    END
  END mprj_adr_o[17]
  PIN mprj_adr_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2231.090 736.000 2231.370 740.000 ;
    END
  END mprj_adr_o[18]
  PIN mprj_adr_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2242.130 736.000 2242.410 740.000 ;
    END
  END mprj_adr_o[19]
  PIN mprj_adr_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 2032.370 736.000 2032.650 740.000 ;
    END
  END mprj_adr_o[1]
  PIN mprj_adr_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2253.170 736.000 2253.450 740.000 ;
    END
  END mprj_adr_o[20]
  PIN mprj_adr_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2264.210 736.000 2264.490 740.000 ;
    END
  END mprj_adr_o[21]
  PIN mprj_adr_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2275.250 736.000 2275.530 740.000 ;
    END
  END mprj_adr_o[22]
  PIN mprj_adr_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2286.290 736.000 2286.570 740.000 ;
    END
  END mprj_adr_o[23]
  PIN mprj_adr_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2297.330 736.000 2297.610 740.000 ;
    END
  END mprj_adr_o[24]
  PIN mprj_adr_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2308.370 736.000 2308.650 740.000 ;
    END
  END mprj_adr_o[25]
  PIN mprj_adr_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2319.410 736.000 2319.690 740.000 ;
    END
  END mprj_adr_o[26]
  PIN mprj_adr_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2330.450 736.000 2330.730 740.000 ;
    END
  END mprj_adr_o[27]
  PIN mprj_adr_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2341.490 736.000 2341.770 740.000 ;
    END
  END mprj_adr_o[28]
  PIN mprj_adr_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2352.530 736.000 2352.810 740.000 ;
    END
  END mprj_adr_o[29]
  PIN mprj_adr_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2047.090 736.000 2047.370 740.000 ;
    END
  END mprj_adr_o[2]
  PIN mprj_adr_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2363.570 736.000 2363.850 740.000 ;
    END
  END mprj_adr_o[30]
  PIN mprj_adr_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2374.610 736.000 2374.890 740.000 ;
    END
  END mprj_adr_o[31]
  PIN mprj_adr_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2061.810 736.000 2062.090 740.000 ;
    END
  END mprj_adr_o[3]
  PIN mprj_adr_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2076.530 736.000 2076.810 740.000 ;
    END
  END mprj_adr_o[4]
  PIN mprj_adr_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2087.570 736.000 2087.850 740.000 ;
    END
  END mprj_adr_o[5]
  PIN mprj_adr_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2098.610 736.000 2098.890 740.000 ;
    END
  END mprj_adr_o[6]
  PIN mprj_adr_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2109.650 736.000 2109.930 740.000 ;
    END
  END mprj_adr_o[7]
  PIN mprj_adr_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2120.690 736.000 2120.970 740.000 ;
    END
  END mprj_adr_o[8]
  PIN mprj_adr_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2131.730 736.000 2132.010 740.000 ;
    END
  END mprj_adr_o[9]
  PIN mprj_cyc_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2002.930 736.000 2003.210 740.000 ;
    END
  END mprj_cyc_o
  PIN mprj_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2021.330 736.000 2021.610 740.000 ;
    END
  END mprj_dat_i[0]
  PIN mprj_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2146.450 736.000 2146.730 740.000 ;
    END
  END mprj_dat_i[10]
  PIN mprj_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2157.490 736.000 2157.770 740.000 ;
    END
  END mprj_dat_i[11]
  PIN mprj_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2168.530 736.000 2168.810 740.000 ;
    END
  END mprj_dat_i[12]
  PIN mprj_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2179.570 736.000 2179.850 740.000 ;
    END
  END mprj_dat_i[13]
  PIN mprj_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2190.610 736.000 2190.890 740.000 ;
    END
  END mprj_dat_i[14]
  PIN mprj_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2201.650 736.000 2201.930 740.000 ;
    END
  END mprj_dat_i[15]
  PIN mprj_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2212.690 736.000 2212.970 740.000 ;
    END
  END mprj_dat_i[16]
  PIN mprj_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2223.730 736.000 2224.010 740.000 ;
    END
  END mprj_dat_i[17]
  PIN mprj_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2234.770 736.000 2235.050 740.000 ;
    END
  END mprj_dat_i[18]
  PIN mprj_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2245.810 736.000 2246.090 740.000 ;
    END
  END mprj_dat_i[19]
  PIN mprj_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2036.050 736.000 2036.330 740.000 ;
    END
  END mprj_dat_i[1]
  PIN mprj_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2256.850 736.000 2257.130 740.000 ;
    END
  END mprj_dat_i[20]
  PIN mprj_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2267.890 736.000 2268.170 740.000 ;
    END
  END mprj_dat_i[21]
  PIN mprj_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2278.930 736.000 2279.210 740.000 ;
    END
  END mprj_dat_i[22]
  PIN mprj_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2289.970 736.000 2290.250 740.000 ;
    END
  END mprj_dat_i[23]
  PIN mprj_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2301.010 736.000 2301.290 740.000 ;
    END
  END mprj_dat_i[24]
  PIN mprj_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2312.050 736.000 2312.330 740.000 ;
    END
  END mprj_dat_i[25]
  PIN mprj_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2323.090 736.000 2323.370 740.000 ;
    END
  END mprj_dat_i[26]
  PIN mprj_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2334.130 736.000 2334.410 740.000 ;
    END
  END mprj_dat_i[27]
  PIN mprj_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2345.170 736.000 2345.450 740.000 ;
    END
  END mprj_dat_i[28]
  PIN mprj_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2356.210 736.000 2356.490 740.000 ;
    END
  END mprj_dat_i[29]
  PIN mprj_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2050.770 736.000 2051.050 740.000 ;
    END
  END mprj_dat_i[2]
  PIN mprj_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2367.250 736.000 2367.530 740.000 ;
    END
  END mprj_dat_i[30]
  PIN mprj_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2378.290 736.000 2378.570 740.000 ;
    END
  END mprj_dat_i[31]
  PIN mprj_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2065.490 736.000 2065.770 740.000 ;
    END
  END mprj_dat_i[3]
  PIN mprj_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2080.210 736.000 2080.490 740.000 ;
    END
  END mprj_dat_i[4]
  PIN mprj_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2091.250 736.000 2091.530 740.000 ;
    END
  END mprj_dat_i[5]
  PIN mprj_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2102.290 736.000 2102.570 740.000 ;
    END
  END mprj_dat_i[6]
  PIN mprj_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2113.330 736.000 2113.610 740.000 ;
    END
  END mprj_dat_i[7]
  PIN mprj_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2124.370 736.000 2124.650 740.000 ;
    END
  END mprj_dat_i[8]
  PIN mprj_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2135.410 736.000 2135.690 740.000 ;
    END
  END mprj_dat_i[9]
  PIN mprj_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2025.010 736.000 2025.290 740.000 ;
    END
  END mprj_dat_o[0]
  PIN mprj_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2150.130 736.000 2150.410 740.000 ;
    END
  END mprj_dat_o[10]
  PIN mprj_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2161.170 736.000 2161.450 740.000 ;
    END
  END mprj_dat_o[11]
  PIN mprj_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2172.210 736.000 2172.490 740.000 ;
    END
  END mprj_dat_o[12]
  PIN mprj_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2183.250 736.000 2183.530 740.000 ;
    END
  END mprj_dat_o[13]
  PIN mprj_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2194.290 736.000 2194.570 740.000 ;
    END
  END mprj_dat_o[14]
  PIN mprj_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2205.330 736.000 2205.610 740.000 ;
    END
  END mprj_dat_o[15]
  PIN mprj_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2216.370 736.000 2216.650 740.000 ;
    END
  END mprj_dat_o[16]
  PIN mprj_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2227.410 736.000 2227.690 740.000 ;
    END
  END mprj_dat_o[17]
  PIN mprj_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2238.450 736.000 2238.730 740.000 ;
    END
  END mprj_dat_o[18]
  PIN mprj_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2249.490 736.000 2249.770 740.000 ;
    END
  END mprj_dat_o[19]
  PIN mprj_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2039.730 736.000 2040.010 740.000 ;
    END
  END mprj_dat_o[1]
  PIN mprj_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2260.530 736.000 2260.810 740.000 ;
    END
  END mprj_dat_o[20]
  PIN mprj_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2271.570 736.000 2271.850 740.000 ;
    END
  END mprj_dat_o[21]
  PIN mprj_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2282.610 736.000 2282.890 740.000 ;
    END
  END mprj_dat_o[22]
  PIN mprj_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2293.650 736.000 2293.930 740.000 ;
    END
  END mprj_dat_o[23]
  PIN mprj_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2304.690 736.000 2304.970 740.000 ;
    END
  END mprj_dat_o[24]
  PIN mprj_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2315.730 736.000 2316.010 740.000 ;
    END
  END mprj_dat_o[25]
  PIN mprj_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2326.770 736.000 2327.050 740.000 ;
    END
  END mprj_dat_o[26]
  PIN mprj_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2337.810 736.000 2338.090 740.000 ;
    END
  END mprj_dat_o[27]
  PIN mprj_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2348.850 736.000 2349.130 740.000 ;
    END
  END mprj_dat_o[28]
  PIN mprj_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2359.890 736.000 2360.170 740.000 ;
    END
  END mprj_dat_o[29]
  PIN mprj_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2054.450 736.000 2054.730 740.000 ;
    END
  END mprj_dat_o[2]
  PIN mprj_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2370.930 736.000 2371.210 740.000 ;
    END
  END mprj_dat_o[30]
  PIN mprj_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2381.970 736.000 2382.250 740.000 ;
    END
  END mprj_dat_o[31]
  PIN mprj_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2069.170 736.000 2069.450 740.000 ;
    END
  END mprj_dat_o[3]
  PIN mprj_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2083.890 736.000 2084.170 740.000 ;
    END
  END mprj_dat_o[4]
  PIN mprj_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2094.930 736.000 2095.210 740.000 ;
    END
  END mprj_dat_o[5]
  PIN mprj_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2105.970 736.000 2106.250 740.000 ;
    END
  END mprj_dat_o[6]
  PIN mprj_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2117.010 736.000 2117.290 740.000 ;
    END
  END mprj_dat_o[7]
  PIN mprj_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2128.050 736.000 2128.330 740.000 ;
    END
  END mprj_dat_o[8]
  PIN mprj_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2139.090 736.000 2139.370 740.000 ;
    END
  END mprj_dat_o[9]
  PIN mprj_sel_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2028.690 736.000 2028.970 740.000 ;
    END
  END mprj_sel_o[0]
  PIN mprj_sel_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2043.410 736.000 2043.690 740.000 ;
    END
  END mprj_sel_o[1]
  PIN mprj_sel_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2058.130 736.000 2058.410 740.000 ;
    END
  END mprj_sel_o[2]
  PIN mprj_sel_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2072.850 736.000 2073.130 740.000 ;
    END
  END mprj_sel_o[3]
  PIN mprj_stb_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2006.610 736.000 2006.890 740.000 ;
    END
  END mprj_stb_o
  PIN mprj_wb_iena
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2010.290 736.000 2010.570 740.000 ;
    END
  END mprj_wb_iena
  PIN mprj_we_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2013.970 736.000 2014.250 740.000 ;
    END
  END mprj_we_o
  PIN qspi_enabled
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 194.520 2520.000 195.120 ;
    END
  END qspi_enabled
  PIN ser_rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 151.000 2520.000 151.600 ;
    END
  END ser_rx
  PIN ser_tx
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 161.880 2520.000 162.480 ;
    END
  END ser_tx
  PIN spi_csb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 129.240 2520.000 129.840 ;
    END
  END spi_csb
  PIN spi_enabled
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 172.760 2520.000 173.360 ;
    END
  END spi_enabled
  PIN spi_sck
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 118.360 2520.000 118.960 ;
    END
  END spi_sck
  PIN spi_sdi
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 140.120 2520.000 140.720 ;
    END
  END spi_sdi
  PIN spi_sdo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 107.480 2520.000 108.080 ;
    END
  END spi_sdo
  PIN spi_sdoenb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 96.600 2520.000 97.200 ;
    END
  END spi_sdoenb
  PIN tck
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END tck
  PIN tdi
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END tdi
  PIN tdo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.800 4.000 430.400 ;
    END
  END tdo
  PIN tdo_paden_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 674.600 4.000 675.200 ;
    END
  END tdo_paden_o
  PIN tms
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.746000 ;
    ANTENNADIFFAREA 3.477600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END tms
  PIN trap
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2516.000 53.080 2520.000 53.680 ;
    END
  END trap
  PIN trst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.200 4.000 552.800 ;
    END
  END trst
  PIN uart_enabled
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 2516.000 183.640 2520.000 184.240 ;
    END
  END uart_enabled
  PIN user_irq_ena[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2385.650 736.000 2385.930 740.000 ;
    END
  END user_irq_ena[0]
  PIN user_irq_ena[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2389.330 736.000 2389.610 740.000 ;
    END
  END user_irq_ena[1]
  PIN user_irq_ena[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 2393.010 736.000 2393.290 740.000 ;
    END
  END user_irq_ena[2]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2514.360 729.045 ;
      LAYER met1 ;
        RECT 5.520 1.060 2519.810 733.680 ;
      LAYER met2 ;
        RECT 6.070 735.720 114.810 736.170 ;
        RECT 115.650 735.720 118.490 736.170 ;
        RECT 119.330 735.720 122.170 736.170 ;
        RECT 123.010 735.720 125.850 736.170 ;
        RECT 126.690 735.720 129.530 736.170 ;
        RECT 130.370 735.720 133.210 736.170 ;
        RECT 134.050 735.720 136.890 736.170 ;
        RECT 137.730 735.720 140.570 736.170 ;
        RECT 141.410 735.720 144.250 736.170 ;
        RECT 145.090 735.720 147.930 736.170 ;
        RECT 148.770 735.720 151.610 736.170 ;
        RECT 152.450 735.720 155.290 736.170 ;
        RECT 156.130 735.720 158.970 736.170 ;
        RECT 159.810 735.720 162.650 736.170 ;
        RECT 163.490 735.720 166.330 736.170 ;
        RECT 167.170 735.720 170.010 736.170 ;
        RECT 170.850 735.720 173.690 736.170 ;
        RECT 174.530 735.720 177.370 736.170 ;
        RECT 178.210 735.720 181.050 736.170 ;
        RECT 181.890 735.720 184.730 736.170 ;
        RECT 185.570 735.720 188.410 736.170 ;
        RECT 189.250 735.720 192.090 736.170 ;
        RECT 192.930 735.720 195.770 736.170 ;
        RECT 196.610 735.720 199.450 736.170 ;
        RECT 200.290 735.720 203.130 736.170 ;
        RECT 203.970 735.720 206.810 736.170 ;
        RECT 207.650 735.720 210.490 736.170 ;
        RECT 211.330 735.720 214.170 736.170 ;
        RECT 215.010 735.720 217.850 736.170 ;
        RECT 218.690 735.720 221.530 736.170 ;
        RECT 222.370 735.720 225.210 736.170 ;
        RECT 226.050 735.720 228.890 736.170 ;
        RECT 229.730 735.720 232.570 736.170 ;
        RECT 233.410 735.720 236.250 736.170 ;
        RECT 237.090 735.720 239.930 736.170 ;
        RECT 240.770 735.720 243.610 736.170 ;
        RECT 244.450 735.720 247.290 736.170 ;
        RECT 248.130 735.720 250.970 736.170 ;
        RECT 251.810 735.720 254.650 736.170 ;
        RECT 255.490 735.720 258.330 736.170 ;
        RECT 259.170 735.720 262.010 736.170 ;
        RECT 262.850 735.720 265.690 736.170 ;
        RECT 266.530 735.720 269.370 736.170 ;
        RECT 270.210 735.720 273.050 736.170 ;
        RECT 273.890 735.720 276.730 736.170 ;
        RECT 277.570 735.720 280.410 736.170 ;
        RECT 281.250 735.720 284.090 736.170 ;
        RECT 284.930 735.720 287.770 736.170 ;
        RECT 288.610 735.720 291.450 736.170 ;
        RECT 292.290 735.720 295.130 736.170 ;
        RECT 295.970 735.720 298.810 736.170 ;
        RECT 299.650 735.720 302.490 736.170 ;
        RECT 303.330 735.720 306.170 736.170 ;
        RECT 307.010 735.720 309.850 736.170 ;
        RECT 310.690 735.720 313.530 736.170 ;
        RECT 314.370 735.720 317.210 736.170 ;
        RECT 318.050 735.720 320.890 736.170 ;
        RECT 321.730 735.720 324.570 736.170 ;
        RECT 325.410 735.720 328.250 736.170 ;
        RECT 329.090 735.720 331.930 736.170 ;
        RECT 332.770 735.720 335.610 736.170 ;
        RECT 336.450 735.720 339.290 736.170 ;
        RECT 340.130 735.720 342.970 736.170 ;
        RECT 343.810 735.720 346.650 736.170 ;
        RECT 347.490 735.720 350.330 736.170 ;
        RECT 351.170 735.720 354.010 736.170 ;
        RECT 354.850 735.720 357.690 736.170 ;
        RECT 358.530 735.720 361.370 736.170 ;
        RECT 362.210 735.720 365.050 736.170 ;
        RECT 365.890 735.720 368.730 736.170 ;
        RECT 369.570 735.720 372.410 736.170 ;
        RECT 373.250 735.720 376.090 736.170 ;
        RECT 376.930 735.720 379.770 736.170 ;
        RECT 380.610 735.720 383.450 736.170 ;
        RECT 384.290 735.720 387.130 736.170 ;
        RECT 387.970 735.720 390.810 736.170 ;
        RECT 391.650 735.720 394.490 736.170 ;
        RECT 395.330 735.720 398.170 736.170 ;
        RECT 399.010 735.720 401.850 736.170 ;
        RECT 402.690 735.720 405.530 736.170 ;
        RECT 406.370 735.720 409.210 736.170 ;
        RECT 410.050 735.720 412.890 736.170 ;
        RECT 413.730 735.720 416.570 736.170 ;
        RECT 417.410 735.720 420.250 736.170 ;
        RECT 421.090 735.720 423.930 736.170 ;
        RECT 424.770 735.720 427.610 736.170 ;
        RECT 428.450 735.720 431.290 736.170 ;
        RECT 432.130 735.720 434.970 736.170 ;
        RECT 435.810 735.720 438.650 736.170 ;
        RECT 439.490 735.720 442.330 736.170 ;
        RECT 443.170 735.720 446.010 736.170 ;
        RECT 446.850 735.720 449.690 736.170 ;
        RECT 450.530 735.720 453.370 736.170 ;
        RECT 454.210 735.720 457.050 736.170 ;
        RECT 457.890 735.720 460.730 736.170 ;
        RECT 461.570 735.720 464.410 736.170 ;
        RECT 465.250 735.720 468.090 736.170 ;
        RECT 468.930 735.720 471.770 736.170 ;
        RECT 472.610 735.720 475.450 736.170 ;
        RECT 476.290 735.720 479.130 736.170 ;
        RECT 479.970 735.720 482.810 736.170 ;
        RECT 483.650 735.720 486.490 736.170 ;
        RECT 487.330 735.720 490.170 736.170 ;
        RECT 491.010 735.720 493.850 736.170 ;
        RECT 494.690 735.720 497.530 736.170 ;
        RECT 498.370 735.720 501.210 736.170 ;
        RECT 502.050 735.720 504.890 736.170 ;
        RECT 505.730 735.720 508.570 736.170 ;
        RECT 509.410 735.720 512.250 736.170 ;
        RECT 513.090 735.720 515.930 736.170 ;
        RECT 516.770 735.720 519.610 736.170 ;
        RECT 520.450 735.720 523.290 736.170 ;
        RECT 524.130 735.720 526.970 736.170 ;
        RECT 527.810 735.720 530.650 736.170 ;
        RECT 531.490 735.720 534.330 736.170 ;
        RECT 535.170 735.720 538.010 736.170 ;
        RECT 538.850 735.720 541.690 736.170 ;
        RECT 542.530 735.720 545.370 736.170 ;
        RECT 546.210 735.720 549.050 736.170 ;
        RECT 549.890 735.720 552.730 736.170 ;
        RECT 553.570 735.720 556.410 736.170 ;
        RECT 557.250 735.720 560.090 736.170 ;
        RECT 560.930 735.720 563.770 736.170 ;
        RECT 564.610 735.720 567.450 736.170 ;
        RECT 568.290 735.720 571.130 736.170 ;
        RECT 571.970 735.720 574.810 736.170 ;
        RECT 575.650 735.720 578.490 736.170 ;
        RECT 579.330 735.720 582.170 736.170 ;
        RECT 583.010 735.720 585.850 736.170 ;
        RECT 586.690 735.720 589.530 736.170 ;
        RECT 590.370 735.720 593.210 736.170 ;
        RECT 594.050 735.720 596.890 736.170 ;
        RECT 597.730 735.720 600.570 736.170 ;
        RECT 601.410 735.720 604.250 736.170 ;
        RECT 605.090 735.720 607.930 736.170 ;
        RECT 608.770 735.720 611.610 736.170 ;
        RECT 612.450 735.720 615.290 736.170 ;
        RECT 616.130 735.720 618.970 736.170 ;
        RECT 619.810 735.720 622.650 736.170 ;
        RECT 623.490 735.720 626.330 736.170 ;
        RECT 627.170 735.720 630.010 736.170 ;
        RECT 630.850 735.720 633.690 736.170 ;
        RECT 634.530 735.720 637.370 736.170 ;
        RECT 638.210 735.720 641.050 736.170 ;
        RECT 641.890 735.720 644.730 736.170 ;
        RECT 645.570 735.720 648.410 736.170 ;
        RECT 649.250 735.720 652.090 736.170 ;
        RECT 652.930 735.720 655.770 736.170 ;
        RECT 656.610 735.720 659.450 736.170 ;
        RECT 660.290 735.720 663.130 736.170 ;
        RECT 663.970 735.720 666.810 736.170 ;
        RECT 667.650 735.720 670.490 736.170 ;
        RECT 671.330 735.720 674.170 736.170 ;
        RECT 675.010 735.720 677.850 736.170 ;
        RECT 678.690 735.720 681.530 736.170 ;
        RECT 682.370 735.720 685.210 736.170 ;
        RECT 686.050 735.720 688.890 736.170 ;
        RECT 689.730 735.720 692.570 736.170 ;
        RECT 693.410 735.720 696.250 736.170 ;
        RECT 697.090 735.720 699.930 736.170 ;
        RECT 700.770 735.720 703.610 736.170 ;
        RECT 704.450 735.720 707.290 736.170 ;
        RECT 708.130 735.720 710.970 736.170 ;
        RECT 711.810 735.720 714.650 736.170 ;
        RECT 715.490 735.720 718.330 736.170 ;
        RECT 719.170 735.720 722.010 736.170 ;
        RECT 722.850 735.720 725.690 736.170 ;
        RECT 726.530 735.720 729.370 736.170 ;
        RECT 730.210 735.720 733.050 736.170 ;
        RECT 733.890 735.720 736.730 736.170 ;
        RECT 737.570 735.720 740.410 736.170 ;
        RECT 741.250 735.720 744.090 736.170 ;
        RECT 744.930 735.720 747.770 736.170 ;
        RECT 748.610 735.720 751.450 736.170 ;
        RECT 752.290 735.720 755.130 736.170 ;
        RECT 755.970 735.720 758.810 736.170 ;
        RECT 759.650 735.720 762.490 736.170 ;
        RECT 763.330 735.720 766.170 736.170 ;
        RECT 767.010 735.720 769.850 736.170 ;
        RECT 770.690 735.720 773.530 736.170 ;
        RECT 774.370 735.720 777.210 736.170 ;
        RECT 778.050 735.720 780.890 736.170 ;
        RECT 781.730 735.720 784.570 736.170 ;
        RECT 785.410 735.720 788.250 736.170 ;
        RECT 789.090 735.720 791.930 736.170 ;
        RECT 792.770 735.720 795.610 736.170 ;
        RECT 796.450 735.720 799.290 736.170 ;
        RECT 800.130 735.720 802.970 736.170 ;
        RECT 803.810 735.720 806.650 736.170 ;
        RECT 807.490 735.720 810.330 736.170 ;
        RECT 811.170 735.720 814.010 736.170 ;
        RECT 814.850 735.720 817.690 736.170 ;
        RECT 818.530 735.720 821.370 736.170 ;
        RECT 822.210 735.720 825.050 736.170 ;
        RECT 825.890 735.720 828.730 736.170 ;
        RECT 829.570 735.720 832.410 736.170 ;
        RECT 833.250 735.720 836.090 736.170 ;
        RECT 836.930 735.720 839.770 736.170 ;
        RECT 840.610 735.720 843.450 736.170 ;
        RECT 844.290 735.720 847.130 736.170 ;
        RECT 847.970 735.720 850.810 736.170 ;
        RECT 851.650 735.720 854.490 736.170 ;
        RECT 855.330 735.720 858.170 736.170 ;
        RECT 859.010 735.720 861.850 736.170 ;
        RECT 862.690 735.720 865.530 736.170 ;
        RECT 866.370 735.720 869.210 736.170 ;
        RECT 870.050 735.720 872.890 736.170 ;
        RECT 873.730 735.720 876.570 736.170 ;
        RECT 877.410 735.720 880.250 736.170 ;
        RECT 881.090 735.720 883.930 736.170 ;
        RECT 884.770 735.720 887.610 736.170 ;
        RECT 888.450 735.720 891.290 736.170 ;
        RECT 892.130 735.720 894.970 736.170 ;
        RECT 895.810 735.720 898.650 736.170 ;
        RECT 899.490 735.720 902.330 736.170 ;
        RECT 903.170 735.720 906.010 736.170 ;
        RECT 906.850 735.720 909.690 736.170 ;
        RECT 910.530 735.720 913.370 736.170 ;
        RECT 914.210 735.720 917.050 736.170 ;
        RECT 917.890 735.720 920.730 736.170 ;
        RECT 921.570 735.720 924.410 736.170 ;
        RECT 925.250 735.720 928.090 736.170 ;
        RECT 928.930 735.720 931.770 736.170 ;
        RECT 932.610 735.720 935.450 736.170 ;
        RECT 936.290 735.720 939.130 736.170 ;
        RECT 939.970 735.720 942.810 736.170 ;
        RECT 943.650 735.720 946.490 736.170 ;
        RECT 947.330 735.720 950.170 736.170 ;
        RECT 951.010 735.720 953.850 736.170 ;
        RECT 954.690 735.720 957.530 736.170 ;
        RECT 958.370 735.720 961.210 736.170 ;
        RECT 962.050 735.720 964.890 736.170 ;
        RECT 965.730 735.720 968.570 736.170 ;
        RECT 969.410 735.720 972.250 736.170 ;
        RECT 973.090 735.720 975.930 736.170 ;
        RECT 976.770 735.720 979.610 736.170 ;
        RECT 980.450 735.720 983.290 736.170 ;
        RECT 984.130 735.720 986.970 736.170 ;
        RECT 987.810 735.720 990.650 736.170 ;
        RECT 991.490 735.720 994.330 736.170 ;
        RECT 995.170 735.720 998.010 736.170 ;
        RECT 998.850 735.720 1001.690 736.170 ;
        RECT 1002.530 735.720 1005.370 736.170 ;
        RECT 1006.210 735.720 1009.050 736.170 ;
        RECT 1009.890 735.720 1012.730 736.170 ;
        RECT 1013.570 735.720 1016.410 736.170 ;
        RECT 1017.250 735.720 1020.090 736.170 ;
        RECT 1020.930 735.720 1023.770 736.170 ;
        RECT 1024.610 735.720 1027.450 736.170 ;
        RECT 1028.290 735.720 1031.130 736.170 ;
        RECT 1031.970 735.720 1034.810 736.170 ;
        RECT 1035.650 735.720 1038.490 736.170 ;
        RECT 1039.330 735.720 1042.170 736.170 ;
        RECT 1043.010 735.720 1045.850 736.170 ;
        RECT 1046.690 735.720 1049.530 736.170 ;
        RECT 1050.370 735.720 1053.210 736.170 ;
        RECT 1054.050 735.720 1056.890 736.170 ;
        RECT 1057.730 735.720 1060.570 736.170 ;
        RECT 1061.410 735.720 1064.250 736.170 ;
        RECT 1065.090 735.720 1067.930 736.170 ;
        RECT 1068.770 735.720 1071.610 736.170 ;
        RECT 1072.450 735.720 1075.290 736.170 ;
        RECT 1076.130 735.720 1078.970 736.170 ;
        RECT 1079.810 735.720 1082.650 736.170 ;
        RECT 1083.490 735.720 1086.330 736.170 ;
        RECT 1087.170 735.720 1090.010 736.170 ;
        RECT 1090.850 735.720 1093.690 736.170 ;
        RECT 1094.530 735.720 1097.370 736.170 ;
        RECT 1098.210 735.720 1101.050 736.170 ;
        RECT 1101.890 735.720 1104.730 736.170 ;
        RECT 1105.570 735.720 1108.410 736.170 ;
        RECT 1109.250 735.720 1112.090 736.170 ;
        RECT 1112.930 735.720 1115.770 736.170 ;
        RECT 1116.610 735.720 1119.450 736.170 ;
        RECT 1120.290 735.720 1123.130 736.170 ;
        RECT 1123.970 735.720 1126.810 736.170 ;
        RECT 1127.650 735.720 1130.490 736.170 ;
        RECT 1131.330 735.720 1134.170 736.170 ;
        RECT 1135.010 735.720 1137.850 736.170 ;
        RECT 1138.690 735.720 1141.530 736.170 ;
        RECT 1142.370 735.720 1145.210 736.170 ;
        RECT 1146.050 735.720 1148.890 736.170 ;
        RECT 1149.730 735.720 1152.570 736.170 ;
        RECT 1153.410 735.720 1156.250 736.170 ;
        RECT 1157.090 735.720 1159.930 736.170 ;
        RECT 1160.770 735.720 1163.610 736.170 ;
        RECT 1164.450 735.720 1167.290 736.170 ;
        RECT 1168.130 735.720 1170.970 736.170 ;
        RECT 1171.810 735.720 1174.650 736.170 ;
        RECT 1175.490 735.720 1178.330 736.170 ;
        RECT 1179.170 735.720 1182.010 736.170 ;
        RECT 1182.850 735.720 1185.690 736.170 ;
        RECT 1186.530 735.720 1189.370 736.170 ;
        RECT 1190.210 735.720 1193.050 736.170 ;
        RECT 1193.890 735.720 1196.730 736.170 ;
        RECT 1197.570 735.720 1200.410 736.170 ;
        RECT 1201.250 735.720 1204.090 736.170 ;
        RECT 1204.930 735.720 1207.770 736.170 ;
        RECT 1208.610 735.720 1211.450 736.170 ;
        RECT 1212.290 735.720 1215.130 736.170 ;
        RECT 1215.970 735.720 1218.810 736.170 ;
        RECT 1219.650 735.720 1222.490 736.170 ;
        RECT 1223.330 735.720 1226.170 736.170 ;
        RECT 1227.010 735.720 1229.850 736.170 ;
        RECT 1230.690 735.720 1233.530 736.170 ;
        RECT 1234.370 735.720 1237.210 736.170 ;
        RECT 1238.050 735.720 1240.890 736.170 ;
        RECT 1241.730 735.720 1244.570 736.170 ;
        RECT 1245.410 735.720 1248.250 736.170 ;
        RECT 1249.090 735.720 1251.930 736.170 ;
        RECT 1252.770 735.720 1255.610 736.170 ;
        RECT 1256.450 735.720 1259.290 736.170 ;
        RECT 1260.130 735.720 1262.970 736.170 ;
        RECT 1263.810 735.720 1266.650 736.170 ;
        RECT 1267.490 735.720 1270.330 736.170 ;
        RECT 1271.170 735.720 1274.010 736.170 ;
        RECT 1274.850 735.720 1277.690 736.170 ;
        RECT 1278.530 735.720 1281.370 736.170 ;
        RECT 1282.210 735.720 1285.050 736.170 ;
        RECT 1285.890 735.720 1288.730 736.170 ;
        RECT 1289.570 735.720 1292.410 736.170 ;
        RECT 1293.250 735.720 1296.090 736.170 ;
        RECT 1296.930 735.720 1299.770 736.170 ;
        RECT 1300.610 735.720 1303.450 736.170 ;
        RECT 1304.290 735.720 1307.130 736.170 ;
        RECT 1307.970 735.720 1310.810 736.170 ;
        RECT 1311.650 735.720 1314.490 736.170 ;
        RECT 1315.330 735.720 1318.170 736.170 ;
        RECT 1319.010 735.720 1321.850 736.170 ;
        RECT 1322.690 735.720 1325.530 736.170 ;
        RECT 1326.370 735.720 1329.210 736.170 ;
        RECT 1330.050 735.720 1332.890 736.170 ;
        RECT 1333.730 735.720 1336.570 736.170 ;
        RECT 1337.410 735.720 1340.250 736.170 ;
        RECT 1341.090 735.720 1343.930 736.170 ;
        RECT 1344.770 735.720 1347.610 736.170 ;
        RECT 1348.450 735.720 1351.290 736.170 ;
        RECT 1352.130 735.720 1354.970 736.170 ;
        RECT 1355.810 735.720 1358.650 736.170 ;
        RECT 1359.490 735.720 1362.330 736.170 ;
        RECT 1363.170 735.720 1366.010 736.170 ;
        RECT 1366.850 735.720 1369.690 736.170 ;
        RECT 1370.530 735.720 1373.370 736.170 ;
        RECT 1374.210 735.720 1377.050 736.170 ;
        RECT 1377.890 735.720 1380.730 736.170 ;
        RECT 1381.570 735.720 1384.410 736.170 ;
        RECT 1385.250 735.720 1388.090 736.170 ;
        RECT 1388.930 735.720 1391.770 736.170 ;
        RECT 1392.610 735.720 1395.450 736.170 ;
        RECT 1396.290 735.720 1399.130 736.170 ;
        RECT 1399.970 735.720 1402.810 736.170 ;
        RECT 1403.650 735.720 1406.490 736.170 ;
        RECT 1407.330 735.720 1410.170 736.170 ;
        RECT 1411.010 735.720 1413.850 736.170 ;
        RECT 1414.690 735.720 1417.530 736.170 ;
        RECT 1418.370 735.720 1421.210 736.170 ;
        RECT 1422.050 735.720 1424.890 736.170 ;
        RECT 1425.730 735.720 1428.570 736.170 ;
        RECT 1429.410 735.720 1432.250 736.170 ;
        RECT 1433.090 735.720 1435.930 736.170 ;
        RECT 1436.770 735.720 1439.610 736.170 ;
        RECT 1440.450 735.720 1443.290 736.170 ;
        RECT 1444.130 735.720 1446.970 736.170 ;
        RECT 1447.810 735.720 1450.650 736.170 ;
        RECT 1451.490 735.720 1454.330 736.170 ;
        RECT 1455.170 735.720 1458.010 736.170 ;
        RECT 1458.850 735.720 1461.690 736.170 ;
        RECT 1462.530 735.720 1465.370 736.170 ;
        RECT 1466.210 735.720 1469.050 736.170 ;
        RECT 1469.890 735.720 1472.730 736.170 ;
        RECT 1473.570 735.720 1476.410 736.170 ;
        RECT 1477.250 735.720 1480.090 736.170 ;
        RECT 1480.930 735.720 1483.770 736.170 ;
        RECT 1484.610 735.720 1487.450 736.170 ;
        RECT 1488.290 735.720 1491.130 736.170 ;
        RECT 1491.970 735.720 1494.810 736.170 ;
        RECT 1495.650 735.720 1498.490 736.170 ;
        RECT 1499.330 735.720 1502.170 736.170 ;
        RECT 1503.010 735.720 1505.850 736.170 ;
        RECT 1506.690 735.720 1509.530 736.170 ;
        RECT 1510.370 735.720 1513.210 736.170 ;
        RECT 1514.050 735.720 1516.890 736.170 ;
        RECT 1517.730 735.720 1520.570 736.170 ;
        RECT 1521.410 735.720 1524.250 736.170 ;
        RECT 1525.090 735.720 1527.930 736.170 ;
        RECT 1528.770 735.720 1531.610 736.170 ;
        RECT 1532.450 735.720 1535.290 736.170 ;
        RECT 1536.130 735.720 1538.970 736.170 ;
        RECT 1539.810 735.720 1542.650 736.170 ;
        RECT 1543.490 735.720 1546.330 736.170 ;
        RECT 1547.170 735.720 1550.010 736.170 ;
        RECT 1550.850 735.720 1553.690 736.170 ;
        RECT 1554.530 735.720 1557.370 736.170 ;
        RECT 1558.210 735.720 1561.050 736.170 ;
        RECT 1561.890 735.720 1564.730 736.170 ;
        RECT 1565.570 735.720 1568.410 736.170 ;
        RECT 1569.250 735.720 1572.090 736.170 ;
        RECT 1572.930 735.720 1575.770 736.170 ;
        RECT 1576.610 735.720 1579.450 736.170 ;
        RECT 1580.290 735.720 1583.130 736.170 ;
        RECT 1583.970 735.720 1586.810 736.170 ;
        RECT 1587.650 735.720 1590.490 736.170 ;
        RECT 1591.330 735.720 1594.170 736.170 ;
        RECT 1595.010 735.720 1597.850 736.170 ;
        RECT 1598.690 735.720 1601.530 736.170 ;
        RECT 1602.370 735.720 1605.210 736.170 ;
        RECT 1606.050 735.720 1608.890 736.170 ;
        RECT 1609.730 735.720 1612.570 736.170 ;
        RECT 1613.410 735.720 1616.250 736.170 ;
        RECT 1617.090 735.720 1619.930 736.170 ;
        RECT 1620.770 735.720 1623.610 736.170 ;
        RECT 1624.450 735.720 1627.290 736.170 ;
        RECT 1628.130 735.720 1630.970 736.170 ;
        RECT 1631.810 735.720 1634.650 736.170 ;
        RECT 1635.490 735.720 1638.330 736.170 ;
        RECT 1639.170 735.720 1642.010 736.170 ;
        RECT 1642.850 735.720 1645.690 736.170 ;
        RECT 1646.530 735.720 1649.370 736.170 ;
        RECT 1650.210 735.720 1653.050 736.170 ;
        RECT 1653.890 735.720 1656.730 736.170 ;
        RECT 1657.570 735.720 1660.410 736.170 ;
        RECT 1661.250 735.720 1664.090 736.170 ;
        RECT 1664.930 735.720 1667.770 736.170 ;
        RECT 1668.610 735.720 1671.450 736.170 ;
        RECT 1672.290 735.720 1675.130 736.170 ;
        RECT 1675.970 735.720 1678.810 736.170 ;
        RECT 1679.650 735.720 1682.490 736.170 ;
        RECT 1683.330 735.720 1686.170 736.170 ;
        RECT 1687.010 735.720 1689.850 736.170 ;
        RECT 1690.690 735.720 1693.530 736.170 ;
        RECT 1694.370 735.720 1697.210 736.170 ;
        RECT 1698.050 735.720 1700.890 736.170 ;
        RECT 1701.730 735.720 1704.570 736.170 ;
        RECT 1705.410 735.720 1708.250 736.170 ;
        RECT 1709.090 735.720 1711.930 736.170 ;
        RECT 1712.770 735.720 1715.610 736.170 ;
        RECT 1716.450 735.720 1719.290 736.170 ;
        RECT 1720.130 735.720 1722.970 736.170 ;
        RECT 1723.810 735.720 1726.650 736.170 ;
        RECT 1727.490 735.720 1730.330 736.170 ;
        RECT 1731.170 735.720 1734.010 736.170 ;
        RECT 1734.850 735.720 1737.690 736.170 ;
        RECT 1738.530 735.720 1741.370 736.170 ;
        RECT 1742.210 735.720 1745.050 736.170 ;
        RECT 1745.890 735.720 1748.730 736.170 ;
        RECT 1749.570 735.720 1752.410 736.170 ;
        RECT 1753.250 735.720 1756.090 736.170 ;
        RECT 1756.930 735.720 1759.770 736.170 ;
        RECT 1760.610 735.720 1763.450 736.170 ;
        RECT 1764.290 735.720 1767.130 736.170 ;
        RECT 1767.970 735.720 1770.810 736.170 ;
        RECT 1771.650 735.720 1774.490 736.170 ;
        RECT 1775.330 735.720 1778.170 736.170 ;
        RECT 1779.010 735.720 1781.850 736.170 ;
        RECT 1782.690 735.720 1785.530 736.170 ;
        RECT 1786.370 735.720 1789.210 736.170 ;
        RECT 1790.050 735.720 1792.890 736.170 ;
        RECT 1793.730 735.720 1796.570 736.170 ;
        RECT 1797.410 735.720 1800.250 736.170 ;
        RECT 1801.090 735.720 1803.930 736.170 ;
        RECT 1804.770 735.720 1807.610 736.170 ;
        RECT 1808.450 735.720 1811.290 736.170 ;
        RECT 1812.130 735.720 1814.970 736.170 ;
        RECT 1815.810 735.720 1818.650 736.170 ;
        RECT 1819.490 735.720 1822.330 736.170 ;
        RECT 1823.170 735.720 1826.010 736.170 ;
        RECT 1826.850 735.720 1829.690 736.170 ;
        RECT 1830.530 735.720 1833.370 736.170 ;
        RECT 1834.210 735.720 1837.050 736.170 ;
        RECT 1837.890 735.720 1840.730 736.170 ;
        RECT 1841.570 735.720 1844.410 736.170 ;
        RECT 1845.250 735.720 1848.090 736.170 ;
        RECT 1848.930 735.720 1851.770 736.170 ;
        RECT 1852.610 735.720 1855.450 736.170 ;
        RECT 1856.290 735.720 1859.130 736.170 ;
        RECT 1859.970 735.720 1862.810 736.170 ;
        RECT 1863.650 735.720 1866.490 736.170 ;
        RECT 1867.330 735.720 1870.170 736.170 ;
        RECT 1871.010 735.720 1873.850 736.170 ;
        RECT 1874.690 735.720 1877.530 736.170 ;
        RECT 1878.370 735.720 1881.210 736.170 ;
        RECT 1882.050 735.720 1884.890 736.170 ;
        RECT 1885.730 735.720 1888.570 736.170 ;
        RECT 1889.410 735.720 1892.250 736.170 ;
        RECT 1893.090 735.720 1895.930 736.170 ;
        RECT 1896.770 735.720 1899.610 736.170 ;
        RECT 1900.450 735.720 1903.290 736.170 ;
        RECT 1904.130 735.720 1906.970 736.170 ;
        RECT 1907.810 735.720 1910.650 736.170 ;
        RECT 1911.490 735.720 1914.330 736.170 ;
        RECT 1915.170 735.720 1918.010 736.170 ;
        RECT 1918.850 735.720 1921.690 736.170 ;
        RECT 1922.530 735.720 1925.370 736.170 ;
        RECT 1926.210 735.720 1929.050 736.170 ;
        RECT 1929.890 735.720 1932.730 736.170 ;
        RECT 1933.570 735.720 1936.410 736.170 ;
        RECT 1937.250 735.720 1940.090 736.170 ;
        RECT 1940.930 735.720 1943.770 736.170 ;
        RECT 1944.610 735.720 1947.450 736.170 ;
        RECT 1948.290 735.720 1951.130 736.170 ;
        RECT 1951.970 735.720 1954.810 736.170 ;
        RECT 1955.650 735.720 1958.490 736.170 ;
        RECT 1959.330 735.720 1962.170 736.170 ;
        RECT 1963.010 735.720 1965.850 736.170 ;
        RECT 1966.690 735.720 1969.530 736.170 ;
        RECT 1970.370 735.720 1973.210 736.170 ;
        RECT 1974.050 735.720 1976.890 736.170 ;
        RECT 1977.730 735.720 1980.570 736.170 ;
        RECT 1981.410 735.720 1984.250 736.170 ;
        RECT 1985.090 735.720 1987.930 736.170 ;
        RECT 1988.770 735.720 1991.610 736.170 ;
        RECT 1992.450 735.720 1995.290 736.170 ;
        RECT 1996.130 735.720 1998.970 736.170 ;
        RECT 1999.810 735.720 2002.650 736.170 ;
        RECT 2003.490 735.720 2006.330 736.170 ;
        RECT 2007.170 735.720 2010.010 736.170 ;
        RECT 2010.850 735.720 2013.690 736.170 ;
        RECT 2014.530 735.720 2017.370 736.170 ;
        RECT 2018.210 735.720 2021.050 736.170 ;
        RECT 2021.890 735.720 2024.730 736.170 ;
        RECT 2025.570 735.720 2028.410 736.170 ;
        RECT 2029.250 735.720 2032.090 736.170 ;
        RECT 2032.930 735.720 2035.770 736.170 ;
        RECT 2036.610 735.720 2039.450 736.170 ;
        RECT 2040.290 735.720 2043.130 736.170 ;
        RECT 2043.970 735.720 2046.810 736.170 ;
        RECT 2047.650 735.720 2050.490 736.170 ;
        RECT 2051.330 735.720 2054.170 736.170 ;
        RECT 2055.010 735.720 2057.850 736.170 ;
        RECT 2058.690 735.720 2061.530 736.170 ;
        RECT 2062.370 735.720 2065.210 736.170 ;
        RECT 2066.050 735.720 2068.890 736.170 ;
        RECT 2069.730 735.720 2072.570 736.170 ;
        RECT 2073.410 735.720 2076.250 736.170 ;
        RECT 2077.090 735.720 2079.930 736.170 ;
        RECT 2080.770 735.720 2083.610 736.170 ;
        RECT 2084.450 735.720 2087.290 736.170 ;
        RECT 2088.130 735.720 2090.970 736.170 ;
        RECT 2091.810 735.720 2094.650 736.170 ;
        RECT 2095.490 735.720 2098.330 736.170 ;
        RECT 2099.170 735.720 2102.010 736.170 ;
        RECT 2102.850 735.720 2105.690 736.170 ;
        RECT 2106.530 735.720 2109.370 736.170 ;
        RECT 2110.210 735.720 2113.050 736.170 ;
        RECT 2113.890 735.720 2116.730 736.170 ;
        RECT 2117.570 735.720 2120.410 736.170 ;
        RECT 2121.250 735.720 2124.090 736.170 ;
        RECT 2124.930 735.720 2127.770 736.170 ;
        RECT 2128.610 735.720 2131.450 736.170 ;
        RECT 2132.290 735.720 2135.130 736.170 ;
        RECT 2135.970 735.720 2138.810 736.170 ;
        RECT 2139.650 735.720 2142.490 736.170 ;
        RECT 2143.330 735.720 2146.170 736.170 ;
        RECT 2147.010 735.720 2149.850 736.170 ;
        RECT 2150.690 735.720 2153.530 736.170 ;
        RECT 2154.370 735.720 2157.210 736.170 ;
        RECT 2158.050 735.720 2160.890 736.170 ;
        RECT 2161.730 735.720 2164.570 736.170 ;
        RECT 2165.410 735.720 2168.250 736.170 ;
        RECT 2169.090 735.720 2171.930 736.170 ;
        RECT 2172.770 735.720 2175.610 736.170 ;
        RECT 2176.450 735.720 2179.290 736.170 ;
        RECT 2180.130 735.720 2182.970 736.170 ;
        RECT 2183.810 735.720 2186.650 736.170 ;
        RECT 2187.490 735.720 2190.330 736.170 ;
        RECT 2191.170 735.720 2194.010 736.170 ;
        RECT 2194.850 735.720 2197.690 736.170 ;
        RECT 2198.530 735.720 2201.370 736.170 ;
        RECT 2202.210 735.720 2205.050 736.170 ;
        RECT 2205.890 735.720 2208.730 736.170 ;
        RECT 2209.570 735.720 2212.410 736.170 ;
        RECT 2213.250 735.720 2216.090 736.170 ;
        RECT 2216.930 735.720 2219.770 736.170 ;
        RECT 2220.610 735.720 2223.450 736.170 ;
        RECT 2224.290 735.720 2227.130 736.170 ;
        RECT 2227.970 735.720 2230.810 736.170 ;
        RECT 2231.650 735.720 2234.490 736.170 ;
        RECT 2235.330 735.720 2238.170 736.170 ;
        RECT 2239.010 735.720 2241.850 736.170 ;
        RECT 2242.690 735.720 2245.530 736.170 ;
        RECT 2246.370 735.720 2249.210 736.170 ;
        RECT 2250.050 735.720 2252.890 736.170 ;
        RECT 2253.730 735.720 2256.570 736.170 ;
        RECT 2257.410 735.720 2260.250 736.170 ;
        RECT 2261.090 735.720 2263.930 736.170 ;
        RECT 2264.770 735.720 2267.610 736.170 ;
        RECT 2268.450 735.720 2271.290 736.170 ;
        RECT 2272.130 735.720 2274.970 736.170 ;
        RECT 2275.810 735.720 2278.650 736.170 ;
        RECT 2279.490 735.720 2282.330 736.170 ;
        RECT 2283.170 735.720 2286.010 736.170 ;
        RECT 2286.850 735.720 2289.690 736.170 ;
        RECT 2290.530 735.720 2293.370 736.170 ;
        RECT 2294.210 735.720 2297.050 736.170 ;
        RECT 2297.890 735.720 2300.730 736.170 ;
        RECT 2301.570 735.720 2304.410 736.170 ;
        RECT 2305.250 735.720 2308.090 736.170 ;
        RECT 2308.930 735.720 2311.770 736.170 ;
        RECT 2312.610 735.720 2315.450 736.170 ;
        RECT 2316.290 735.720 2319.130 736.170 ;
        RECT 2319.970 735.720 2322.810 736.170 ;
        RECT 2323.650 735.720 2326.490 736.170 ;
        RECT 2327.330 735.720 2330.170 736.170 ;
        RECT 2331.010 735.720 2333.850 736.170 ;
        RECT 2334.690 735.720 2337.530 736.170 ;
        RECT 2338.370 735.720 2341.210 736.170 ;
        RECT 2342.050 735.720 2344.890 736.170 ;
        RECT 2345.730 735.720 2348.570 736.170 ;
        RECT 2349.410 735.720 2352.250 736.170 ;
        RECT 2353.090 735.720 2355.930 736.170 ;
        RECT 2356.770 735.720 2359.610 736.170 ;
        RECT 2360.450 735.720 2363.290 736.170 ;
        RECT 2364.130 735.720 2366.970 736.170 ;
        RECT 2367.810 735.720 2370.650 736.170 ;
        RECT 2371.490 735.720 2374.330 736.170 ;
        RECT 2375.170 735.720 2378.010 736.170 ;
        RECT 2378.850 735.720 2381.690 736.170 ;
        RECT 2382.530 735.720 2385.370 736.170 ;
        RECT 2386.210 735.720 2389.050 736.170 ;
        RECT 2389.890 735.720 2392.730 736.170 ;
        RECT 2393.570 735.720 2396.410 736.170 ;
        RECT 2397.250 735.720 2400.090 736.170 ;
        RECT 2400.930 735.720 2403.770 736.170 ;
        RECT 2404.610 735.720 2519.780 736.170 ;
        RECT 6.070 4.280 2519.780 735.720 ;
        RECT 6.070 1.030 1384.870 4.280 ;
        RECT 1385.710 1.030 1468.590 4.280 ;
        RECT 1469.430 1.030 1887.190 4.280 ;
        RECT 1888.030 1.030 1970.910 4.280 ;
        RECT 1971.750 1.030 2054.630 4.280 ;
        RECT 2055.470 1.030 2138.350 4.280 ;
        RECT 2139.190 1.030 2222.070 4.280 ;
        RECT 2222.910 1.030 2305.790 4.280 ;
        RECT 2306.630 1.030 2519.780 4.280 ;
      LAYER met3 ;
        RECT 3.990 728.640 2519.355 731.505 ;
        RECT 3.990 727.240 2515.600 728.640 ;
        RECT 3.990 717.760 2519.355 727.240 ;
        RECT 3.990 716.360 2515.600 717.760 ;
        RECT 3.990 706.880 2519.355 716.360 ;
        RECT 3.990 705.480 2515.600 706.880 ;
        RECT 3.990 696.000 2519.355 705.480 ;
        RECT 3.990 694.600 2515.600 696.000 ;
        RECT 3.990 685.120 2519.355 694.600 ;
        RECT 3.990 683.720 2515.600 685.120 ;
        RECT 3.990 675.600 2519.355 683.720 ;
        RECT 4.400 674.240 2519.355 675.600 ;
        RECT 4.400 674.200 2515.600 674.240 ;
        RECT 3.990 672.840 2515.600 674.200 ;
        RECT 3.990 663.360 2519.355 672.840 ;
        RECT 3.990 661.960 2515.600 663.360 ;
        RECT 3.990 652.480 2519.355 661.960 ;
        RECT 3.990 651.080 2515.600 652.480 ;
        RECT 3.990 641.600 2519.355 651.080 ;
        RECT 3.990 640.200 2515.600 641.600 ;
        RECT 3.990 630.720 2519.355 640.200 ;
        RECT 3.990 629.320 2515.600 630.720 ;
        RECT 3.990 619.840 2519.355 629.320 ;
        RECT 3.990 618.440 2515.600 619.840 ;
        RECT 3.990 608.960 2519.355 618.440 ;
        RECT 3.990 607.560 2515.600 608.960 ;
        RECT 3.990 598.080 2519.355 607.560 ;
        RECT 3.990 596.680 2515.600 598.080 ;
        RECT 3.990 587.200 2519.355 596.680 ;
        RECT 3.990 585.800 2515.600 587.200 ;
        RECT 3.990 576.320 2519.355 585.800 ;
        RECT 3.990 574.920 2515.600 576.320 ;
        RECT 3.990 565.440 2519.355 574.920 ;
        RECT 3.990 564.040 2515.600 565.440 ;
        RECT 3.990 554.560 2519.355 564.040 ;
        RECT 3.990 553.200 2515.600 554.560 ;
        RECT 4.400 553.160 2515.600 553.200 ;
        RECT 4.400 551.800 2519.355 553.160 ;
        RECT 3.990 543.680 2519.355 551.800 ;
        RECT 3.990 542.280 2515.600 543.680 ;
        RECT 3.990 532.800 2519.355 542.280 ;
        RECT 3.990 531.400 2515.600 532.800 ;
        RECT 3.990 521.920 2519.355 531.400 ;
        RECT 3.990 520.520 2515.600 521.920 ;
        RECT 3.990 511.040 2519.355 520.520 ;
        RECT 3.990 509.640 2515.600 511.040 ;
        RECT 3.990 500.160 2519.355 509.640 ;
        RECT 3.990 498.760 2515.600 500.160 ;
        RECT 3.990 489.280 2519.355 498.760 ;
        RECT 3.990 487.880 2515.600 489.280 ;
        RECT 3.990 478.400 2519.355 487.880 ;
        RECT 3.990 477.000 2515.600 478.400 ;
        RECT 3.990 467.520 2519.355 477.000 ;
        RECT 3.990 466.120 2515.600 467.520 ;
        RECT 3.990 456.640 2519.355 466.120 ;
        RECT 3.990 455.240 2515.600 456.640 ;
        RECT 3.990 445.760 2519.355 455.240 ;
        RECT 3.990 444.360 2515.600 445.760 ;
        RECT 3.990 434.880 2519.355 444.360 ;
        RECT 3.990 433.480 2515.600 434.880 ;
        RECT 3.990 430.800 2519.355 433.480 ;
        RECT 4.400 429.400 2519.355 430.800 ;
        RECT 3.990 424.000 2519.355 429.400 ;
        RECT 3.990 422.600 2515.600 424.000 ;
        RECT 3.990 413.120 2519.355 422.600 ;
        RECT 3.990 411.720 2515.600 413.120 ;
        RECT 3.990 402.240 2519.355 411.720 ;
        RECT 3.990 400.840 2515.600 402.240 ;
        RECT 3.990 391.360 2519.355 400.840 ;
        RECT 3.990 389.960 2515.600 391.360 ;
        RECT 3.990 380.480 2519.355 389.960 ;
        RECT 3.990 379.080 2515.600 380.480 ;
        RECT 3.990 369.600 2519.355 379.080 ;
        RECT 3.990 368.200 2515.600 369.600 ;
        RECT 3.990 358.720 2519.355 368.200 ;
        RECT 3.990 357.320 2515.600 358.720 ;
        RECT 3.990 347.840 2519.355 357.320 ;
        RECT 3.990 346.440 2515.600 347.840 ;
        RECT 3.990 336.960 2519.355 346.440 ;
        RECT 3.990 335.560 2515.600 336.960 ;
        RECT 3.990 326.080 2519.355 335.560 ;
        RECT 3.990 324.680 2515.600 326.080 ;
        RECT 3.990 315.200 2519.355 324.680 ;
        RECT 3.990 313.800 2515.600 315.200 ;
        RECT 3.990 308.400 2519.355 313.800 ;
        RECT 4.400 307.000 2519.355 308.400 ;
        RECT 3.990 304.320 2519.355 307.000 ;
        RECT 3.990 302.920 2515.600 304.320 ;
        RECT 3.990 293.440 2519.355 302.920 ;
        RECT 3.990 292.040 2515.600 293.440 ;
        RECT 3.990 282.560 2519.355 292.040 ;
        RECT 3.990 281.160 2515.600 282.560 ;
        RECT 3.990 271.680 2519.355 281.160 ;
        RECT 3.990 270.280 2515.600 271.680 ;
        RECT 3.990 260.800 2519.355 270.280 ;
        RECT 3.990 259.400 2515.600 260.800 ;
        RECT 3.990 249.920 2519.355 259.400 ;
        RECT 3.990 248.520 2515.600 249.920 ;
        RECT 3.990 239.040 2519.355 248.520 ;
        RECT 3.990 237.640 2515.600 239.040 ;
        RECT 3.990 228.160 2519.355 237.640 ;
        RECT 3.990 226.760 2515.600 228.160 ;
        RECT 3.990 217.280 2519.355 226.760 ;
        RECT 3.990 215.880 2515.600 217.280 ;
        RECT 3.990 206.400 2519.355 215.880 ;
        RECT 3.990 205.000 2515.600 206.400 ;
        RECT 3.990 195.520 2519.355 205.000 ;
        RECT 3.990 194.120 2515.600 195.520 ;
        RECT 3.990 186.000 2519.355 194.120 ;
        RECT 4.400 184.640 2519.355 186.000 ;
        RECT 4.400 184.600 2515.600 184.640 ;
        RECT 3.990 183.240 2515.600 184.600 ;
        RECT 3.990 173.760 2519.355 183.240 ;
        RECT 3.990 172.360 2515.600 173.760 ;
        RECT 3.990 162.880 2519.355 172.360 ;
        RECT 3.990 161.480 2515.600 162.880 ;
        RECT 3.990 152.000 2519.355 161.480 ;
        RECT 3.990 150.600 2515.600 152.000 ;
        RECT 3.990 141.120 2519.355 150.600 ;
        RECT 3.990 139.720 2515.600 141.120 ;
        RECT 3.990 130.240 2519.355 139.720 ;
        RECT 3.990 128.840 2515.600 130.240 ;
        RECT 3.990 119.360 2519.355 128.840 ;
        RECT 3.990 117.960 2515.600 119.360 ;
        RECT 3.990 108.480 2519.355 117.960 ;
        RECT 3.990 107.080 2515.600 108.480 ;
        RECT 3.990 97.600 2519.355 107.080 ;
        RECT 3.990 96.200 2515.600 97.600 ;
        RECT 3.990 86.720 2519.355 96.200 ;
        RECT 3.990 85.320 2515.600 86.720 ;
        RECT 3.990 75.840 2519.355 85.320 ;
        RECT 3.990 74.440 2515.600 75.840 ;
        RECT 3.990 64.960 2519.355 74.440 ;
        RECT 3.990 63.600 2515.600 64.960 ;
        RECT 4.400 63.560 2515.600 63.600 ;
        RECT 4.400 62.200 2519.355 63.560 ;
        RECT 3.990 54.080 2519.355 62.200 ;
        RECT 3.990 52.680 2515.600 54.080 ;
        RECT 3.990 43.200 2519.355 52.680 ;
        RECT 3.990 41.800 2515.600 43.200 ;
        RECT 3.990 32.320 2519.355 41.800 ;
        RECT 3.990 30.920 2515.600 32.320 ;
        RECT 3.990 21.440 2519.355 30.920 ;
        RECT 3.990 20.040 2515.600 21.440 ;
        RECT 3.990 10.560 2519.355 20.040 ;
        RECT 3.990 9.160 2515.600 10.560 ;
        RECT 3.990 5.615 2519.355 9.160 ;
      LAYER met4 ;
        RECT 16.855 5.615 20.640 724.705 ;
        RECT 23.040 5.615 32.240 724.705 ;
        RECT 34.640 585.110 70.640 724.705 ;
        RECT 73.040 585.110 82.240 724.705 ;
        RECT 34.640 52.870 82.240 585.110 ;
        RECT 34.640 5.615 70.640 52.870 ;
        RECT 73.040 5.615 82.240 52.870 ;
        RECT 84.640 5.615 120.640 724.705 ;
        RECT 123.040 585.110 132.240 724.705 ;
        RECT 134.640 585.110 170.640 724.705 ;
        RECT 123.040 52.870 170.640 585.110 ;
        RECT 123.040 5.615 132.240 52.870 ;
        RECT 134.640 5.615 170.640 52.870 ;
        RECT 173.040 5.615 182.240 724.705 ;
        RECT 184.640 585.110 220.640 724.705 ;
        RECT 223.040 585.110 232.240 724.705 ;
        RECT 184.640 554.475 232.240 585.110 ;
        RECT 234.640 554.475 270.640 724.705 ;
        RECT 273.040 585.110 282.240 724.705 ;
        RECT 284.640 585.110 320.640 724.705 ;
        RECT 273.040 554.475 320.640 585.110 ;
        RECT 323.040 554.475 332.240 724.705 ;
        RECT 334.640 585.110 370.640 724.705 ;
        RECT 373.040 585.110 382.240 724.705 ;
        RECT 334.640 554.475 382.240 585.110 ;
        RECT 384.640 554.475 420.640 724.705 ;
        RECT 423.040 585.110 432.240 724.705 ;
        RECT 434.640 585.110 470.640 724.705 ;
        RECT 423.040 554.475 470.640 585.110 ;
        RECT 473.040 554.475 482.240 724.705 ;
        RECT 484.640 585.110 520.640 724.705 ;
        RECT 523.040 585.110 532.240 724.705 ;
        RECT 484.640 554.475 532.240 585.110 ;
        RECT 534.640 554.475 570.640 724.705 ;
        RECT 573.040 585.110 582.240 724.705 ;
        RECT 584.640 585.110 620.640 724.705 ;
        RECT 573.040 554.475 620.640 585.110 ;
        RECT 623.040 554.475 632.240 724.705 ;
        RECT 634.640 585.110 670.640 724.705 ;
        RECT 673.040 585.110 682.240 724.705 ;
        RECT 634.640 554.475 682.240 585.110 ;
        RECT 684.640 554.475 720.640 724.705 ;
        RECT 723.040 585.110 732.240 724.705 ;
        RECT 734.640 585.110 770.640 724.705 ;
        RECT 723.040 554.475 770.640 585.110 ;
        RECT 773.040 554.475 782.240 724.705 ;
        RECT 784.640 585.110 820.640 724.705 ;
        RECT 823.040 585.110 832.240 724.705 ;
        RECT 784.640 554.475 832.240 585.110 ;
        RECT 834.640 554.475 870.640 724.705 ;
        RECT 873.040 585.110 882.240 724.705 ;
        RECT 884.640 585.110 920.640 724.705 ;
        RECT 873.040 554.475 920.640 585.110 ;
        RECT 923.040 554.475 932.240 724.705 ;
        RECT 934.640 585.110 970.640 724.705 ;
        RECT 973.040 585.110 982.240 724.705 ;
        RECT 934.640 554.475 982.240 585.110 ;
        RECT 984.640 554.475 1020.640 724.705 ;
        RECT 1023.040 585.110 1032.240 724.705 ;
        RECT 1034.640 585.110 1070.640 724.705 ;
        RECT 1023.040 554.475 1070.640 585.110 ;
        RECT 1073.040 554.475 1082.240 724.705 ;
        RECT 1084.640 585.110 1120.640 724.705 ;
        RECT 1123.040 585.110 1132.240 724.705 ;
        RECT 1084.640 554.475 1132.240 585.110 ;
        RECT 1134.640 554.475 1170.640 724.705 ;
        RECT 1173.040 585.110 1182.240 724.705 ;
        RECT 1184.640 585.110 1220.640 724.705 ;
        RECT 1173.040 554.475 1220.640 585.110 ;
        RECT 184.640 104.585 1220.640 554.475 ;
        RECT 184.640 52.870 232.240 104.585 ;
        RECT 184.640 5.615 220.640 52.870 ;
        RECT 223.040 5.615 232.240 52.870 ;
        RECT 234.640 5.615 270.640 104.585 ;
        RECT 273.040 52.870 320.640 104.585 ;
        RECT 273.040 5.615 282.240 52.870 ;
        RECT 284.640 5.615 320.640 52.870 ;
        RECT 323.040 5.615 332.240 104.585 ;
        RECT 334.640 52.870 382.240 104.585 ;
        RECT 334.640 5.615 370.640 52.870 ;
        RECT 373.040 5.615 382.240 52.870 ;
        RECT 384.640 5.615 420.640 104.585 ;
        RECT 423.040 52.870 470.640 104.585 ;
        RECT 423.040 5.615 432.240 52.870 ;
        RECT 434.640 5.615 470.640 52.870 ;
        RECT 473.040 5.615 482.240 104.585 ;
        RECT 484.640 52.870 532.240 104.585 ;
        RECT 484.640 5.615 520.640 52.870 ;
        RECT 523.040 5.615 532.240 52.870 ;
        RECT 534.640 5.615 570.640 104.585 ;
        RECT 573.040 52.870 620.640 104.585 ;
        RECT 573.040 5.615 582.240 52.870 ;
        RECT 584.640 5.615 620.640 52.870 ;
        RECT 623.040 5.615 632.240 104.585 ;
        RECT 634.640 52.870 682.240 104.585 ;
        RECT 634.640 5.615 670.640 52.870 ;
        RECT 673.040 5.615 682.240 52.870 ;
        RECT 684.640 5.615 720.640 104.585 ;
        RECT 723.040 52.870 770.640 104.585 ;
        RECT 723.040 5.615 732.240 52.870 ;
        RECT 734.640 5.615 770.640 52.870 ;
        RECT 773.040 5.615 782.240 104.585 ;
        RECT 784.640 52.870 832.240 104.585 ;
        RECT 784.640 5.615 820.640 52.870 ;
        RECT 823.040 5.615 832.240 52.870 ;
        RECT 834.640 5.615 870.640 104.585 ;
        RECT 873.040 52.870 920.640 104.585 ;
        RECT 873.040 5.615 882.240 52.870 ;
        RECT 884.640 5.615 920.640 52.870 ;
        RECT 923.040 5.615 932.240 104.585 ;
        RECT 934.640 52.870 982.240 104.585 ;
        RECT 934.640 5.615 970.640 52.870 ;
        RECT 973.040 5.615 982.240 52.870 ;
        RECT 984.640 5.615 1020.640 104.585 ;
        RECT 1023.040 52.870 1070.640 104.585 ;
        RECT 1023.040 5.615 1032.240 52.870 ;
        RECT 1034.640 5.615 1070.640 52.870 ;
        RECT 1073.040 5.615 1082.240 104.585 ;
        RECT 1084.640 52.870 1132.240 104.585 ;
        RECT 1084.640 5.615 1120.640 52.870 ;
        RECT 1123.040 5.615 1132.240 52.870 ;
        RECT 1134.640 5.615 1170.640 104.585 ;
        RECT 1173.040 52.870 1220.640 104.585 ;
        RECT 1173.040 5.615 1182.240 52.870 ;
        RECT 1184.640 5.615 1220.640 52.870 ;
        RECT 1223.040 5.615 1232.240 724.705 ;
        RECT 1234.640 5.615 1270.640 724.705 ;
        RECT 1273.040 5.615 1282.240 724.705 ;
        RECT 1284.640 5.615 1320.640 724.705 ;
        RECT 1323.040 5.615 1332.240 724.705 ;
        RECT 1334.640 5.615 1370.640 724.705 ;
        RECT 1373.040 5.615 1382.240 724.705 ;
        RECT 1384.640 5.615 1420.640 724.705 ;
        RECT 1423.040 5.615 1432.240 724.705 ;
        RECT 1434.640 5.615 1470.640 724.705 ;
        RECT 1473.040 5.615 1482.240 724.705 ;
        RECT 1484.640 5.615 1520.640 724.705 ;
        RECT 1523.040 5.615 1532.240 724.705 ;
        RECT 1534.640 5.615 1570.640 724.705 ;
        RECT 1573.040 5.615 1582.240 724.705 ;
        RECT 1584.640 5.615 1620.640 724.705 ;
        RECT 1623.040 5.615 1632.240 724.705 ;
        RECT 1634.640 5.615 1670.640 724.705 ;
        RECT 1673.040 5.615 1682.240 724.705 ;
        RECT 1684.640 5.615 1720.640 724.705 ;
        RECT 1723.040 5.615 1732.240 724.705 ;
        RECT 1734.640 5.615 1770.640 724.705 ;
        RECT 1773.040 5.615 1782.240 724.705 ;
        RECT 1784.640 5.615 1820.640 724.705 ;
        RECT 1823.040 5.615 1832.240 724.705 ;
        RECT 1834.640 5.615 1870.640 724.705 ;
        RECT 1873.040 5.615 1882.240 724.705 ;
        RECT 1884.640 5.615 1920.640 724.705 ;
        RECT 1923.040 5.615 1932.240 724.705 ;
        RECT 1934.640 5.615 1970.640 724.705 ;
        RECT 1973.040 5.615 1982.240 724.705 ;
        RECT 1984.640 580.760 2020.640 724.705 ;
        RECT 2023.040 580.760 2032.240 724.705 ;
        RECT 2034.640 580.760 2070.640 724.705 ;
        RECT 2073.040 580.760 2082.240 724.705 ;
        RECT 2084.640 580.760 2120.640 724.705 ;
        RECT 2123.040 580.760 2132.240 724.705 ;
        RECT 2134.640 580.760 2170.640 724.705 ;
        RECT 2173.040 580.760 2182.240 724.705 ;
        RECT 2184.640 580.760 2220.640 724.705 ;
        RECT 2223.040 580.760 2232.240 724.705 ;
        RECT 2234.640 580.760 2270.640 724.705 ;
        RECT 2273.040 580.760 2282.240 724.705 ;
        RECT 2284.640 580.760 2320.640 724.705 ;
        RECT 2323.040 580.760 2332.240 724.705 ;
        RECT 2334.640 580.760 2370.640 724.705 ;
        RECT 2373.040 580.760 2382.240 724.705 ;
        RECT 2384.640 580.760 2420.640 724.705 ;
        RECT 2423.040 580.760 2432.240 724.705 ;
        RECT 2434.640 580.760 2470.640 724.705 ;
        RECT 1984.640 70.350 2470.640 580.760 ;
        RECT 1984.640 5.615 2020.640 70.350 ;
        RECT 2023.040 5.615 2032.240 70.350 ;
        RECT 2034.640 5.615 2070.640 70.350 ;
        RECT 2073.040 5.615 2082.240 70.350 ;
        RECT 2084.640 5.615 2120.640 70.350 ;
        RECT 2123.040 5.615 2132.240 70.350 ;
        RECT 2134.640 5.615 2170.640 70.350 ;
        RECT 2173.040 5.615 2182.240 70.350 ;
        RECT 2184.640 5.615 2220.640 70.350 ;
        RECT 2223.040 5.615 2232.240 70.350 ;
        RECT 2234.640 5.615 2270.640 70.350 ;
        RECT 2273.040 5.615 2282.240 70.350 ;
        RECT 2284.640 5.615 2320.640 70.350 ;
        RECT 2323.040 5.615 2332.240 70.350 ;
        RECT 2334.640 5.615 2370.640 70.350 ;
        RECT 2373.040 5.615 2382.240 70.350 ;
        RECT 2384.640 5.615 2420.640 70.350 ;
        RECT 2423.040 5.615 2432.240 70.350 ;
        RECT 2434.640 5.615 2470.640 70.350 ;
        RECT 2473.040 5.615 2482.240 724.705 ;
        RECT 2484.640 626.240 2514.490 724.705 ;
        RECT 2484.640 34.720 2493.380 626.240 ;
        RECT 2495.780 34.720 2505.340 626.240 ;
        RECT 2507.740 34.720 2514.490 626.240 ;
        RECT 2484.640 5.615 2514.490 34.720 ;
      LAYER met5 ;
        RECT 473.460 691.530 2514.700 702.900 ;
        RECT 473.460 679.930 2514.700 686.730 ;
        RECT 473.460 641.530 2514.700 675.130 ;
        RECT 473.460 629.930 2514.700 636.730 ;
        RECT 473.460 591.530 2514.700 625.130 ;
        RECT 473.460 579.930 2514.700 586.730 ;
        RECT 473.460 541.530 2514.700 575.130 ;
        RECT 473.460 529.930 2514.700 536.730 ;
        RECT 473.460 491.530 2514.700 525.130 ;
        RECT 473.460 479.930 2514.700 486.730 ;
        RECT 473.460 441.530 2514.700 475.130 ;
        RECT 473.460 429.930 2514.700 436.730 ;
        RECT 473.460 391.530 2514.700 425.130 ;
        RECT 473.460 379.930 2514.700 386.730 ;
        RECT 473.460 341.530 2514.700 375.130 ;
        RECT 473.460 329.930 2514.700 336.730 ;
        RECT 473.460 291.530 2514.700 325.130 ;
        RECT 473.460 279.930 2514.700 286.730 ;
        RECT 473.460 241.530 2514.700 275.130 ;
        RECT 473.460 229.930 2514.700 236.730 ;
        RECT 473.460 191.530 2514.700 225.130 ;
        RECT 473.460 179.930 2514.700 186.730 ;
        RECT 473.460 141.530 2514.700 175.130 ;
        RECT 473.460 129.930 2514.700 136.730 ;
        RECT 473.460 91.530 2514.700 125.130 ;
        RECT 473.460 79.930 2514.700 86.730 ;
        RECT 473.460 41.530 2514.700 75.130 ;
        RECT 473.460 31.500 2514.700 36.730 ;
  END
END mgmt_core_wrapper
END LIBRARY

