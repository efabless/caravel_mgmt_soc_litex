magic
tech sky130A
magscale 1 2
timestamp 1637325823
<< obsli1 >>
rect 1869 2159 107916 145809
<< obsm1 >>
rect 1670 1980 108270 146192
<< metal2 >>
rect 1674 147200 1730 148000
rect 5078 147200 5134 148000
rect 8482 147200 8538 148000
rect 11978 147200 12034 148000
rect 15382 147200 15438 148000
rect 18786 147200 18842 148000
rect 22282 147200 22338 148000
rect 25686 147200 25742 148000
rect 29182 147200 29238 148000
rect 32586 147200 32642 148000
rect 35990 147200 36046 148000
rect 39486 147200 39542 148000
rect 42890 147200 42946 148000
rect 46294 147200 46350 148000
rect 49790 147200 49846 148000
rect 53194 147200 53250 148000
rect 56690 147200 56746 148000
rect 60094 147200 60150 148000
rect 63498 147200 63554 148000
rect 66994 147200 67050 148000
rect 70398 147200 70454 148000
rect 73802 147200 73858 148000
rect 77298 147200 77354 148000
rect 80702 147200 80758 148000
rect 84198 147200 84254 148000
rect 87602 147200 87658 148000
rect 91006 147200 91062 148000
rect 94502 147200 94558 148000
rect 97906 147200 97962 148000
rect 101310 147200 101366 148000
rect 104806 147200 104862 148000
rect 108210 147200 108266 148000
rect 1674 0 1730 800
rect 4986 0 5042 800
rect 8298 0 8354 800
rect 11610 0 11666 800
rect 14922 0 14978 800
rect 18326 0 18382 800
rect 21638 0 21694 800
rect 24950 0 25006 800
rect 28262 0 28318 800
rect 31666 0 31722 800
rect 34978 0 35034 800
rect 38290 0 38346 800
rect 41602 0 41658 800
rect 45006 0 45062 800
rect 48318 0 48374 800
rect 51630 0 51686 800
rect 54942 0 54998 800
rect 58346 0 58402 800
rect 61658 0 61714 800
rect 64970 0 65026 800
rect 68282 0 68338 800
rect 71686 0 71742 800
rect 74998 0 75054 800
rect 78310 0 78366 800
rect 81622 0 81678 800
rect 85026 0 85082 800
rect 88338 0 88394 800
rect 91650 0 91706 800
rect 94962 0 95018 800
rect 98366 0 98422 800
rect 101678 0 101734 800
rect 104990 0 105046 800
rect 108302 0 108358 800
<< obsm2 >>
rect 1786 147144 5022 147234
rect 5190 147144 8426 147234
rect 8594 147144 11922 147234
rect 12090 147144 15326 147234
rect 15494 147144 18730 147234
rect 18898 147144 22226 147234
rect 22394 147144 25630 147234
rect 25798 147144 29126 147234
rect 29294 147144 32530 147234
rect 32698 147144 35934 147234
rect 36102 147144 39430 147234
rect 39598 147144 42834 147234
rect 43002 147144 46238 147234
rect 46406 147144 49734 147234
rect 49902 147144 53138 147234
rect 53306 147144 56634 147234
rect 56802 147144 60038 147234
rect 60206 147144 63442 147234
rect 63610 147144 66938 147234
rect 67106 147144 70342 147234
rect 70510 147144 73746 147234
rect 73914 147144 77242 147234
rect 77410 147144 80646 147234
rect 80814 147144 84142 147234
rect 84310 147144 87546 147234
rect 87714 147144 90950 147234
rect 91118 147144 94446 147234
rect 94614 147144 97850 147234
rect 98018 147144 101254 147234
rect 101422 147144 104750 147234
rect 104918 147144 108154 147234
rect 108322 147144 108344 147234
rect 1674 856 108344 147144
rect 1786 734 4930 856
rect 5098 734 8242 856
rect 8410 734 11554 856
rect 11722 734 14866 856
rect 15034 734 18270 856
rect 18438 734 21582 856
rect 21750 734 24894 856
rect 25062 734 28206 856
rect 28374 734 31610 856
rect 31778 734 34922 856
rect 35090 734 38234 856
rect 38402 734 41546 856
rect 41714 734 44950 856
rect 45118 734 48262 856
rect 48430 734 51574 856
rect 51742 734 54886 856
rect 55054 734 58290 856
rect 58458 734 61602 856
rect 61770 734 64914 856
rect 65082 734 68226 856
rect 68394 734 71630 856
rect 71798 734 74942 856
rect 75110 734 78254 856
rect 78422 734 81566 856
rect 81734 734 84970 856
rect 85138 734 88282 856
rect 88450 734 91594 856
rect 91762 734 94906 856
rect 95074 734 98310 856
rect 98478 734 101622 856
rect 101790 734 104934 856
rect 105102 734 108246 856
<< metal3 >>
rect 109200 142128 110000 142248
rect 109200 130704 110000 130824
rect 109200 119280 110000 119400
rect 109200 107992 110000 108112
rect 109200 96568 110000 96688
rect 109200 85144 110000 85264
rect 109200 73856 110000 73976
rect 109200 62432 110000 62552
rect 109200 51008 110000 51128
rect 109200 39720 110000 39840
rect 109200 28296 110000 28416
rect 109200 16872 110000 16992
rect 109200 5584 110000 5704
<< obsm3 >>
rect 1669 142328 109200 145825
rect 1669 142048 109120 142328
rect 1669 130904 109200 142048
rect 1669 130624 109120 130904
rect 1669 119480 109200 130624
rect 1669 119200 109120 119480
rect 1669 108192 109200 119200
rect 1669 107912 109120 108192
rect 1669 96768 109200 107912
rect 1669 96488 109120 96768
rect 1669 85344 109200 96488
rect 1669 85064 109120 85344
rect 1669 74056 109200 85064
rect 1669 73776 109120 74056
rect 1669 62632 109200 73776
rect 1669 62352 109120 62632
rect 1669 51208 109200 62352
rect 1669 50928 109120 51208
rect 1669 39920 109200 50928
rect 1669 39640 109120 39920
rect 1669 28496 109200 39640
rect 1669 28216 109120 28496
rect 1669 17072 109200 28216
rect 1669 16792 109120 17072
rect 1669 5784 109200 16792
rect 1669 5504 109120 5784
rect 1669 2143 109200 5504
<< metal4 >>
rect 4 156 324 147812
rect 664 816 984 147152
rect 5128 156 5448 147812
rect 20488 156 20808 147812
rect 35848 156 36168 147812
rect 51208 156 51528 147812
rect 66568 156 66888 147812
rect 81928 156 82248 147812
rect 97288 156 97608 147812
rect 108956 816 109276 147152
rect 109616 156 109936 147812
<< obsm4 >>
rect 4475 2891 5048 145485
rect 5528 2891 20408 145485
rect 20888 2891 35768 145485
rect 36248 2891 51128 145485
rect 51608 2891 66488 145485
rect 66968 2891 81848 145485
rect 82328 2891 97208 145485
rect 97688 2891 100037 145485
<< metal5 >>
rect 4 147492 109936 147812
rect 664 146832 109276 147152
rect 4 135298 109936 135618
rect 4 122298 109936 122618
rect 4 109298 109936 109618
rect 4 96298 109936 96618
rect 4 83298 109936 83618
rect 4 70298 109936 70618
rect 4 57298 109936 57618
rect 4 44298 109936 44618
rect 4 31298 109936 31618
rect 4 18298 109936 18618
rect 4 5298 109936 5618
rect 664 816 109276 1136
rect 4 156 109936 476
<< labels >>
rlabel metal3 s 109200 5584 110000 5704 6 A[0]
port 1 nsew signal input
rlabel metal3 s 109200 16872 110000 16992 6 A[1]
port 2 nsew signal input
rlabel metal3 s 109200 28296 110000 28416 6 A[2]
port 3 nsew signal input
rlabel metal3 s 109200 39720 110000 39840 6 A[3]
port 4 nsew signal input
rlabel metal3 s 109200 51008 110000 51128 6 A[4]
port 5 nsew signal input
rlabel metal3 s 109200 62432 110000 62552 6 A[5]
port 6 nsew signal input
rlabel metal3 s 109200 73856 110000 73976 6 A[6]
port 7 nsew signal input
rlabel metal3 s 109200 85144 110000 85264 6 A[7]
port 8 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 CLK
port 9 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 Di[0]
port 10 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 Di[10]
port 11 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 Di[11]
port 12 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 Di[12]
port 13 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 Di[13]
port 14 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 Di[14]
port 15 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 Di[15]
port 16 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 Di[16]
port 17 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 Di[17]
port 18 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 Di[18]
port 19 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 Di[19]
port 20 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 Di[1]
port 21 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 Di[20]
port 22 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 Di[21]
port 23 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 Di[22]
port 24 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 Di[23]
port 25 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 Di[24]
port 26 nsew signal input
rlabel metal2 s 88338 0 88394 800 6 Di[25]
port 27 nsew signal input
rlabel metal2 s 91650 0 91706 800 6 Di[26]
port 28 nsew signal input
rlabel metal2 s 94962 0 95018 800 6 Di[27]
port 29 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 Di[28]
port 30 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 Di[29]
port 31 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 Di[2]
port 32 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 Di[30]
port 33 nsew signal input
rlabel metal2 s 108302 0 108358 800 6 Di[31]
port 34 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 Di[3]
port 35 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 Di[4]
port 36 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 Di[5]
port 37 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 Di[6]
port 38 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 Di[7]
port 39 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 Di[8]
port 40 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 Di[9]
port 41 nsew signal input
rlabel metal2 s 1674 147200 1730 148000 6 Do[0]
port 42 nsew signal output
rlabel metal2 s 35990 147200 36046 148000 6 Do[10]
port 43 nsew signal output
rlabel metal2 s 39486 147200 39542 148000 6 Do[11]
port 44 nsew signal output
rlabel metal2 s 42890 147200 42946 148000 6 Do[12]
port 45 nsew signal output
rlabel metal2 s 46294 147200 46350 148000 6 Do[13]
port 46 nsew signal output
rlabel metal2 s 49790 147200 49846 148000 6 Do[14]
port 47 nsew signal output
rlabel metal2 s 53194 147200 53250 148000 6 Do[15]
port 48 nsew signal output
rlabel metal2 s 56690 147200 56746 148000 6 Do[16]
port 49 nsew signal output
rlabel metal2 s 60094 147200 60150 148000 6 Do[17]
port 50 nsew signal output
rlabel metal2 s 63498 147200 63554 148000 6 Do[18]
port 51 nsew signal output
rlabel metal2 s 66994 147200 67050 148000 6 Do[19]
port 52 nsew signal output
rlabel metal2 s 5078 147200 5134 148000 6 Do[1]
port 53 nsew signal output
rlabel metal2 s 70398 147200 70454 148000 6 Do[20]
port 54 nsew signal output
rlabel metal2 s 73802 147200 73858 148000 6 Do[21]
port 55 nsew signal output
rlabel metal2 s 77298 147200 77354 148000 6 Do[22]
port 56 nsew signal output
rlabel metal2 s 80702 147200 80758 148000 6 Do[23]
port 57 nsew signal output
rlabel metal2 s 84198 147200 84254 148000 6 Do[24]
port 58 nsew signal output
rlabel metal2 s 87602 147200 87658 148000 6 Do[25]
port 59 nsew signal output
rlabel metal2 s 91006 147200 91062 148000 6 Do[26]
port 60 nsew signal output
rlabel metal2 s 94502 147200 94558 148000 6 Do[27]
port 61 nsew signal output
rlabel metal2 s 97906 147200 97962 148000 6 Do[28]
port 62 nsew signal output
rlabel metal2 s 101310 147200 101366 148000 6 Do[29]
port 63 nsew signal output
rlabel metal2 s 8482 147200 8538 148000 6 Do[2]
port 64 nsew signal output
rlabel metal2 s 104806 147200 104862 148000 6 Do[30]
port 65 nsew signal output
rlabel metal2 s 108210 147200 108266 148000 6 Do[31]
port 66 nsew signal output
rlabel metal2 s 11978 147200 12034 148000 6 Do[3]
port 67 nsew signal output
rlabel metal2 s 15382 147200 15438 148000 6 Do[4]
port 68 nsew signal output
rlabel metal2 s 18786 147200 18842 148000 6 Do[5]
port 69 nsew signal output
rlabel metal2 s 22282 147200 22338 148000 6 Do[6]
port 70 nsew signal output
rlabel metal2 s 25686 147200 25742 148000 6 Do[7]
port 71 nsew signal output
rlabel metal2 s 29182 147200 29238 148000 6 Do[8]
port 72 nsew signal output
rlabel metal2 s 32586 147200 32642 148000 6 Do[9]
port 73 nsew signal output
rlabel metal3 s 109200 142128 110000 142248 6 EN
port 74 nsew signal input
rlabel metal5 s 4 156 109936 476 6 VGND
port 75 nsew ground input
rlabel metal5 s 4 18298 109936 18618 6 VGND
port 75 nsew ground input
rlabel metal5 s 4 44298 109936 44618 6 VGND
port 75 nsew ground input
rlabel metal5 s 4 70298 109936 70618 6 VGND
port 75 nsew ground input
rlabel metal5 s 4 96298 109936 96618 6 VGND
port 75 nsew ground input
rlabel metal5 s 4 122298 109936 122618 6 VGND
port 75 nsew ground input
rlabel metal5 s 4 147492 109936 147812 6 VGND
port 75 nsew ground input
rlabel metal4 s 4 156 324 147812 6 VGND
port 75 nsew ground input
rlabel metal4 s 20488 156 20808 147812 6 VGND
port 75 nsew ground input
rlabel metal4 s 51208 156 51528 147812 6 VGND
port 75 nsew ground input
rlabel metal4 s 81928 156 82248 147812 6 VGND
port 75 nsew ground input
rlabel metal4 s 109616 156 109936 147812 6 VGND
port 75 nsew ground input
rlabel metal5 s 664 816 109276 1136 6 VPWR
port 76 nsew power input
rlabel metal5 s 4 5298 109936 5618 6 VPWR
port 76 nsew power input
rlabel metal5 s 4 31298 109936 31618 6 VPWR
port 76 nsew power input
rlabel metal5 s 4 57298 109936 57618 6 VPWR
port 76 nsew power input
rlabel metal5 s 4 83298 109936 83618 6 VPWR
port 76 nsew power input
rlabel metal5 s 4 109298 109936 109618 6 VPWR
port 76 nsew power input
rlabel metal5 s 4 135298 109936 135618 6 VPWR
port 76 nsew power input
rlabel metal5 s 664 146832 109276 147152 6 VPWR
port 76 nsew power input
rlabel metal4 s 664 816 984 147152 6 VPWR
port 76 nsew power input
rlabel metal4 s 108956 816 109276 147152 6 VPWR
port 76 nsew power input
rlabel metal4 s 5128 156 5448 147812 6 VPWR
port 76 nsew power input
rlabel metal4 s 35848 156 36168 147812 6 VPWR
port 76 nsew power input
rlabel metal4 s 66568 156 66888 147812 6 VPWR
port 76 nsew power input
rlabel metal4 s 97288 156 97608 147812 6 VPWR
port 76 nsew power input
rlabel metal3 s 109200 96568 110000 96688 6 WE[0]
port 77 nsew signal input
rlabel metal3 s 109200 107992 110000 108112 6 WE[1]
port 78 nsew signal input
rlabel metal3 s 109200 119280 110000 119400 6 WE[2]
port 79 nsew signal input
rlabel metal3 s 109200 130704 110000 130824 6 WE[3]
port 80 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 110000 148000
string LEFview TRUE
string GDS_FILE ../gds/DFFRAM.gds
string GDS_END 59531056
string GDS_START 181858
<< end >>

