magic
tech sky130A
magscale 1 2
timestamp 1648060287
<< metal1 >>
rect 168558 160284 168564 160336
rect 168616 160324 168622 160336
rect 173342 160324 173348 160336
rect 168616 160296 173348 160324
rect 168616 160284 168622 160296
rect 173342 160284 173348 160296
rect 173400 160284 173406 160336
rect 63402 160012 63408 160064
rect 63460 160052 63466 160064
rect 146478 160052 146484 160064
rect 63460 160024 146484 160052
rect 63460 160012 63466 160024
rect 146478 160012 146484 160024
rect 146536 160012 146542 160064
rect 146938 160012 146944 160064
rect 146996 160052 147002 160064
rect 154482 160052 154488 160064
rect 146996 160024 154488 160052
rect 146996 160012 147002 160024
rect 154482 160012 154488 160024
rect 154540 160012 154546 160064
rect 156782 160012 156788 160064
rect 156840 160052 156846 160064
rect 191650 160052 191656 160064
rect 156840 160024 191656 160052
rect 156840 160012 156846 160024
rect 191650 160012 191656 160024
rect 191708 160012 191714 160064
rect 197170 160012 197176 160064
rect 197228 160052 197234 160064
rect 207014 160052 207020 160064
rect 197228 160024 207020 160052
rect 197228 160012 197234 160024
rect 207014 160012 207020 160024
rect 207072 160012 207078 160064
rect 211430 160012 211436 160064
rect 211488 160052 211494 160064
rect 280338 160052 280344 160064
rect 211488 160024 280344 160052
rect 211488 160012 211494 160024
rect 280338 160012 280344 160024
rect 280396 160012 280402 160064
rect 281258 160012 281264 160064
rect 281316 160052 281322 160064
rect 332686 160052 332692 160064
rect 281316 160024 332692 160052
rect 281316 160012 281322 160024
rect 332686 160012 332692 160024
rect 332744 160012 332750 160064
rect 334250 160012 334256 160064
rect 334308 160052 334314 160064
rect 374086 160052 374092 160064
rect 334308 160024 374092 160052
rect 334308 160012 334314 160024
rect 374086 160012 374092 160024
rect 374144 160012 374150 160064
rect 378870 160012 378876 160064
rect 378928 160052 378934 160064
rect 391382 160052 391388 160064
rect 378928 160024 391388 160052
rect 378928 160012 378934 160024
rect 391382 160012 391388 160024
rect 391440 160012 391446 160064
rect 391474 160012 391480 160064
rect 391532 160052 391538 160064
rect 394602 160052 394608 160064
rect 391532 160024 394608 160052
rect 391532 160012 391538 160024
rect 394602 160012 394608 160024
rect 394660 160012 394666 160064
rect 400766 160012 400772 160064
rect 400824 160052 400830 160064
rect 424870 160052 424876 160064
rect 400824 160024 424876 160052
rect 400824 160012 400830 160024
rect 424870 160012 424876 160024
rect 424928 160012 424934 160064
rect 25590 159944 25596 159996
rect 25648 159984 25654 159996
rect 110322 159984 110328 159996
rect 25648 159956 110328 159984
rect 25648 159944 25654 159956
rect 110322 159944 110328 159956
rect 110380 159944 110386 159996
rect 117222 159944 117228 159996
rect 117280 159984 117286 159996
rect 191466 159984 191472 159996
rect 117280 159956 191472 159984
rect 117280 159944 117286 159956
rect 191466 159944 191472 159956
rect 191524 159944 191530 159996
rect 197998 159944 198004 159996
rect 198056 159984 198062 159996
rect 269114 159984 269120 159996
rect 198056 159956 269120 159984
rect 198056 159944 198062 159956
rect 269114 159944 269120 159956
rect 269172 159944 269178 159996
rect 271230 159944 271236 159996
rect 271288 159984 271294 159996
rect 272794 159984 272800 159996
rect 271288 159956 272800 159984
rect 271288 159944 271294 159956
rect 272794 159944 272800 159956
rect 272852 159944 272858 159996
rect 275370 159944 275376 159996
rect 275428 159984 275434 159996
rect 328454 159984 328460 159996
rect 275428 159956 328460 159984
rect 275428 159944 275434 159956
rect 328454 159944 328460 159956
rect 328512 159944 328518 159996
rect 329190 159944 329196 159996
rect 329248 159984 329254 159996
rect 369946 159984 369952 159996
rect 329248 159956 369952 159984
rect 329248 159944 329254 159956
rect 369946 159944 369952 159956
rect 370004 159944 370010 159996
rect 372154 159944 372160 159996
rect 372212 159984 372218 159996
rect 396166 159984 396172 159996
rect 372212 159956 396172 159984
rect 372212 159944 372218 159956
rect 396166 159944 396172 159956
rect 396224 159944 396230 159996
rect 403250 159944 403256 159996
rect 403308 159984 403314 159996
rect 415854 159984 415860 159996
rect 403308 159956 415860 159984
rect 403308 159944 403314 159956
rect 415854 159944 415860 159956
rect 415912 159944 415918 159996
rect 76926 159876 76932 159928
rect 76984 159916 76990 159928
rect 162486 159916 162492 159928
rect 76984 159888 162492 159916
rect 76984 159876 76990 159888
rect 162486 159876 162492 159888
rect 162544 159876 162550 159928
rect 166902 159876 166908 159928
rect 166960 159916 166966 159928
rect 186406 159916 186412 159928
rect 166960 159888 186412 159916
rect 166960 159876 166966 159888
rect 186406 159876 186412 159888
rect 186464 159876 186470 159928
rect 191282 159876 191288 159928
rect 191340 159916 191346 159928
rect 264882 159916 264888 159928
rect 191340 159888 264888 159916
rect 191340 159876 191346 159888
rect 264882 159876 264888 159888
rect 264940 159876 264946 159928
rect 268654 159876 268660 159928
rect 268712 159916 268718 159928
rect 324038 159916 324044 159928
rect 268712 159888 324044 159916
rect 268712 159876 268718 159888
rect 324038 159876 324044 159888
rect 324096 159876 324102 159928
rect 328362 159876 328368 159928
rect 328420 159916 328426 159928
rect 369486 159916 369492 159928
rect 328420 159888 369492 159916
rect 328420 159876 328426 159888
rect 369486 159876 369492 159888
rect 369544 159876 369550 159928
rect 379698 159876 379704 159928
rect 379756 159916 379762 159928
rect 405826 159916 405832 159928
rect 379756 159888 405832 159916
rect 379756 159876 379762 159888
rect 405826 159876 405832 159888
rect 405884 159876 405890 159928
rect 457070 159876 457076 159928
rect 457128 159916 457134 159928
rect 464338 159916 464344 159928
rect 457128 159888 464344 159916
rect 457128 159876 457134 159888
rect 464338 159876 464344 159888
rect 464396 159876 464402 159928
rect 480622 159876 480628 159928
rect 480680 159916 480686 159928
rect 485958 159916 485964 159928
rect 480680 159888 485964 159916
rect 480680 159876 480686 159888
rect 485958 159876 485964 159888
rect 486016 159876 486022 159928
rect 70118 159808 70124 159860
rect 70176 159848 70182 159860
rect 156322 159848 156328 159860
rect 70176 159820 156328 159848
rect 70176 159808 70182 159820
rect 156322 159808 156328 159820
rect 156380 159808 156386 159860
rect 160094 159848 160100 159860
rect 156708 159820 160100 159848
rect 56686 159740 56692 159792
rect 56744 159780 56750 159792
rect 137278 159780 137284 159792
rect 56744 159752 137284 159780
rect 56744 159740 56750 159752
rect 137278 159740 137284 159752
rect 137336 159740 137342 159792
rect 137370 159740 137376 159792
rect 137428 159780 137434 159792
rect 139394 159780 139400 159792
rect 137428 159752 139400 159780
rect 137428 159740 137434 159752
rect 139394 159740 139400 159752
rect 139452 159740 139458 159792
rect 139946 159740 139952 159792
rect 140004 159780 140010 159792
rect 147030 159780 147036 159792
rect 140004 159752 147036 159780
rect 140004 159740 140010 159752
rect 147030 159740 147036 159752
rect 147088 159740 147094 159792
rect 147122 159740 147128 159792
rect 147180 159780 147186 159792
rect 148318 159780 148324 159792
rect 147180 159752 148324 159780
rect 147180 159740 147186 159752
rect 148318 159740 148324 159752
rect 148376 159740 148382 159792
rect 153470 159740 153476 159792
rect 153528 159780 153534 159792
rect 156598 159780 156604 159792
rect 153528 159752 156604 159780
rect 153528 159740 153534 159752
rect 156598 159740 156604 159752
rect 156656 159740 156662 159792
rect 18874 159672 18880 159724
rect 18932 159712 18938 159724
rect 109218 159712 109224 159724
rect 18932 159684 109224 159712
rect 18932 159672 18938 159684
rect 109218 159672 109224 159684
rect 109276 159672 109282 159724
rect 113082 159672 113088 159724
rect 113140 159712 113146 159724
rect 126422 159712 126428 159724
rect 113140 159684 126428 159712
rect 113140 159672 113146 159684
rect 126422 159672 126428 159684
rect 126480 159672 126486 159724
rect 126514 159672 126520 159724
rect 126572 159712 126578 159724
rect 156506 159712 156512 159724
rect 126572 159684 156512 159712
rect 126572 159672 126578 159684
rect 156506 159672 156512 159684
rect 156564 159672 156570 159724
rect 156708 159712 156736 159820
rect 160094 159808 160100 159820
rect 160152 159808 160158 159860
rect 179414 159848 179420 159860
rect 161446 159820 179420 159848
rect 156782 159740 156788 159792
rect 156840 159780 156846 159792
rect 161446 159780 161474 159820
rect 179414 159808 179420 159820
rect 179472 159808 179478 159860
rect 184566 159808 184572 159860
rect 184624 159848 184630 159860
rect 259546 159848 259552 159860
rect 184624 159820 259552 159848
rect 184624 159808 184630 159820
rect 259546 159808 259552 159820
rect 259604 159808 259610 159860
rect 261110 159808 261116 159860
rect 261168 159848 261174 159860
rect 317046 159848 317052 159860
rect 261168 159820 317052 159848
rect 261168 159808 261174 159820
rect 317046 159808 317052 159820
rect 317104 159808 317110 159860
rect 320818 159808 320824 159860
rect 320876 159848 320882 159860
rect 362954 159848 362960 159860
rect 320876 159820 362960 159848
rect 320876 159808 320882 159820
rect 362954 159808 362960 159820
rect 363012 159808 363018 159860
rect 376294 159808 376300 159860
rect 376352 159848 376358 159860
rect 406194 159848 406200 159860
rect 376352 159820 406200 159848
rect 376352 159808 376358 159820
rect 406194 159808 406200 159820
rect 406252 159808 406258 159860
rect 409966 159808 409972 159860
rect 410024 159848 410030 159860
rect 417234 159848 417240 159860
rect 410024 159820 417240 159848
rect 410024 159808 410030 159820
rect 417234 159808 417240 159820
rect 417292 159808 417298 159860
rect 446122 159808 446128 159860
rect 446180 159848 446186 159860
rect 456794 159848 456800 159860
rect 446180 159820 456800 159848
rect 446180 159808 446186 159820
rect 456794 159808 456800 159820
rect 456852 159808 456858 159860
rect 458726 159808 458732 159860
rect 458784 159848 458790 159860
rect 465074 159848 465080 159860
rect 458784 159820 465080 159848
rect 458784 159808 458790 159820
rect 465074 159808 465080 159820
rect 465132 159808 465138 159860
rect 472250 159808 472256 159860
rect 472308 159848 472314 159860
rect 479426 159848 479432 159860
rect 472308 159820 479432 159848
rect 472308 159808 472314 159820
rect 479426 159808 479432 159820
rect 479484 159808 479490 159860
rect 156840 159752 161474 159780
rect 156840 159740 156846 159752
rect 171134 159740 171140 159792
rect 171192 159780 171198 159792
rect 173250 159780 173256 159792
rect 171192 159752 173256 159780
rect 171192 159740 171198 159752
rect 173250 159740 173256 159752
rect 173308 159740 173314 159792
rect 177850 159740 177856 159792
rect 177908 159780 177914 159792
rect 253934 159780 253940 159792
rect 177908 159752 253940 159780
rect 177908 159740 177914 159752
rect 253934 159740 253940 159752
rect 253992 159740 253998 159792
rect 261938 159740 261944 159792
rect 261996 159780 262002 159792
rect 318886 159780 318892 159792
rect 261996 159752 318892 159780
rect 261996 159740 262002 159752
rect 318886 159740 318892 159752
rect 318944 159740 318950 159792
rect 322474 159740 322480 159792
rect 322532 159780 322538 159792
rect 365162 159780 365168 159792
rect 322532 159752 365168 159780
rect 322532 159740 322538 159752
rect 365162 159740 365168 159752
rect 365220 159740 365226 159792
rect 365438 159740 365444 159792
rect 365496 159780 365502 159792
rect 395522 159780 395528 159792
rect 365496 159752 395528 159780
rect 365496 159740 365502 159752
rect 395522 159740 395528 159752
rect 395580 159740 395586 159792
rect 396534 159740 396540 159792
rect 396592 159780 396598 159792
rect 413186 159780 413192 159792
rect 396592 159752 413192 159780
rect 396592 159740 396598 159752
rect 413186 159740 413192 159752
rect 413244 159740 413250 159792
rect 413370 159740 413376 159792
rect 413428 159780 413434 159792
rect 419626 159780 419632 159792
rect 413428 159752 419632 159780
rect 413428 159740 413434 159752
rect 419626 159740 419632 159752
rect 419684 159740 419690 159792
rect 420914 159740 420920 159792
rect 420972 159780 420978 159792
rect 440418 159780 440424 159792
rect 420972 159752 440424 159780
rect 420972 159740 420978 159752
rect 440418 159740 440424 159752
rect 440476 159740 440482 159792
rect 448698 159740 448704 159792
rect 448756 159780 448762 159792
rect 460934 159780 460940 159792
rect 448756 159752 460940 159780
rect 448756 159740 448762 159752
rect 460934 159740 460940 159752
rect 460992 159740 460998 159792
rect 469674 159740 469680 159792
rect 469732 159780 469738 159792
rect 477402 159780 477408 159792
rect 469732 159752 477408 159780
rect 469732 159740 469738 159752
rect 477402 159740 477408 159752
rect 477460 159740 477466 159792
rect 478966 159740 478972 159792
rect 479024 159780 479030 159792
rect 484670 159780 484676 159792
rect 479024 159752 484676 159780
rect 479024 159740 479030 159752
rect 484670 159740 484676 159752
rect 484728 159740 484734 159792
rect 163774 159712 163780 159724
rect 156616 159684 156736 159712
rect 156800 159684 163780 159712
rect 49970 159604 49976 159656
rect 50028 159644 50034 159656
rect 143258 159644 143264 159656
rect 50028 159616 143264 159644
rect 50028 159604 50034 159616
rect 143258 159604 143264 159616
rect 143316 159604 143322 159656
rect 143350 159604 143356 159656
rect 143408 159644 143414 159656
rect 156616 159644 156644 159684
rect 143408 159616 156644 159644
rect 143408 159604 143414 159616
rect 43254 159536 43260 159588
rect 43312 159576 43318 159588
rect 136818 159576 136824 159588
rect 43312 159548 136824 159576
rect 43312 159536 43318 159548
rect 136818 159536 136824 159548
rect 136876 159536 136882 159588
rect 137278 159536 137284 159588
rect 137336 159576 137342 159588
rect 143994 159576 144000 159588
rect 137336 159548 144000 159576
rect 137336 159536 137342 159548
rect 143994 159536 144000 159548
rect 144052 159536 144058 159588
rect 144086 159536 144092 159588
rect 144144 159576 144150 159588
rect 146846 159576 146852 159588
rect 144144 159548 146852 159576
rect 144144 159536 144150 159548
rect 146846 159536 146852 159548
rect 146904 159536 146910 159588
rect 147214 159536 147220 159588
rect 147272 159576 147278 159588
rect 156800 159576 156828 159684
rect 163774 159672 163780 159684
rect 163832 159672 163838 159724
rect 167730 159672 167736 159724
rect 167788 159712 167794 159724
rect 246942 159712 246948 159724
rect 167788 159684 246948 159712
rect 167788 159672 167794 159684
rect 246942 159672 246948 159684
rect 247000 159672 247006 159724
rect 255222 159672 255228 159724
rect 255280 159712 255286 159724
rect 313366 159712 313372 159724
rect 255280 159684 313372 159712
rect 255280 159672 255286 159684
rect 313366 159672 313372 159684
rect 313424 159672 313430 159724
rect 314102 159672 314108 159724
rect 314160 159712 314166 159724
rect 357986 159712 357992 159724
rect 314160 159684 357992 159712
rect 314160 159672 314166 159684
rect 357986 159672 357992 159684
rect 358044 159672 358050 159724
rect 369578 159672 369584 159724
rect 369636 159712 369642 159724
rect 401042 159712 401048 159724
rect 369636 159684 401048 159712
rect 369636 159672 369642 159684
rect 401042 159672 401048 159684
rect 401100 159672 401106 159724
rect 407482 159672 407488 159724
rect 407540 159712 407546 159724
rect 429930 159712 429936 159724
rect 407540 159684 429936 159712
rect 407540 159672 407546 159684
rect 429930 159672 429936 159684
rect 429988 159672 429994 159724
rect 451182 159672 451188 159724
rect 451240 159712 451246 159724
rect 462314 159712 462320 159724
rect 451240 159684 462320 159712
rect 451240 159672 451246 159684
rect 462314 159672 462320 159684
rect 462372 159672 462378 159724
rect 468018 159672 468024 159724
rect 468076 159712 468082 159724
rect 476022 159712 476028 159724
rect 468076 159684 476028 159712
rect 468076 159672 468082 159684
rect 476022 159672 476028 159684
rect 476080 159672 476086 159724
rect 479794 159672 479800 159724
rect 479852 159712 479858 159724
rect 485222 159712 485228 159724
rect 479852 159684 485228 159712
rect 479852 159672 479858 159684
rect 485222 159672 485228 159684
rect 485280 159672 485286 159724
rect 161014 159604 161020 159656
rect 161072 159644 161078 159656
rect 240318 159644 240324 159656
rect 161072 159616 240324 159644
rect 161072 159604 161078 159616
rect 240318 159604 240324 159616
rect 240376 159604 240382 159656
rect 241790 159604 241796 159656
rect 241848 159644 241854 159656
rect 302234 159644 302240 159656
rect 241848 159616 302240 159644
rect 241848 159604 241854 159616
rect 302234 159604 302240 159616
rect 302292 159604 302298 159656
rect 302326 159604 302332 159656
rect 302384 159644 302390 159656
rect 349246 159644 349252 159656
rect 302384 159616 349252 159644
rect 302384 159604 302390 159616
rect 349246 159604 349252 159616
rect 349304 159604 349310 159656
rect 351914 159604 351920 159656
rect 351972 159644 351978 159656
rect 385770 159644 385776 159656
rect 351972 159616 385776 159644
rect 351972 159604 351978 159616
rect 385770 159604 385776 159616
rect 385828 159604 385834 159656
rect 388070 159604 388076 159656
rect 388128 159644 388134 159656
rect 389082 159644 389088 159656
rect 388128 159616 389088 159644
rect 388128 159604 388134 159616
rect 389082 159604 389088 159616
rect 389140 159604 389146 159656
rect 389818 159604 389824 159656
rect 389876 159644 389882 159656
rect 413370 159644 413376 159656
rect 389876 159616 413376 159644
rect 389876 159604 389882 159616
rect 413370 159604 413376 159616
rect 413428 159604 413434 159656
rect 417510 159604 417516 159656
rect 417568 159644 417574 159656
rect 437658 159644 437664 159656
rect 417568 159616 437664 159644
rect 417568 159604 417574 159616
rect 437658 159604 437664 159616
rect 437716 159604 437722 159656
rect 453758 159604 453764 159656
rect 453816 159644 453822 159656
rect 465258 159644 465264 159656
rect 453816 159616 465264 159644
rect 453816 159604 453822 159616
rect 465258 159604 465264 159616
rect 465316 159604 465322 159656
rect 147272 159548 156828 159576
rect 147272 159536 147278 159548
rect 157610 159536 157616 159588
rect 157668 159576 157674 159588
rect 239306 159576 239312 159588
rect 157668 159548 239312 159576
rect 157668 159536 157674 159548
rect 239306 159536 239312 159548
rect 239364 159536 239370 159588
rect 250990 159536 250996 159588
rect 251048 159576 251054 159588
rect 310606 159576 310612 159588
rect 251048 159548 310612 159576
rect 251048 159536 251054 159548
rect 310606 159536 310612 159548
rect 310664 159536 310670 159588
rect 315758 159536 315764 159588
rect 315816 159576 315822 159588
rect 358906 159576 358912 159588
rect 315816 159548 358912 159576
rect 315816 159536 315822 159548
rect 358906 159536 358912 159548
rect 358964 159536 358970 159588
rect 362862 159536 362868 159588
rect 362920 159576 362926 159588
rect 394970 159576 394976 159588
rect 362920 159548 394976 159576
rect 362920 159536 362926 159548
rect 394970 159536 394976 159548
rect 395028 159536 395034 159588
rect 399018 159536 399024 159588
rect 399076 159576 399082 159588
rect 408494 159576 408500 159588
rect 399076 159548 408500 159576
rect 399076 159536 399082 159548
rect 408494 159536 408500 159548
rect 408552 159536 408558 159588
rect 410794 159536 410800 159588
rect 410852 159576 410858 159588
rect 432506 159576 432512 159588
rect 410852 159548 432512 159576
rect 410852 159536 410858 159548
rect 432506 159536 432512 159548
rect 432564 159536 432570 159588
rect 452010 159536 452016 159588
rect 452068 159576 452074 159588
rect 463970 159576 463976 159588
rect 452068 159548 463976 159576
rect 452068 159536 452074 159548
rect 463970 159536 463976 159548
rect 464028 159536 464034 159588
rect 467190 159536 467196 159588
rect 467248 159576 467254 159588
rect 473354 159576 473360 159588
rect 467248 159548 473360 159576
rect 467248 159536 467254 159548
rect 473354 159536 473360 159548
rect 473412 159536 473418 159588
rect 36538 159468 36544 159520
rect 36596 159508 36602 159520
rect 126330 159508 126336 159520
rect 36596 159480 126336 159508
rect 36596 159468 36602 159480
rect 126330 159468 126336 159480
rect 126388 159468 126394 159520
rect 126422 159468 126428 159520
rect 126480 159508 126486 159520
rect 127618 159508 127624 159520
rect 126480 159480 127624 159508
rect 126480 159468 126486 159480
rect 127618 159468 127624 159480
rect 127676 159468 127682 159520
rect 129918 159468 129924 159520
rect 129976 159508 129982 159520
rect 146938 159508 146944 159520
rect 129976 159480 146944 159508
rect 129976 159468 129982 159480
rect 146938 159468 146944 159480
rect 146996 159468 147002 159520
rect 225322 159508 225328 159520
rect 147508 159480 225328 159508
rect 32306 159400 32312 159452
rect 32364 159440 32370 159452
rect 126606 159440 126612 159452
rect 32364 159412 126612 159440
rect 32364 159400 32370 159412
rect 126606 159400 126612 159412
rect 126664 159400 126670 159452
rect 130746 159400 130752 159452
rect 130804 159440 130810 159452
rect 137186 159440 137192 159452
rect 130804 159412 137192 159440
rect 130804 159400 130810 159412
rect 137186 159400 137192 159412
rect 137244 159400 137250 159452
rect 144086 159440 144092 159452
rect 137296 159412 144092 159440
rect 6270 159332 6276 159384
rect 6328 159372 6334 159384
rect 122834 159372 122840 159384
rect 6328 159344 122840 159372
rect 6328 159332 6334 159344
rect 122834 159332 122840 159344
rect 122892 159332 122898 159384
rect 123110 159332 123116 159384
rect 123168 159372 123174 159384
rect 137296 159372 137324 159412
rect 144086 159400 144092 159412
rect 144144 159400 144150 159452
rect 144178 159400 144184 159452
rect 144236 159440 144242 159452
rect 147508 159440 147536 159480
rect 225322 159468 225328 159480
rect 225380 159468 225386 159520
rect 231670 159468 231676 159520
rect 231728 159508 231734 159520
rect 295518 159508 295524 159520
rect 231728 159480 295524 159508
rect 231728 159468 231734 159480
rect 295518 159468 295524 159480
rect 295576 159468 295582 159520
rect 295610 159468 295616 159520
rect 295668 159508 295674 159520
rect 342438 159508 342444 159520
rect 295668 159480 342444 159508
rect 295668 159468 295674 159480
rect 342438 159468 342444 159480
rect 342496 159468 342502 159520
rect 347682 159468 347688 159520
rect 347740 159508 347746 159520
rect 354214 159508 354220 159520
rect 347740 159480 354220 159508
rect 347740 159468 347746 159480
rect 354214 159468 354220 159480
rect 354272 159468 354278 159520
rect 356146 159468 356152 159520
rect 356204 159508 356210 159520
rect 390554 159508 390560 159520
rect 356204 159480 390560 159508
rect 356204 159468 356210 159480
rect 390554 159468 390560 159480
rect 390612 159468 390618 159520
rect 391382 159468 391388 159520
rect 391440 159508 391446 159520
rect 398558 159508 398564 159520
rect 391440 159480 398564 159508
rect 391440 159468 391446 159480
rect 398558 159468 398564 159480
rect 398616 159468 398622 159520
rect 424318 159468 424324 159520
rect 424376 159508 424382 159520
rect 442810 159508 442816 159520
rect 424376 159480 442816 159508
rect 424376 159468 424382 159480
rect 442810 159468 442816 159480
rect 442868 159468 442874 159520
rect 447870 159468 447876 159520
rect 447928 159508 447934 159520
rect 460106 159508 460112 159520
rect 447928 159480 460112 159508
rect 447928 159468 447934 159480
rect 460106 159468 460112 159480
rect 460164 159468 460170 159520
rect 461302 159468 461308 159520
rect 461360 159508 461366 159520
rect 467926 159508 467932 159520
rect 461360 159480 467932 159508
rect 461360 159468 461366 159480
rect 467926 159468 467932 159480
rect 467984 159468 467990 159520
rect 481450 159468 481456 159520
rect 481508 159508 481514 159520
rect 486510 159508 486516 159520
rect 481508 159480 486516 159508
rect 481508 159468 481514 159480
rect 486510 159468 486516 159480
rect 486568 159468 486574 159520
rect 518802 159468 518808 159520
rect 518860 159508 518866 159520
rect 522666 159508 522672 159520
rect 518860 159480 522672 159508
rect 518860 159468 518866 159480
rect 522666 159468 522672 159480
rect 522724 159468 522730 159520
rect 144236 159412 147536 159440
rect 144236 159400 144242 159412
rect 147582 159400 147588 159452
rect 147640 159440 147646 159452
rect 149514 159440 149520 159452
rect 147640 159412 149520 159440
rect 147640 159400 147646 159412
rect 149514 159400 149520 159412
rect 149572 159400 149578 159452
rect 150894 159400 150900 159452
rect 150952 159440 150958 159452
rect 233234 159440 233240 159452
rect 150952 159412 233240 159440
rect 150952 159400 150958 159412
rect 233234 159400 233240 159412
rect 233292 159400 233298 159452
rect 234982 159400 234988 159452
rect 235040 159440 235046 159452
rect 298002 159440 298008 159452
rect 235040 159412 298008 159440
rect 235040 159400 235046 159412
rect 298002 159400 298008 159412
rect 298060 159400 298066 159452
rect 301498 159400 301504 159452
rect 301556 159440 301562 159452
rect 349062 159440 349068 159452
rect 301556 159412 349068 159440
rect 301556 159400 301562 159412
rect 349062 159400 349068 159412
rect 349120 159400 349126 159452
rect 349798 159400 349804 159452
rect 349856 159440 349862 159452
rect 354858 159440 354864 159452
rect 349856 159412 354864 159440
rect 349856 159400 349862 159412
rect 354858 159400 354864 159412
rect 354916 159400 354922 159452
rect 358630 159400 358636 159452
rect 358688 159440 358694 159452
rect 392762 159440 392768 159452
rect 358688 159412 392768 159440
rect 358688 159400 358694 159412
rect 392762 159400 392768 159412
rect 392820 159400 392826 159452
rect 404078 159400 404084 159452
rect 404136 159440 404142 159452
rect 427354 159440 427360 159452
rect 404136 159412 427360 159440
rect 404136 159400 404142 159412
rect 427354 159400 427360 159412
rect 427412 159400 427418 159452
rect 427630 159400 427636 159452
rect 427688 159440 427694 159452
rect 445386 159440 445392 159452
rect 427688 159412 445392 159440
rect 427688 159400 427694 159412
rect 445386 159400 445392 159412
rect 445444 159400 445450 159452
rect 449526 159400 449532 159452
rect 449584 159440 449590 159452
rect 461486 159440 461492 159452
rect 449584 159412 461492 159440
rect 449584 159400 449590 159412
rect 461486 159400 461492 159412
rect 461544 159400 461550 159452
rect 468846 159400 468852 159452
rect 468904 159440 468910 159452
rect 474826 159440 474832 159452
rect 468904 159412 474832 159440
rect 468904 159400 468910 159412
rect 474826 159400 474832 159412
rect 474884 159400 474890 159452
rect 477310 159400 477316 159452
rect 477368 159440 477374 159452
rect 483290 159440 483296 159452
rect 477368 159412 483296 159440
rect 477368 159400 477374 159412
rect 483290 159400 483296 159412
rect 483348 159400 483354 159452
rect 123168 159344 137324 159372
rect 123168 159332 123174 159344
rect 137462 159332 137468 159384
rect 137520 159372 137526 159384
rect 223574 159372 223580 159384
rect 137520 159344 223580 159372
rect 137520 159332 137526 159344
rect 223574 159332 223580 159344
rect 223632 159332 223638 159384
rect 224954 159332 224960 159384
rect 225012 159372 225018 159384
rect 290642 159372 290648 159384
rect 225012 159344 290648 159372
rect 225012 159332 225018 159344
rect 290642 159332 290648 159344
rect 290700 159332 290706 159384
rect 294782 159332 294788 159384
rect 294840 159372 294846 159384
rect 342254 159372 342260 159384
rect 294840 159344 342260 159372
rect 294840 159332 294846 159344
rect 342254 159332 342260 159344
rect 342312 159332 342318 159384
rect 342714 159332 342720 159384
rect 342772 159372 342778 159384
rect 343634 159372 343640 159384
rect 342772 159344 343640 159372
rect 342772 159332 342778 159344
rect 343634 159332 343640 159344
rect 343692 159332 343698 159384
rect 346026 159332 346032 159384
rect 346084 159372 346090 159384
rect 382826 159372 382832 159384
rect 346084 159344 382832 159372
rect 346084 159332 346090 159344
rect 382826 159332 382832 159344
rect 382884 159332 382890 159384
rect 414198 159332 414204 159384
rect 414256 159372 414262 159384
rect 435082 159372 435088 159384
rect 414256 159344 435088 159372
rect 414256 159332 414262 159344
rect 435082 159332 435088 159344
rect 435140 159332 435146 159384
rect 450354 159332 450360 159384
rect 450412 159372 450418 159384
rect 462682 159372 462688 159384
rect 450412 159344 462688 159372
rect 450412 159332 450418 159344
rect 462682 159332 462688 159344
rect 462740 159332 462746 159384
rect 470502 159332 470508 159384
rect 470560 159372 470566 159384
rect 476114 159372 476120 159384
rect 470560 159344 476120 159372
rect 470560 159332 470566 159344
rect 476114 159332 476120 159344
rect 476172 159332 476178 159384
rect 478138 159332 478144 159384
rect 478196 159372 478202 159384
rect 483198 159372 483204 159384
rect 478196 159344 483204 159372
rect 478196 159332 478202 159344
rect 483198 159332 483204 159344
rect 483256 159332 483262 159384
rect 518710 159332 518716 159384
rect 518768 159372 518774 159384
rect 523494 159372 523500 159384
rect 518768 159344 523500 159372
rect 518768 159332 518774 159344
rect 523494 159332 523500 159344
rect 523552 159332 523558 159384
rect 73522 159264 73528 159316
rect 73580 159304 73586 159316
rect 80054 159304 80060 159316
rect 73580 159276 80060 159304
rect 73580 159264 73586 159276
rect 80054 159264 80060 159276
rect 80112 159264 80118 159316
rect 83642 159264 83648 159316
rect 83700 159304 83706 159316
rect 166994 159304 167000 159316
rect 83700 159276 167000 159304
rect 83700 159264 83706 159276
rect 166994 159264 167000 159276
rect 167052 159264 167058 159316
rect 170214 159264 170220 159316
rect 170272 159304 170278 159316
rect 198918 159304 198924 159316
rect 170272 159276 198924 159304
rect 170272 159264 170278 159276
rect 198918 159264 198924 159276
rect 198976 159264 198982 159316
rect 201402 159264 201408 159316
rect 201460 159304 201466 159316
rect 213730 159304 213736 159316
rect 201460 159276 213736 159304
rect 201460 159264 201466 159276
rect 213730 159264 213736 159276
rect 213788 159264 213794 159316
rect 214006 159264 214012 159316
rect 214064 159304 214070 159316
rect 281534 159304 281540 159316
rect 214064 159276 281540 159304
rect 214064 159264 214070 159276
rect 281534 159264 281540 159276
rect 281592 159264 281598 159316
rect 282086 159264 282092 159316
rect 282144 159304 282150 159316
rect 334342 159304 334348 159316
rect 282144 159276 334348 159304
rect 282144 159264 282150 159276
rect 334342 159264 334348 159276
rect 334400 159264 334406 159316
rect 335078 159264 335084 159316
rect 335136 159304 335142 159316
rect 374730 159304 374736 159316
rect 335136 159276 374736 159304
rect 335136 159264 335142 159276
rect 374730 159264 374736 159276
rect 374788 159264 374794 159316
rect 378042 159264 378048 159316
rect 378100 159304 378106 159316
rect 388346 159304 388352 159316
rect 378100 159276 388352 159304
rect 378100 159264 378106 159276
rect 388346 159264 388352 159276
rect 388404 159264 388410 159316
rect 388990 159264 388996 159316
rect 389048 159304 389054 159316
rect 395154 159304 395160 159316
rect 389048 159276 395160 159304
rect 389048 159264 389054 159276
rect 395154 159264 395160 159276
rect 395212 159264 395218 159316
rect 462130 159264 462136 159316
rect 462188 159304 462194 159316
rect 467834 159304 467840 159316
rect 462188 159276 467840 159304
rect 462188 159264 462194 159276
rect 467834 159264 467840 159276
rect 467892 159264 467898 159316
rect 80238 159196 80244 159248
rect 80296 159236 80302 159248
rect 91094 159236 91100 159248
rect 80296 159208 91100 159236
rect 80296 159196 80302 159208
rect 91094 159196 91100 159208
rect 91152 159196 91158 159248
rect 100478 159196 100484 159248
rect 100536 159236 100542 159248
rect 184382 159236 184388 159248
rect 100536 159208 184388 159236
rect 100536 159196 100542 159208
rect 184382 159196 184388 159208
rect 184440 159196 184446 159248
rect 187050 159196 187056 159248
rect 187108 159236 187114 159248
rect 214558 159236 214564 159248
rect 187108 159208 214564 159236
rect 187108 159196 187114 159208
rect 214558 159196 214564 159208
rect 214616 159196 214622 159248
rect 218238 159196 218244 159248
rect 218296 159236 218302 159248
rect 284386 159236 284392 159248
rect 218296 159208 284392 159236
rect 218296 159196 218302 159208
rect 284386 159196 284392 159208
rect 284444 159196 284450 159248
rect 287974 159196 287980 159248
rect 288032 159236 288038 159248
rect 338758 159236 338764 159248
rect 288032 159208 338764 159236
rect 288032 159196 288038 159208
rect 338758 159196 338764 159208
rect 338816 159196 338822 159248
rect 339310 159196 339316 159248
rect 339368 159236 339374 159248
rect 377950 159236 377956 159248
rect 339368 159208 377956 159236
rect 339368 159196 339374 159208
rect 377950 159196 377956 159208
rect 378008 159196 378014 159248
rect 385586 159196 385592 159248
rect 385644 159236 385650 159248
rect 398834 159236 398840 159248
rect 385644 159208 398840 159236
rect 385644 159196 385650 159208
rect 398834 159196 398840 159208
rect 398892 159196 398898 159248
rect 459646 159196 459652 159248
rect 459704 159236 459710 159248
rect 466638 159236 466644 159248
rect 459704 159208 466644 159236
rect 459704 159196 459710 159208
rect 466638 159196 466644 159208
rect 466696 159196 466702 159248
rect 86954 159128 86960 159180
rect 87012 159168 87018 159180
rect 87012 159140 162992 159168
rect 87012 159128 87018 159140
rect 93670 159060 93676 159112
rect 93728 159100 93734 159112
rect 162854 159100 162860 159112
rect 93728 159072 162860 159100
rect 93728 159060 93734 159072
rect 162854 159060 162860 159072
rect 162912 159060 162918 159112
rect 162964 159100 162992 159140
rect 163038 159128 163044 159180
rect 163096 159168 163102 159180
rect 172146 159168 172152 159180
rect 163096 159140 172152 159168
rect 163096 159128 163102 159140
rect 172146 159128 172152 159140
rect 172204 159128 172210 159180
rect 193766 159128 193772 159180
rect 193824 159168 193830 159180
rect 218054 159168 218060 159180
rect 193824 159140 218060 159168
rect 193824 159128 193830 159140
rect 218054 159128 218060 159140
rect 218112 159128 218118 159180
rect 220722 159128 220728 159180
rect 220780 159168 220786 159180
rect 283190 159168 283196 159180
rect 220780 159140 283196 159168
rect 220780 159128 220786 159140
rect 283190 159128 283196 159140
rect 283248 159128 283254 159180
rect 284662 159128 284668 159180
rect 284720 159168 284726 159180
rect 285766 159168 285772 159180
rect 284720 159140 285772 159168
rect 284720 159128 284726 159140
rect 285766 159128 285772 159140
rect 285824 159128 285830 159180
rect 288158 159168 288164 159180
rect 287026 159140 288164 159168
rect 169754 159100 169760 159112
rect 162964 159072 169760 159100
rect 169754 159060 169760 159072
rect 169812 159060 169818 159112
rect 171778 159060 171784 159112
rect 171836 159100 171842 159112
rect 176654 159100 176660 159112
rect 171836 159072 176660 159100
rect 171836 159060 171842 159072
rect 176654 159060 176660 159072
rect 176712 159060 176718 159112
rect 180334 159060 180340 159112
rect 180392 159100 180398 159112
rect 204898 159100 204904 159112
rect 180392 159072 204904 159100
rect 180392 159060 180398 159072
rect 204898 159060 204904 159072
rect 204956 159060 204962 159112
rect 224126 159060 224132 159112
rect 224184 159100 224190 159112
rect 287026 159100 287054 159140
rect 288158 159128 288164 159140
rect 288216 159128 288222 159180
rect 288894 159128 288900 159180
rect 288952 159168 288958 159180
rect 338390 159168 338396 159180
rect 288952 159140 338396 159168
rect 288952 159128 288958 159140
rect 338390 159128 338396 159140
rect 338448 159128 338454 159180
rect 338482 159128 338488 159180
rect 338540 159168 338546 159180
rect 339678 159168 339684 159180
rect 338540 159140 339684 159168
rect 338540 159128 338546 159140
rect 339678 159128 339684 159140
rect 339736 159128 339742 159180
rect 341886 159128 341892 159180
rect 341944 159168 341950 159180
rect 378226 159168 378232 159180
rect 341944 159140 378232 159168
rect 341944 159128 341950 159140
rect 378226 159128 378232 159140
rect 378284 159128 378290 159180
rect 383102 159128 383108 159180
rect 383160 159168 383166 159180
rect 383160 159140 391244 159168
rect 383160 159128 383166 159140
rect 224184 159072 287054 159100
rect 224184 159060 224190 159072
rect 302234 159060 302240 159112
rect 302292 159100 302298 159112
rect 303522 159100 303528 159112
rect 302292 159072 303528 159100
rect 302292 159060 302298 159072
rect 303522 159060 303528 159072
rect 303580 159060 303586 159112
rect 309042 159060 309048 159112
rect 309100 159100 309106 159112
rect 349798 159100 349804 159112
rect 309100 159072 349804 159100
rect 309100 159060 309106 159072
rect 349798 159060 349804 159072
rect 349856 159060 349862 159112
rect 353202 159100 353208 159112
rect 349908 159072 353208 159100
rect 107194 158992 107200 159044
rect 107252 159032 107258 159044
rect 183462 159032 183468 159044
rect 107252 159004 183468 159032
rect 107252 158992 107258 159004
rect 183462 158992 183468 159004
rect 183520 158992 183526 159044
rect 183738 158992 183744 159044
rect 183796 159032 183802 159044
rect 201402 159032 201408 159044
rect 183796 159004 201408 159032
rect 183796 158992 183802 159004
rect 201402 158992 201408 159004
rect 201460 158992 201466 159044
rect 203886 158992 203892 159044
rect 203944 159032 203950 159044
rect 212718 159032 212724 159044
rect 203944 159004 212724 159032
rect 203944 158992 203950 159004
rect 212718 158992 212724 159004
rect 212776 158992 212782 159044
rect 230842 158992 230848 159044
rect 230900 159032 230906 159044
rect 295150 159032 295156 159044
rect 230900 159004 295156 159032
rect 230900 158992 230906 159004
rect 295150 158992 295156 159004
rect 295208 158992 295214 159044
rect 298094 158992 298100 159044
rect 298152 159032 298158 159044
rect 299566 159032 299572 159044
rect 298152 159004 299572 159032
rect 298152 158992 298158 159004
rect 299566 158992 299572 159004
rect 299624 158992 299630 159044
rect 305362 159032 305368 159044
rect 301056 159004 305368 159032
rect 96246 158924 96252 158976
rect 96304 158964 96310 158976
rect 121914 158964 121920 158976
rect 96304 158936 121920 158964
rect 96304 158924 96310 158936
rect 121914 158924 121920 158936
rect 121972 158924 121978 158976
rect 124030 158924 124036 158976
rect 124088 158964 124094 158976
rect 194134 158964 194140 158976
rect 124088 158936 194140 158964
rect 124088 158924 124094 158936
rect 194134 158924 194140 158936
rect 194192 158924 194198 158976
rect 194686 158924 194692 158976
rect 194744 158964 194750 158976
rect 204162 158964 204168 158976
rect 194744 158936 204168 158964
rect 194744 158924 194750 158936
rect 204162 158924 204168 158936
rect 204220 158924 204226 158976
rect 207290 158924 207296 158976
rect 207348 158964 207354 158976
rect 230750 158964 230756 158976
rect 207348 158936 230756 158964
rect 207348 158924 207354 158936
rect 230750 158924 230756 158936
rect 230808 158924 230814 158976
rect 237558 158924 237564 158976
rect 237616 158964 237622 158976
rect 299474 158964 299480 158976
rect 237616 158936 299480 158964
rect 237616 158924 237622 158936
rect 299474 158924 299480 158936
rect 299532 158924 299538 158976
rect 102962 158856 102968 158908
rect 103020 158896 103026 158908
rect 125502 158896 125508 158908
rect 103020 158868 125508 158896
rect 103020 158856 103026 158868
rect 125502 158856 125508 158868
rect 125560 158856 125566 158908
rect 126330 158856 126336 158908
rect 126388 158896 126394 158908
rect 129734 158896 129740 158908
rect 126388 158868 129740 158896
rect 126388 158856 126394 158868
rect 129734 158856 129740 158868
rect 129792 158856 129798 158908
rect 137094 158896 137100 158908
rect 133156 158868 137100 158896
rect 109678 158788 109684 158840
rect 109736 158828 109742 158840
rect 133156 158828 133184 158868
rect 137094 158856 137100 158868
rect 137152 158856 137158 158908
rect 137186 158856 137192 158908
rect 137244 158896 137250 158908
rect 195422 158896 195428 158908
rect 137244 158868 195428 158896
rect 137244 158856 137250 158868
rect 195422 158856 195428 158868
rect 195480 158856 195486 158908
rect 210602 158856 210608 158908
rect 210660 158896 210666 158908
rect 215386 158896 215392 158908
rect 210660 158868 215392 158896
rect 210660 158856 210666 158868
rect 215386 158856 215392 158868
rect 215444 158856 215450 158908
rect 217318 158856 217324 158908
rect 217376 158896 217382 158908
rect 220354 158896 220360 158908
rect 217376 158868 220360 158896
rect 217376 158856 217382 158868
rect 220354 158856 220360 158868
rect 220412 158856 220418 158908
rect 238386 158856 238392 158908
rect 238444 158896 238450 158908
rect 242434 158896 242440 158908
rect 238444 158868 242440 158896
rect 238444 158856 238450 158868
rect 242434 158856 242440 158868
rect 242492 158856 242498 158908
rect 244274 158856 244280 158908
rect 244332 158896 244338 158908
rect 301056 158896 301084 159004
rect 305362 158992 305368 159004
rect 305420 158992 305426 159044
rect 307386 158992 307392 159044
rect 307444 159032 307450 159044
rect 349908 159032 349936 159072
rect 353202 159060 353208 159072
rect 353260 159060 353266 159112
rect 357802 159060 357808 159112
rect 357860 159100 357866 159112
rect 384942 159100 384948 159112
rect 357860 159072 384948 159100
rect 357860 159060 357866 159072
rect 384942 159060 384948 159072
rect 385000 159060 385006 159112
rect 307444 159004 349936 159032
rect 307444 158992 307450 159004
rect 351086 158992 351092 159044
rect 351144 159032 351150 159044
rect 382550 159032 382556 159044
rect 351144 159004 382556 159032
rect 351144 158992 351150 159004
rect 382550 158992 382556 159004
rect 382608 158992 382614 159044
rect 244332 158868 301084 158896
rect 301516 158936 307524 158964
rect 244332 158856 244338 158868
rect 109736 158800 133184 158828
rect 109736 158788 109742 158800
rect 133230 158788 133236 158840
rect 133288 158828 133294 158840
rect 158714 158828 158720 158840
rect 133288 158800 158720 158828
rect 133288 158788 133294 158800
rect 158714 158788 158720 158800
rect 158772 158788 158778 158840
rect 163498 158788 163504 158840
rect 163556 158828 163562 158840
rect 197262 158828 197268 158840
rect 163556 158800 197268 158828
rect 163556 158788 163562 158800
rect 197262 158788 197268 158800
rect 197320 158788 197326 158840
rect 208118 158788 208124 158840
rect 208176 158828 208182 158840
rect 212442 158828 212448 158840
rect 208176 158800 212448 158828
rect 208176 158788 208182 158800
rect 212442 158788 212448 158800
rect 212500 158788 212506 158840
rect 214834 158788 214840 158840
rect 214892 158828 214898 158840
rect 221458 158828 221464 158840
rect 214892 158800 221464 158828
rect 214892 158788 214898 158800
rect 221458 158788 221464 158800
rect 221516 158788 221522 158840
rect 221550 158788 221556 158840
rect 221608 158828 221614 158840
rect 224586 158828 224592 158840
rect 221608 158800 224592 158828
rect 221608 158788 221614 158800
rect 224586 158788 224592 158800
rect 224644 158788 224650 158840
rect 248506 158788 248512 158840
rect 248564 158828 248570 158840
rect 301516 158828 301544 158936
rect 305638 158856 305644 158908
rect 305696 158896 305702 158908
rect 307386 158896 307392 158908
rect 305696 158868 307392 158896
rect 305696 158856 305702 158868
rect 307386 158856 307392 158868
rect 307444 158856 307450 158908
rect 307496 158896 307524 158936
rect 308214 158924 308220 158976
rect 308272 158964 308278 158976
rect 347682 158964 347688 158976
rect 308272 158936 347688 158964
rect 308272 158924 308278 158936
rect 347682 158924 347688 158936
rect 347740 158924 347746 158976
rect 347774 158924 347780 158976
rect 347832 158964 347838 158976
rect 378778 158964 378784 158976
rect 347832 158936 378784 158964
rect 347832 158924 347838 158936
rect 378778 158924 378784 158936
rect 378836 158924 378842 158976
rect 384758 158924 384764 158976
rect 384816 158964 384822 158976
rect 391216 158964 391244 159140
rect 392302 159128 392308 159180
rect 392360 159168 392366 159180
rect 404262 159168 404268 159180
rect 392360 159140 404268 159168
rect 392360 159128 392366 159140
rect 404262 159128 404268 159140
rect 404320 159128 404326 159180
rect 462958 159128 462964 159180
rect 463016 159168 463022 159180
rect 469214 159168 469220 159180
rect 463016 159140 469220 159168
rect 463016 159128 463022 159140
rect 469214 159128 469220 159140
rect 469272 159128 469278 159180
rect 395706 159060 395712 159112
rect 395764 159100 395770 159112
rect 405642 159100 405648 159112
rect 395764 159072 405648 159100
rect 395764 159060 395770 159072
rect 405642 159060 405648 159072
rect 405700 159060 405706 159112
rect 457898 159060 457904 159112
rect 457956 159100 457962 159112
rect 464522 159100 464528 159112
rect 457956 159072 464528 159100
rect 457956 159060 457962 159072
rect 464522 159060 464528 159072
rect 464580 159060 464586 159112
rect 471422 159060 471428 159112
rect 471480 159100 471486 159112
rect 477678 159100 477684 159112
rect 471480 159072 477684 159100
rect 471480 159060 471486 159072
rect 477678 159060 477684 159072
rect 477736 159060 477742 159112
rect 395154 158992 395160 159044
rect 395212 159032 395218 159044
rect 404170 159032 404176 159044
rect 395212 159004 404176 159032
rect 395212 158992 395218 159004
rect 404170 158992 404176 159004
rect 404228 158992 404234 159044
rect 460474 158992 460480 159044
rect 460532 159032 460538 159044
rect 466454 159032 466460 159044
rect 460532 159004 466460 159032
rect 460532 158992 460538 159004
rect 466454 158992 466460 159004
rect 466512 158992 466518 159044
rect 473906 158992 473912 159044
rect 473964 159032 473970 159044
rect 480254 159032 480260 159044
rect 473964 159004 480260 159032
rect 473964 158992 473970 159004
rect 480254 158992 480260 159004
rect 480312 158992 480318 159044
rect 411346 158964 411352 158976
rect 384816 158936 389036 158964
rect 391216 158936 411352 158964
rect 384816 158924 384822 158936
rect 308582 158896 308588 158908
rect 307496 158868 308588 158896
rect 308582 158856 308588 158868
rect 308640 158856 308646 158908
rect 312446 158856 312452 158908
rect 312504 158896 312510 158908
rect 313642 158896 313648 158908
rect 312504 158868 313648 158896
rect 312504 158856 312510 158868
rect 313642 158856 313648 158868
rect 313700 158856 313706 158908
rect 314930 158856 314936 158908
rect 314988 158896 314994 158908
rect 357434 158896 357440 158908
rect 314988 158868 357440 158896
rect 314988 158856 314994 158868
rect 357434 158856 357440 158868
rect 357492 158856 357498 158908
rect 361206 158856 361212 158908
rect 361264 158896 361270 158908
rect 386322 158896 386328 158908
rect 361264 158868 386328 158896
rect 361264 158856 361270 158868
rect 386322 158856 386328 158868
rect 386380 158856 386386 158908
rect 248564 158800 301544 158828
rect 248564 158788 248570 158800
rect 310698 158788 310704 158840
rect 310756 158828 310762 158840
rect 313182 158828 313188 158840
rect 310756 158800 313188 158828
rect 310756 158788 310762 158800
rect 313182 158788 313188 158800
rect 313240 158788 313246 158840
rect 319162 158788 319168 158840
rect 319220 158828 319226 158840
rect 321554 158828 321560 158840
rect 319220 158800 321560 158828
rect 319220 158788 319226 158800
rect 321554 158788 321560 158800
rect 321612 158788 321618 158840
rect 321646 158788 321652 158840
rect 321704 158828 321710 158840
rect 363138 158828 363144 158840
rect 321704 158800 363144 158828
rect 321704 158788 321710 158800
rect 363138 158788 363144 158800
rect 363196 158788 363202 158840
rect 367922 158788 367928 158840
rect 367980 158828 367986 158840
rect 385034 158828 385040 158840
rect 367980 158800 385040 158828
rect 367980 158788 367986 158800
rect 385034 158788 385040 158800
rect 385092 158788 385098 158840
rect 90358 158720 90364 158772
rect 90416 158760 90422 158772
rect 92474 158760 92480 158772
rect 90416 158732 92480 158760
rect 90416 158720 90422 158732
rect 92474 158720 92480 158732
rect 92532 158720 92538 158772
rect 92842 158720 92848 158772
rect 92900 158760 92906 158772
rect 114462 158760 114468 158772
rect 92900 158732 114468 158760
rect 92900 158720 92906 158732
rect 114462 158720 114468 158732
rect 114520 158720 114526 158772
rect 119798 158720 119804 158772
rect 119856 158760 119862 158772
rect 146570 158760 146576 158772
rect 119856 158732 146576 158760
rect 119856 158720 119862 158732
rect 146570 158720 146576 158732
rect 146628 158720 146634 158772
rect 146662 158720 146668 158772
rect 146720 158760 146726 158772
rect 171778 158760 171784 158772
rect 146720 158732 171784 158760
rect 146720 158720 146726 158732
rect 171778 158720 171784 158732
rect 171836 158720 171842 158772
rect 173618 158720 173624 158772
rect 173676 158760 173682 158772
rect 197354 158760 197360 158772
rect 173676 158732 197360 158760
rect 173676 158720 173682 158732
rect 197354 158720 197360 158732
rect 197412 158720 197418 158772
rect 200574 158720 200580 158772
rect 200632 158760 200638 158772
rect 224954 158760 224960 158772
rect 200632 158732 224960 158760
rect 200632 158720 200638 158732
rect 224954 158720 224960 158732
rect 225012 158720 225018 158772
rect 240870 158720 240876 158772
rect 240928 158760 240934 158772
rect 243354 158760 243360 158772
rect 240928 158732 243360 158760
rect 240928 158720 240934 158732
rect 243354 158720 243360 158732
rect 243412 158720 243418 158772
rect 254394 158720 254400 158772
rect 254452 158760 254458 158772
rect 255406 158760 255412 158772
rect 254452 158732 255412 158760
rect 254452 158720 254458 158732
rect 255406 158720 255412 158732
rect 255464 158720 255470 158772
rect 258534 158720 258540 158772
rect 258592 158760 258598 158772
rect 260926 158760 260932 158772
rect 258592 158732 260932 158760
rect 258592 158720 258598 158732
rect 260926 158720 260932 158732
rect 260984 158720 260990 158772
rect 264422 158720 264428 158772
rect 264480 158760 264486 158772
rect 266354 158760 266360 158772
rect 264480 158732 266360 158760
rect 264480 158720 264486 158732
rect 266354 158720 266360 158732
rect 266412 158720 266418 158772
rect 267826 158720 267832 158772
rect 267884 158760 267890 158772
rect 320266 158760 320272 158772
rect 267884 158732 320272 158760
rect 267884 158720 267890 158732
rect 320266 158720 320272 158732
rect 320324 158720 320330 158772
rect 327534 158720 327540 158772
rect 327592 158760 327598 158772
rect 367186 158760 367192 158772
rect 327592 158732 367192 158760
rect 327592 158720 327598 158732
rect 367186 158720 367192 158732
rect 367244 158720 367250 158772
rect 374638 158720 374644 158772
rect 374696 158760 374702 158772
rect 388438 158760 388444 158772
rect 374696 158732 388444 158760
rect 374696 158720 374702 158732
rect 388438 158720 388444 158732
rect 388496 158720 388502 158772
rect 389008 158760 389036 158936
rect 411346 158924 411352 158936
rect 411404 158924 411410 158976
rect 416682 158924 416688 158976
rect 416740 158964 416746 158976
rect 419534 158964 419540 158976
rect 416740 158936 419540 158964
rect 416740 158924 416746 158936
rect 419534 158924 419540 158936
rect 419592 158924 419598 158976
rect 420086 158924 420092 158976
rect 420144 158964 420150 158976
rect 423582 158964 423588 158976
rect 420144 158936 423588 158964
rect 420144 158924 420150 158936
rect 423582 158924 423588 158936
rect 423640 158924 423646 158976
rect 456242 158924 456248 158976
rect 456300 158964 456306 158976
rect 463142 158964 463148 158976
rect 456300 158936 463148 158964
rect 456300 158924 456306 158936
rect 463142 158924 463148 158936
rect 463200 158924 463206 158976
rect 466362 158924 466368 158976
rect 466420 158964 466426 158976
rect 472342 158964 472348 158976
rect 466420 158936 472348 158964
rect 466420 158924 466426 158936
rect 472342 158924 472348 158936
rect 472400 158924 472406 158976
rect 475562 158924 475568 158976
rect 475620 158964 475626 158976
rect 482002 158964 482008 158976
rect 475620 158936 482008 158964
rect 475620 158924 475626 158936
rect 482002 158924 482008 158936
rect 482060 158924 482066 158976
rect 412542 158856 412548 158908
rect 412600 158896 412606 158908
rect 412818 158896 412824 158908
rect 412600 158868 412824 158896
rect 412600 158856 412606 158868
rect 412818 158856 412824 158868
rect 412876 158856 412882 158908
rect 454586 158856 454592 158908
rect 454644 158896 454650 158908
rect 461670 158896 461676 158908
rect 454644 158868 461676 158896
rect 454644 158856 454650 158868
rect 461670 158856 461676 158868
rect 461728 158856 461734 158908
rect 465534 158856 465540 158908
rect 465592 158896 465598 158908
rect 472158 158896 472164 158908
rect 465592 158868 472164 158896
rect 465592 158856 465598 158868
rect 472158 158856 472164 158868
rect 472216 158856 472222 158908
rect 474734 158856 474740 158908
rect 474792 158896 474798 158908
rect 481358 158896 481364 158908
rect 474792 158868 481364 158896
rect 474792 158856 474798 158868
rect 481358 158856 481364 158868
rect 481416 158856 481422 158908
rect 508314 158856 508320 158908
rect 508372 158896 508378 158908
rect 510062 158896 510068 158908
rect 508372 158868 510068 158896
rect 508372 158856 508378 158868
rect 510062 158856 510068 158868
rect 510120 158856 510126 158908
rect 389082 158788 389088 158840
rect 389140 158828 389146 158840
rect 390370 158828 390376 158840
rect 389140 158800 390376 158828
rect 389140 158788 389146 158800
rect 390370 158788 390376 158800
rect 390428 158788 390434 158840
rect 409138 158788 409144 158840
rect 409196 158828 409202 158840
rect 410702 158828 410708 158840
rect 409196 158800 410708 158828
rect 409196 158788 409202 158800
rect 410702 158788 410708 158800
rect 410760 158788 410766 158840
rect 455414 158788 455420 158840
rect 455472 158828 455478 158840
rect 463602 158828 463608 158840
rect 455472 158800 463608 158828
rect 455472 158788 455478 158800
rect 463602 158788 463608 158800
rect 463660 158788 463666 158840
rect 464614 158788 464620 158840
rect 464672 158828 464678 158840
rect 471422 158828 471428 158840
rect 464672 158800 471428 158828
rect 464672 158788 464678 158800
rect 471422 158788 471428 158800
rect 471480 158788 471486 158840
rect 476390 158788 476396 158840
rect 476448 158828 476454 158840
rect 481634 158828 481640 158840
rect 476448 158800 481640 158828
rect 476448 158788 476454 158800
rect 481634 158788 481640 158800
rect 481692 158788 481698 158840
rect 506382 158788 506388 158840
rect 506440 158828 506446 158840
rect 507578 158828 507584 158840
rect 506440 158800 507584 158828
rect 506440 158788 506446 158800
rect 507578 158788 507584 158800
rect 507636 158788 507642 158840
rect 389174 158760 389180 158772
rect 389008 158732 389180 158760
rect 389174 158720 389180 158732
rect 389232 158720 389238 158772
rect 405734 158720 405740 158772
rect 405792 158760 405798 158772
rect 409230 158760 409236 158772
rect 405792 158732 409236 158760
rect 405792 158720 405798 158732
rect 409230 158720 409236 158732
rect 409288 158720 409294 158772
rect 452838 158720 452844 158772
rect 452896 158760 452902 158772
rect 459554 158760 459560 158772
rect 452896 158732 459560 158760
rect 452896 158720 452902 158732
rect 459554 158720 459560 158732
rect 459612 158720 459618 158772
rect 463786 158720 463792 158772
rect 463844 158760 463850 158772
rect 471790 158760 471796 158772
rect 463844 158732 471796 158760
rect 463844 158720 463850 158732
rect 471790 158720 471796 158732
rect 471848 158720 471854 158772
rect 473078 158720 473084 158772
rect 473136 158760 473142 158772
rect 478966 158760 478972 158772
rect 473136 158732 478972 158760
rect 473136 158720 473142 158732
rect 478966 158720 478972 158732
rect 479024 158720 479030 158772
rect 482278 158720 482284 158772
rect 482336 158760 482342 158772
rect 487246 158760 487252 158772
rect 482336 158732 487252 158760
rect 482336 158720 482342 158732
rect 487246 158720 487252 158732
rect 487304 158720 487310 158772
rect 505278 158720 505284 158772
rect 505336 158760 505342 158772
rect 506750 158760 506756 158772
rect 505336 158732 506756 158760
rect 505336 158720 505342 158732
rect 506750 158720 506756 158732
rect 506808 158720 506814 158772
rect 507026 158720 507032 158772
rect 507084 158760 507090 158772
rect 508406 158760 508412 158772
rect 507084 158732 508412 158760
rect 507084 158720 507090 158732
rect 508406 158720 508412 158732
rect 508464 158720 508470 158772
rect 509418 158720 509424 158772
rect 509476 158760 509482 158772
rect 511718 158760 511724 158772
rect 509476 158732 511724 158760
rect 509476 158720 509482 158732
rect 511718 158720 511724 158732
rect 511776 158720 511782 158772
rect 514938 158720 514944 158772
rect 514996 158760 515002 158772
rect 518526 158760 518532 158772
rect 514996 158732 518532 158760
rect 514996 158720 515002 158732
rect 518526 158720 518532 158732
rect 518584 158720 518590 158772
rect 81066 158652 81072 158704
rect 81124 158692 81130 158704
rect 180886 158692 180892 158704
rect 81124 158664 180892 158692
rect 81124 158652 81130 158664
rect 180886 158652 180892 158664
rect 180944 158652 180950 158704
rect 181990 158652 181996 158704
rect 182048 158692 182054 158704
rect 256786 158692 256792 158704
rect 182048 158664 256792 158692
rect 182048 158652 182054 158664
rect 256786 158652 256792 158664
rect 256844 158652 256850 158704
rect 67634 158584 67640 158636
rect 67692 158624 67698 158636
rect 166074 158624 166080 158636
rect 67692 158596 166080 158624
rect 67692 158584 67698 158596
rect 166074 158584 166080 158596
rect 166132 158584 166138 158636
rect 166534 158584 166540 158636
rect 166592 158624 166598 158636
rect 172974 158624 172980 158636
rect 166592 158596 172980 158624
rect 166592 158584 166598 158596
rect 172974 158584 172980 158596
rect 173032 158584 173038 158636
rect 173342 158584 173348 158636
rect 173400 158624 173406 158636
rect 247126 158624 247132 158636
rect 173400 158596 247132 158624
rect 173400 158584 173406 158596
rect 247126 158584 247132 158596
rect 247184 158584 247190 158636
rect 74350 158516 74356 158568
rect 74408 158556 74414 158568
rect 172882 158556 172888 158568
rect 74408 158528 172888 158556
rect 74408 158516 74414 158528
rect 172882 158516 172888 158528
rect 172940 158516 172946 158568
rect 178678 158516 178684 158568
rect 178736 158556 178742 158568
rect 255590 158556 255596 158568
rect 178736 158528 255596 158556
rect 178736 158516 178742 158528
rect 255590 158516 255596 158528
rect 255648 158516 255654 158568
rect 71038 158448 71044 158500
rect 71096 158488 71102 158500
rect 165982 158488 165988 158500
rect 71096 158460 165988 158488
rect 71096 158448 71102 158460
rect 165982 158448 165988 158460
rect 166040 158448 166046 158500
rect 166442 158448 166448 158500
rect 166500 158488 166506 158500
rect 170398 158488 170404 158500
rect 166500 158460 170404 158488
rect 166500 158448 166506 158460
rect 170398 158448 170404 158460
rect 170456 158448 170462 158500
rect 173158 158448 173164 158500
rect 173216 158488 173222 158500
rect 175182 158488 175188 158500
rect 173216 158460 175188 158488
rect 173216 158448 173222 158460
rect 175182 158448 175188 158460
rect 175240 158448 175246 158500
rect 175274 158448 175280 158500
rect 175332 158488 175338 158500
rect 252738 158488 252744 158500
rect 175332 158460 252744 158488
rect 175332 158448 175338 158460
rect 252738 158448 252744 158460
rect 252796 158448 252802 158500
rect 64230 158380 64236 158432
rect 64288 158420 64294 158432
rect 167546 158420 167552 158432
rect 64288 158392 167552 158420
rect 64288 158380 64294 158392
rect 167546 158380 167552 158392
rect 167604 158380 167610 158432
rect 171962 158380 171968 158432
rect 172020 158420 172026 158432
rect 250070 158420 250076 158432
rect 172020 158392 250076 158420
rect 172020 158380 172026 158392
rect 250070 158380 250076 158392
rect 250128 158380 250134 158432
rect 60918 158312 60924 158364
rect 60976 158352 60982 158364
rect 164326 158352 164332 158364
rect 60976 158324 164332 158352
rect 60976 158312 60982 158324
rect 164326 158312 164332 158324
rect 164384 158312 164390 158364
rect 165246 158312 165252 158364
rect 165304 158352 165310 158364
rect 245010 158352 245016 158364
rect 165304 158324 245016 158352
rect 165304 158312 165310 158324
rect 245010 158312 245016 158324
rect 245068 158312 245074 158364
rect 54202 158244 54208 158296
rect 54260 158284 54266 158296
rect 160278 158284 160284 158296
rect 54260 158256 160284 158284
rect 54260 158244 54266 158256
rect 160278 158244 160284 158256
rect 160336 158244 160342 158296
rect 161842 158244 161848 158296
rect 161900 158284 161906 158296
rect 242066 158284 242072 158296
rect 161900 158256 242072 158284
rect 161900 158244 161906 158256
rect 242066 158244 242072 158256
rect 242124 158244 242130 158296
rect 50798 158176 50804 158228
rect 50856 158216 50862 158228
rect 157702 158216 157708 158228
rect 50856 158188 157708 158216
rect 50856 158176 50862 158188
rect 157702 158176 157708 158188
rect 157760 158176 157766 158228
rect 158438 158176 158444 158228
rect 158496 158216 158502 158228
rect 238938 158216 238944 158228
rect 158496 158188 238944 158216
rect 158496 158176 158502 158188
rect 238938 158176 238944 158188
rect 238996 158176 239002 158228
rect 256878 158176 256884 158228
rect 256936 158216 256942 158228
rect 315022 158216 315028 158228
rect 256936 158188 315028 158216
rect 256936 158176 256942 158188
rect 315022 158176 315028 158188
rect 315080 158176 315086 158228
rect 47486 158108 47492 158160
rect 47544 158148 47550 158160
rect 155034 158148 155040 158160
rect 47544 158120 155040 158148
rect 47544 158108 47550 158120
rect 155034 158108 155040 158120
rect 155092 158108 155098 158160
rect 155126 158108 155132 158160
rect 155184 158148 155190 158160
rect 237374 158148 237380 158160
rect 155184 158120 237380 158148
rect 155184 158108 155190 158120
rect 237374 158108 237380 158120
rect 237432 158108 237438 158160
rect 246758 158108 246764 158160
rect 246816 158148 246822 158160
rect 306926 158148 306932 158160
rect 246816 158120 306932 158148
rect 246816 158108 246822 158120
rect 306926 158108 306932 158120
rect 306984 158108 306990 158160
rect 37366 158040 37372 158092
rect 37424 158080 37430 158092
rect 146386 158080 146392 158092
rect 37424 158052 146392 158080
rect 37424 158040 37430 158052
rect 146386 158040 146392 158052
rect 146444 158040 146450 158092
rect 148410 158040 148416 158092
rect 148468 158080 148474 158092
rect 231946 158080 231952 158092
rect 148468 158052 231952 158080
rect 148468 158040 148474 158052
rect 231946 158040 231952 158052
rect 232004 158040 232010 158092
rect 243446 158040 243452 158092
rect 243504 158080 243510 158092
rect 304718 158080 304724 158092
rect 243504 158052 304724 158080
rect 243504 158040 243510 158052
rect 304718 158040 304724 158052
rect 304776 158040 304782 158092
rect 382 157972 388 158024
rect 440 158012 446 158024
rect 118878 158012 118884 158024
rect 440 157984 118884 158012
rect 440 157972 446 157984
rect 118878 157972 118884 157984
rect 118936 157972 118942 158024
rect 131574 157972 131580 158024
rect 131632 158012 131638 158024
rect 219342 158012 219348 158024
rect 131632 157984 219348 158012
rect 131632 157972 131638 157984
rect 219342 157972 219348 157984
rect 219400 157972 219406 158024
rect 236730 157972 236736 158024
rect 236788 158012 236794 158024
rect 299658 158012 299664 158024
rect 236788 157984 299664 158012
rect 236788 157972 236794 157984
rect 299658 157972 299664 157984
rect 299716 157972 299722 158024
rect 77754 157904 77760 157956
rect 77812 157944 77818 157956
rect 77812 157916 170168 157944
rect 77812 157904 77818 157916
rect 87782 157836 87788 157888
rect 87840 157876 87846 157888
rect 164878 157876 164884 157888
rect 87840 157848 164884 157876
rect 87840 157836 87846 157848
rect 164878 157836 164884 157848
rect 164936 157836 164942 157888
rect 84470 157768 84476 157820
rect 84528 157808 84534 157820
rect 170030 157808 170036 157820
rect 84528 157780 170036 157808
rect 84528 157768 84534 157780
rect 170030 157768 170036 157780
rect 170088 157768 170094 157820
rect 170140 157808 170168 157916
rect 170214 157904 170220 157956
rect 170272 157944 170278 157956
rect 182266 157944 182272 157956
rect 170272 157916 182272 157944
rect 170272 157904 170278 157916
rect 182266 157904 182272 157916
rect 182324 157904 182330 157956
rect 185302 157944 185308 157956
rect 185228 157916 185308 157944
rect 170490 157836 170496 157888
rect 170548 157876 170554 157888
rect 185118 157876 185124 157888
rect 170548 157848 185124 157876
rect 170548 157836 170554 157848
rect 185118 157836 185124 157848
rect 185176 157836 185182 157888
rect 178034 157808 178040 157820
rect 170140 157780 178040 157808
rect 178034 157768 178040 157780
rect 178092 157768 178098 157820
rect 179414 157768 179420 157820
rect 179472 157808 179478 157820
rect 185228 157808 185256 157916
rect 185302 157904 185308 157916
rect 185360 157904 185366 157956
rect 185394 157904 185400 157956
rect 185452 157944 185458 157956
rect 260466 157944 260472 157956
rect 185452 157916 260472 157944
rect 185452 157904 185458 157916
rect 260466 157904 260472 157916
rect 260524 157904 260530 157956
rect 188798 157836 188804 157888
rect 188856 157876 188862 157888
rect 263042 157876 263048 157888
rect 188856 157848 263048 157876
rect 188856 157836 188862 157848
rect 263042 157836 263048 157848
rect 263100 157836 263106 157888
rect 190638 157808 190644 157820
rect 179472 157780 185256 157808
rect 185504 157780 190644 157808
rect 179472 157768 179478 157780
rect 91186 157700 91192 157752
rect 91244 157740 91250 157752
rect 185302 157740 185308 157752
rect 91244 157712 185308 157740
rect 91244 157700 91250 157712
rect 185302 157700 185308 157712
rect 185360 157700 185366 157752
rect 94590 157632 94596 157684
rect 94648 157672 94654 157684
rect 185504 157672 185532 157780
rect 190638 157768 190644 157780
rect 190696 157768 190702 157820
rect 195514 157768 195520 157820
rect 195572 157808 195578 157820
rect 267734 157808 267740 157820
rect 195572 157780 267740 157808
rect 195572 157768 195578 157780
rect 267734 157768 267740 157780
rect 267792 157768 267798 157820
rect 185670 157700 185676 157752
rect 185728 157740 185734 157752
rect 188522 157740 188528 157752
rect 185728 157712 188528 157740
rect 185728 157700 185734 157712
rect 188522 157700 188528 157712
rect 188580 157700 188586 157752
rect 190454 157700 190460 157752
rect 190512 157740 190518 157752
rect 263686 157740 263692 157752
rect 190512 157712 263692 157740
rect 190512 157700 190518 157712
rect 263686 157700 263692 157712
rect 263744 157700 263750 157752
rect 94648 157644 185532 157672
rect 94648 157632 94654 157644
rect 185578 157632 185584 157684
rect 185636 157672 185642 157684
rect 236086 157672 236092 157684
rect 185636 157644 236092 157672
rect 185636 157632 185642 157644
rect 236086 157632 236092 157644
rect 236144 157632 236150 157684
rect 97902 157564 97908 157616
rect 97960 157604 97966 157616
rect 193214 157604 193220 157616
rect 97960 157576 193220 157604
rect 97960 157564 97966 157576
rect 193214 157564 193220 157576
rect 193272 157564 193278 157616
rect 197354 157564 197360 157616
rect 197412 157604 197418 157616
rect 251450 157604 251456 157616
rect 197412 157576 251456 157604
rect 197412 157564 197418 157576
rect 251450 157564 251456 157576
rect 251508 157564 251514 157616
rect 111334 157496 111340 157548
rect 111392 157536 111398 157548
rect 203978 157536 203984 157548
rect 111392 157508 203984 157536
rect 111392 157496 111398 157508
rect 203978 157496 203984 157508
rect 204036 157496 204042 157548
rect 204898 157496 204904 157548
rect 204956 157536 204962 157548
rect 255866 157536 255872 157548
rect 204956 157508 255872 157536
rect 204956 157496 204962 157508
rect 255866 157496 255872 157508
rect 255924 157496 255930 157548
rect 114738 157428 114744 157480
rect 114796 157468 114802 157480
rect 206554 157468 206560 157480
rect 114796 157440 206560 157468
rect 114796 157428 114802 157440
rect 206554 157428 206560 157440
rect 206612 157428 206618 157480
rect 141694 157360 141700 157412
rect 141752 157400 141758 157412
rect 227070 157400 227076 157412
rect 141752 157372 227076 157400
rect 141752 157360 141758 157372
rect 227070 157360 227076 157372
rect 227128 157360 227134 157412
rect 49142 157292 49148 157344
rect 49200 157332 49206 157344
rect 156414 157332 156420 157344
rect 49200 157304 156420 157332
rect 49200 157292 49206 157304
rect 156414 157292 156420 157304
rect 156472 157292 156478 157344
rect 158714 157292 158720 157344
rect 158772 157332 158778 157344
rect 219986 157332 219992 157344
rect 158772 157304 219992 157332
rect 158772 157292 158778 157304
rect 219986 157292 219992 157304
rect 220044 157292 220050 157344
rect 45738 157224 45744 157276
rect 45796 157264 45802 157276
rect 153838 157264 153844 157276
rect 45796 157236 153844 157264
rect 45796 157224 45802 157236
rect 153838 157224 153844 157236
rect 153896 157224 153902 157276
rect 163774 157224 163780 157276
rect 163832 157264 163838 157276
rect 166442 157264 166448 157276
rect 163832 157236 166448 157264
rect 163832 157224 163838 157236
rect 166442 157224 166448 157236
rect 166500 157224 166506 157276
rect 192110 157224 192116 157276
rect 192168 157264 192174 157276
rect 265158 157264 265164 157276
rect 192168 157236 265164 157264
rect 192168 157224 192174 157236
rect 265158 157224 265164 157236
rect 265216 157224 265222 157276
rect 283834 157224 283840 157276
rect 283892 157264 283898 157276
rect 335538 157264 335544 157276
rect 283892 157236 335544 157264
rect 283892 157224 283898 157236
rect 335538 157224 335544 157236
rect 335596 157224 335602 157276
rect 42426 157156 42432 157208
rect 42484 157196 42490 157208
rect 151262 157196 151268 157208
rect 42484 157168 151268 157196
rect 42484 157156 42490 157168
rect 151262 157156 151268 157168
rect 151320 157156 151326 157208
rect 156506 157156 156512 157208
rect 156564 157196 156570 157208
rect 159082 157196 159088 157208
rect 156564 157168 159088 157196
rect 156564 157156 156570 157168
rect 159082 157156 159088 157168
rect 159140 157156 159146 157208
rect 160094 157156 160100 157208
rect 160152 157196 160158 157208
rect 166166 157196 166172 157208
rect 160152 157168 166172 157196
rect 160152 157156 160158 157168
rect 166166 157156 166172 157168
rect 166224 157156 166230 157208
rect 166258 157156 166264 157208
rect 166316 157196 166322 157208
rect 171134 157196 171140 157208
rect 166316 157168 171140 157196
rect 166316 157156 166322 157168
rect 171134 157156 171140 157168
rect 171192 157156 171198 157208
rect 177022 157156 177028 157208
rect 177080 157196 177086 157208
rect 254026 157196 254032 157208
rect 177080 157168 254032 157196
rect 177080 157156 177086 157168
rect 254026 157156 254032 157168
rect 254084 157156 254090 157208
rect 300670 157156 300676 157208
rect 300728 157196 300734 157208
rect 348050 157196 348056 157208
rect 300728 157168 348056 157196
rect 300728 157156 300734 157168
rect 348050 157156 348056 157168
rect 348108 157156 348114 157208
rect 39022 157088 39028 157140
rect 39080 157128 39086 157140
rect 148778 157128 148784 157140
rect 39080 157100 148784 157128
rect 39080 157088 39086 157100
rect 148778 157088 148784 157100
rect 148836 157088 148842 157140
rect 150066 157088 150072 157140
rect 150124 157128 150130 157140
rect 233510 157128 233516 157140
rect 150124 157100 233516 157128
rect 150124 157088 150130 157100
rect 233510 157088 233516 157100
rect 233568 157088 233574 157140
rect 280430 157088 280436 157140
rect 280488 157128 280494 157140
rect 333054 157128 333060 157140
rect 280488 157100 333060 157128
rect 280488 157088 280494 157100
rect 333054 157088 333060 157100
rect 333112 157088 333118 157140
rect 35710 157020 35716 157072
rect 35768 157060 35774 157072
rect 146202 157060 146208 157072
rect 35768 157032 146208 157060
rect 35768 157020 35774 157032
rect 146202 157020 146208 157032
rect 146260 157020 146266 157072
rect 151722 157020 151728 157072
rect 151780 157060 151786 157072
rect 234798 157060 234804 157072
rect 151780 157032 234804 157060
rect 151780 157020 151786 157032
rect 234798 157020 234804 157032
rect 234856 157020 234862 157072
rect 273714 157020 273720 157072
rect 273772 157060 273778 157072
rect 327902 157060 327908 157072
rect 273772 157032 327908 157060
rect 273772 157020 273778 157032
rect 327902 157020 327908 157032
rect 327960 157020 327966 157072
rect 24762 156952 24768 157004
rect 24820 156992 24826 157004
rect 137370 156992 137376 157004
rect 24820 156964 137376 156992
rect 24820 156952 24826 156964
rect 137370 156952 137376 156964
rect 137428 156952 137434 157004
rect 138290 156952 138296 157004
rect 138348 156992 138354 157004
rect 224126 156992 224132 157004
rect 138348 156964 224132 156992
rect 138348 156952 138354 156964
rect 224126 156952 224132 156964
rect 224184 156952 224190 157004
rect 224954 156952 224960 157004
rect 225012 156992 225018 157004
rect 272058 156992 272064 157004
rect 225012 156964 272064 156992
rect 225012 156952 225018 156964
rect 272058 156952 272064 156964
rect 272116 156952 272122 157004
rect 277118 156952 277124 157004
rect 277176 156992 277182 157004
rect 330478 156992 330484 157004
rect 277176 156964 330484 156992
rect 277176 156952 277182 156964
rect 330478 156952 330484 156964
rect 330536 156952 330542 157004
rect 21358 156884 21364 156936
rect 21416 156924 21422 156936
rect 135254 156924 135260 156936
rect 21416 156896 135260 156924
rect 21416 156884 21422 156896
rect 135254 156884 135260 156896
rect 135312 156884 135318 156936
rect 135806 156884 135812 156936
rect 135864 156924 135870 156936
rect 222562 156924 222568 156936
rect 135864 156896 222568 156924
rect 135864 156884 135870 156896
rect 222562 156884 222568 156896
rect 222620 156884 222626 156936
rect 226610 156884 226616 156936
rect 226668 156924 226674 156936
rect 291930 156924 291936 156936
rect 226668 156896 291936 156924
rect 226668 156884 226674 156896
rect 291930 156884 291936 156896
rect 291988 156884 291994 156936
rect 293862 156884 293868 156936
rect 293920 156924 293926 156936
rect 342714 156924 342720 156936
rect 293920 156896 342720 156924
rect 293920 156884 293926 156896
rect 342714 156884 342720 156896
rect 342772 156884 342778 156936
rect 18046 156816 18052 156868
rect 18104 156856 18110 156868
rect 132494 156856 132500 156868
rect 18104 156828 132500 156856
rect 18104 156816 18110 156828
rect 132494 156816 132500 156828
rect 132552 156816 132558 156868
rect 134886 156816 134892 156868
rect 134944 156856 134950 156868
rect 221366 156856 221372 156868
rect 134944 156828 221372 156856
rect 134944 156816 134950 156828
rect 221366 156816 221372 156828
rect 221424 156816 221430 156868
rect 223206 156816 223212 156868
rect 223264 156856 223270 156868
rect 289354 156856 289360 156868
rect 223264 156828 289360 156856
rect 223264 156816 223270 156828
rect 289354 156816 289360 156828
rect 289412 156816 289418 156868
rect 290550 156816 290556 156868
rect 290608 156856 290614 156868
rect 340046 156856 340052 156868
rect 290608 156828 340052 156856
rect 290608 156816 290614 156828
rect 340046 156816 340052 156828
rect 340104 156816 340110 156868
rect 14642 156748 14648 156800
rect 14700 156788 14706 156800
rect 130102 156788 130108 156800
rect 14700 156760 130108 156788
rect 14700 156748 14706 156760
rect 130102 156748 130108 156760
rect 130160 156748 130166 156800
rect 139118 156748 139124 156800
rect 139176 156788 139182 156800
rect 225138 156788 225144 156800
rect 139176 156760 225144 156788
rect 139176 156748 139182 156760
rect 225138 156748 225144 156760
rect 225196 156748 225202 156800
rect 230014 156748 230020 156800
rect 230072 156788 230078 156800
rect 294046 156788 294052 156800
rect 230072 156760 294052 156788
rect 230072 156748 230078 156760
rect 294046 156748 294052 156760
rect 294104 156748 294110 156800
rect 297266 156748 297272 156800
rect 297324 156788 297330 156800
rect 345106 156788 345112 156800
rect 297324 156760 345112 156788
rect 297324 156748 297330 156760
rect 345106 156748 345112 156760
rect 345164 156748 345170 156800
rect 11238 156680 11244 156732
rect 11296 156720 11302 156732
rect 127526 156720 127532 156732
rect 11296 156692 127532 156720
rect 11296 156680 11302 156692
rect 127526 156680 127532 156692
rect 127584 156680 127590 156732
rect 128170 156680 128176 156732
rect 128228 156720 128234 156732
rect 212534 156720 212540 156732
rect 128228 156692 212540 156720
rect 128228 156680 128234 156692
rect 212534 156680 212540 156692
rect 212592 156680 212598 156732
rect 215478 156720 215484 156732
rect 212644 156692 215484 156720
rect 2038 156612 2044 156664
rect 2096 156652 2102 156664
rect 120442 156652 120448 156664
rect 2096 156624 120448 156652
rect 2096 156612 2102 156624
rect 120442 156612 120448 156624
rect 120500 156612 120506 156664
rect 124858 156612 124864 156664
rect 124916 156652 124922 156664
rect 211798 156652 211804 156664
rect 124916 156624 211804 156652
rect 124916 156612 124922 156624
rect 211798 156612 211804 156624
rect 211856 156612 211862 156664
rect 52454 156544 52460 156596
rect 52512 156584 52518 156596
rect 158990 156584 158996 156596
rect 52512 156556 158996 156584
rect 52512 156544 52518 156556
rect 158990 156544 158996 156556
rect 159048 156544 159054 156596
rect 159082 156544 159088 156596
rect 159140 156584 159146 156596
rect 212644 156584 212672 156692
rect 215478 156680 215484 156692
rect 215536 156680 215542 156732
rect 219894 156680 219900 156732
rect 219952 156720 219958 156732
rect 286226 156720 286232 156732
rect 219952 156692 286232 156720
rect 219952 156680 219958 156692
rect 286226 156680 286232 156692
rect 286284 156680 286290 156732
rect 287146 156680 287152 156732
rect 287204 156720 287210 156732
rect 338114 156720 338120 156732
rect 287204 156692 338120 156720
rect 287204 156680 287210 156692
rect 338114 156680 338120 156692
rect 338172 156680 338178 156732
rect 216490 156612 216496 156664
rect 216548 156652 216554 156664
rect 283098 156652 283104 156664
rect 216548 156624 283104 156652
rect 216548 156612 216554 156624
rect 283098 156612 283104 156624
rect 283156 156612 283162 156664
rect 498286 156612 498292 156664
rect 498344 156652 498350 156664
rect 499298 156652 499304 156664
rect 498344 156624 499304 156652
rect 498344 156612 498350 156624
rect 499298 156612 499304 156624
rect 499356 156612 499362 156664
rect 159140 156556 212672 156584
rect 159140 156544 159146 156556
rect 213822 156544 213828 156596
rect 213880 156584 213886 156596
rect 281626 156584 281632 156596
rect 213880 156556 281632 156584
rect 213880 156544 213886 156556
rect 281626 156544 281632 156556
rect 281684 156544 281690 156596
rect 59262 156476 59268 156528
rect 59320 156516 59326 156528
rect 164142 156516 164148 156528
rect 59320 156488 164148 156516
rect 59320 156476 59326 156488
rect 164142 156476 164148 156488
rect 164200 156476 164206 156528
rect 166166 156476 166172 156528
rect 166224 156516 166230 156528
rect 166224 156488 166396 156516
rect 166224 156476 166230 156488
rect 69290 156408 69296 156460
rect 69348 156448 69354 156460
rect 166258 156448 166264 156460
rect 69348 156420 166264 156448
rect 69348 156408 69354 156420
rect 166258 156408 166264 156420
rect 166316 156408 166322 156460
rect 166368 156448 166396 156488
rect 166442 156476 166448 156528
rect 166500 156516 166506 156528
rect 225046 156516 225052 156528
rect 166500 156488 225052 156516
rect 166500 156476 166506 156488
rect 225046 156476 225052 156488
rect 225104 156476 225110 156528
rect 228358 156448 228364 156460
rect 166368 156420 228364 156448
rect 228358 156408 228364 156420
rect 228416 156408 228422 156460
rect 82814 156340 82820 156392
rect 82872 156380 82878 156392
rect 182082 156380 182088 156392
rect 82872 156352 182088 156380
rect 82872 156340 82878 156352
rect 182082 156340 182088 156352
rect 182140 156340 182146 156392
rect 198826 156340 198832 156392
rect 198884 156380 198890 156392
rect 200850 156380 200856 156392
rect 198884 156352 200856 156380
rect 198884 156340 198890 156352
rect 200850 156340 200856 156352
rect 200908 156340 200914 156392
rect 209774 156340 209780 156392
rect 209832 156380 209838 156392
rect 279050 156380 279056 156392
rect 209832 156352 279056 156380
rect 209832 156340 209838 156352
rect 279050 156340 279056 156352
rect 279108 156340 279114 156392
rect 99558 156272 99564 156324
rect 99616 156312 99622 156324
rect 194962 156312 194968 156324
rect 99616 156284 194968 156312
rect 99616 156272 99622 156284
rect 194962 156272 194968 156284
rect 195020 156272 195026 156324
rect 209130 156312 209136 156324
rect 200592 156284 209136 156312
rect 101306 156204 101312 156256
rect 101364 156244 101370 156256
rect 196250 156244 196256 156256
rect 101364 156216 196256 156244
rect 101364 156204 101370 156216
rect 196250 156204 196256 156216
rect 196308 156204 196314 156256
rect 108022 156136 108028 156188
rect 108080 156176 108086 156188
rect 200390 156176 200396 156188
rect 108080 156148 200396 156176
rect 108080 156136 108086 156148
rect 200390 156136 200396 156148
rect 200448 156136 200454 156188
rect 118142 156068 118148 156120
rect 118200 156108 118206 156120
rect 200592 156108 200620 156284
rect 209130 156272 209136 156284
rect 209188 156272 209194 156324
rect 212534 156272 212540 156324
rect 212592 156312 212598 156324
rect 216766 156312 216772 156324
rect 212592 156284 216772 156312
rect 212592 156272 212598 156284
rect 216766 156272 216772 156284
rect 216824 156272 216830 156324
rect 218054 156272 218060 156324
rect 218112 156312 218118 156324
rect 266906 156312 266912 156324
rect 218112 156284 266912 156312
rect 218112 156272 218118 156284
rect 266906 156272 266912 156284
rect 266964 156272 266970 156324
rect 200666 156204 200672 156256
rect 200724 156244 200730 156256
rect 201310 156244 201316 156256
rect 200724 156216 201316 156244
rect 200724 156204 200730 156216
rect 201310 156204 201316 156216
rect 201368 156204 201374 156256
rect 203058 156204 203064 156256
rect 203116 156244 203122 156256
rect 203116 156216 219434 156244
rect 203116 156204 203122 156216
rect 211614 156176 211620 156188
rect 118200 156080 200620 156108
rect 200776 156148 211620 156176
rect 118200 156068 118206 156080
rect 121454 156000 121460 156052
rect 121512 156040 121518 156052
rect 200776 156040 200804 156148
rect 211614 156136 211620 156148
rect 211672 156136 211678 156188
rect 211798 156136 211804 156188
rect 211856 156176 211862 156188
rect 213914 156176 213920 156188
rect 211856 156148 213920 156176
rect 211856 156136 211862 156148
rect 213914 156136 213920 156148
rect 213972 156136 213978 156188
rect 219406 156176 219434 156216
rect 230750 156204 230756 156256
rect 230808 156244 230814 156256
rect 277118 156244 277124 156256
rect 230808 156216 277124 156244
rect 230808 156204 230814 156216
rect 277118 156204 277124 156216
rect 277176 156204 277182 156256
rect 273898 156176 273904 156188
rect 219406 156148 273904 156176
rect 273898 156136 273904 156148
rect 273956 156136 273962 156188
rect 202322 156068 202328 156120
rect 202380 156108 202386 156120
rect 273254 156108 273260 156120
rect 202380 156080 273260 156108
rect 202380 156068 202386 156080
rect 273254 156068 273260 156080
rect 273312 156068 273318 156120
rect 121512 156012 200804 156040
rect 121512 156000 121518 156012
rect 200850 156000 200856 156052
rect 200908 156040 200914 156052
rect 270494 156040 270500 156052
rect 200908 156012 270500 156040
rect 200908 156000 200914 156012
rect 270494 156000 270500 156012
rect 270552 156000 270558 156052
rect 145006 155932 145012 155984
rect 145064 155972 145070 155984
rect 229646 155972 229652 155984
rect 145064 155944 229652 155972
rect 145064 155932 145070 155944
rect 229646 155932 229652 155944
rect 229704 155932 229710 155984
rect 66806 155864 66812 155916
rect 66864 155904 66870 155916
rect 82814 155904 82820 155916
rect 66864 155876 82820 155904
rect 66864 155864 66870 155876
rect 82814 155864 82820 155876
rect 82872 155864 82878 155916
rect 89530 155864 89536 155916
rect 89588 155904 89594 155916
rect 186314 155904 186320 155916
rect 89588 155876 186320 155904
rect 89588 155864 89594 155876
rect 186314 155864 186320 155876
rect 186372 155864 186378 155916
rect 186406 155864 186412 155916
rect 186464 155904 186470 155916
rect 192846 155904 192852 155916
rect 186464 155876 192852 155904
rect 186464 155864 186470 155876
rect 192846 155864 192852 155876
rect 192904 155864 192910 155916
rect 192938 155864 192944 155916
rect 192996 155904 193002 155916
rect 266262 155904 266268 155916
rect 192996 155876 266268 155904
rect 192996 155864 193002 155876
rect 266262 155864 266268 155876
rect 266320 155864 266326 155916
rect 296438 155864 296444 155916
rect 296496 155904 296502 155916
rect 345198 155904 345204 155916
rect 296496 155876 345204 155904
rect 296496 155864 296502 155876
rect 345198 155864 345204 155876
rect 345256 155864 345262 155916
rect 60090 155796 60096 155848
rect 60148 155836 60154 155848
rect 79318 155836 79324 155848
rect 60148 155808 79324 155836
rect 60148 155796 60154 155808
rect 79318 155796 79324 155808
rect 79376 155796 79382 155848
rect 88702 155796 88708 155848
rect 88760 155836 88766 155848
rect 186866 155836 186872 155848
rect 88760 155808 186872 155836
rect 88760 155796 88766 155808
rect 186866 155796 186872 155808
rect 186924 155796 186930 155848
rect 189626 155796 189632 155848
rect 189684 155836 189690 155848
rect 263778 155836 263784 155848
rect 189684 155808 263784 155836
rect 189684 155796 189690 155808
rect 263778 155796 263784 155808
rect 263836 155796 263842 155848
rect 293034 155796 293040 155848
rect 293092 155836 293098 155848
rect 342346 155836 342352 155848
rect 293092 155808 342352 155836
rect 293092 155796 293098 155808
rect 342346 155796 342352 155808
rect 342404 155796 342410 155848
rect 12158 155728 12164 155780
rect 12216 155768 12222 155780
rect 109126 155768 109132 155780
rect 12216 155740 109132 155768
rect 12216 155728 12222 155740
rect 109126 155728 109132 155740
rect 109184 155728 109190 155780
rect 112254 155728 112260 155780
rect 112312 155768 112318 155780
rect 204622 155768 204628 155780
rect 112312 155740 204628 155768
rect 112312 155728 112318 155740
rect 204622 155728 204628 155740
rect 204680 155728 204686 155780
rect 206462 155728 206468 155780
rect 206520 155768 206526 155780
rect 276106 155768 276112 155780
rect 206520 155740 276112 155768
rect 206520 155728 206526 155740
rect 276106 155728 276112 155740
rect 276164 155728 276170 155780
rect 289722 155728 289728 155780
rect 289780 155768 289786 155780
rect 339586 155768 339592 155780
rect 289780 155740 339592 155768
rect 289780 155728 289786 155740
rect 339586 155728 339592 155740
rect 339644 155728 339650 155780
rect 46566 155660 46572 155712
rect 46624 155700 46630 155712
rect 75454 155700 75460 155712
rect 46624 155672 75460 155700
rect 46624 155660 46630 155672
rect 75454 155660 75460 155672
rect 75512 155660 75518 155712
rect 81894 155660 81900 155712
rect 81952 155700 81958 155712
rect 180978 155700 180984 155712
rect 81952 155672 180984 155700
rect 81952 155660 81958 155672
rect 180978 155660 180984 155672
rect 181036 155660 181042 155712
rect 186222 155660 186228 155712
rect 186280 155700 186286 155712
rect 260834 155700 260840 155712
rect 186280 155672 260840 155700
rect 186280 155660 186286 155672
rect 260834 155660 260840 155672
rect 260892 155660 260898 155712
rect 270310 155660 270316 155712
rect 270368 155700 270374 155712
rect 325326 155700 325332 155712
rect 270368 155672 325332 155700
rect 270368 155660 270374 155672
rect 325326 155660 325332 155672
rect 325384 155660 325390 155712
rect 344370 155660 344376 155712
rect 344428 155700 344434 155712
rect 381814 155700 381820 155712
rect 344428 155672 381820 155700
rect 344428 155660 344434 155672
rect 381814 155660 381820 155672
rect 381872 155660 381878 155712
rect 53374 155592 53380 155644
rect 53432 155632 53438 155644
rect 67082 155632 67088 155644
rect 53432 155604 67088 155632
rect 53432 155592 53438 155604
rect 67082 155592 67088 155604
rect 67140 155592 67146 155644
rect 71866 155592 71872 155644
rect 71924 155632 71930 155644
rect 172698 155632 172704 155644
rect 71924 155604 172704 155632
rect 71924 155592 71930 155604
rect 172698 155592 172704 155604
rect 172756 155592 172762 155644
rect 176286 155592 176292 155644
rect 176344 155632 176350 155644
rect 253382 155632 253388 155644
rect 176344 155604 253388 155632
rect 176344 155592 176350 155604
rect 253382 155592 253388 155604
rect 253440 155592 253446 155644
rect 266998 155592 267004 155644
rect 267056 155632 267062 155644
rect 321738 155632 321744 155644
rect 267056 155604 321744 155632
rect 267056 155592 267062 155604
rect 321738 155592 321744 155604
rect 321796 155592 321802 155644
rect 340966 155592 340972 155644
rect 341024 155632 341030 155644
rect 378134 155632 378140 155644
rect 341024 155604 378140 155632
rect 341024 155592 341030 155604
rect 378134 155592 378140 155604
rect 378192 155592 378198 155644
rect 39850 155524 39856 155576
rect 39908 155564 39914 155576
rect 68830 155564 68836 155576
rect 39908 155536 68836 155564
rect 39908 155524 39914 155536
rect 68830 155524 68836 155536
rect 68888 155524 68894 155576
rect 75178 155524 75184 155576
rect 75236 155564 75242 155576
rect 176378 155564 176384 155576
rect 75236 155536 176384 155564
rect 75236 155524 75242 155536
rect 176378 155524 176384 155536
rect 176436 155524 176442 155576
rect 179506 155524 179512 155576
rect 179564 155564 179570 155576
rect 255774 155564 255780 155576
rect 179564 155536 255780 155564
rect 179564 155524 179570 155536
rect 255774 155524 255780 155536
rect 255832 155524 255838 155576
rect 263594 155524 263600 155576
rect 263652 155564 263658 155576
rect 320174 155564 320180 155576
rect 263652 155536 320180 155564
rect 263652 155524 263658 155536
rect 320174 155524 320180 155536
rect 320232 155524 320238 155576
rect 337654 155524 337660 155576
rect 337712 155564 337718 155576
rect 375558 155564 375564 155576
rect 337712 155536 375564 155564
rect 337712 155524 337718 155536
rect 375558 155524 375564 155536
rect 375616 155524 375622 155576
rect 65150 155456 65156 155508
rect 65208 155496 65214 155508
rect 168650 155496 168656 155508
rect 65208 155468 168656 155496
rect 65208 155456 65214 155468
rect 168650 155456 168656 155468
rect 168708 155456 168714 155508
rect 169386 155456 169392 155508
rect 169444 155496 169450 155508
rect 248230 155496 248236 155508
rect 169444 155468 248236 155496
rect 169444 155456 169450 155468
rect 248230 155456 248236 155468
rect 248288 155456 248294 155508
rect 260282 155456 260288 155508
rect 260340 155496 260346 155508
rect 317598 155496 317604 155508
rect 260340 155468 317604 155496
rect 260340 155456 260346 155468
rect 317598 155456 317604 155468
rect 317656 155456 317662 155508
rect 333422 155456 333428 155508
rect 333480 155496 333486 155508
rect 373442 155496 373448 155508
rect 333480 155468 373448 155496
rect 333480 155456 333486 155468
rect 373442 155456 373448 155468
rect 373500 155456 373506 155508
rect 8754 155388 8760 155440
rect 8812 155428 8818 155440
rect 125686 155428 125692 155440
rect 8812 155400 125692 155428
rect 8812 155388 8818 155400
rect 125686 155388 125692 155400
rect 125744 155388 125750 155440
rect 145834 155388 145840 155440
rect 145892 155428 145898 155440
rect 229186 155428 229192 155440
rect 145892 155400 229192 155428
rect 145892 155388 145898 155400
rect 229186 155388 229192 155400
rect 229244 155388 229250 155440
rect 253566 155388 253572 155440
rect 253624 155428 253630 155440
rect 312446 155428 312452 155440
rect 253624 155400 312452 155428
rect 253624 155388 253630 155400
rect 312446 155388 312452 155400
rect 312504 155388 312510 155440
rect 330110 155388 330116 155440
rect 330168 155428 330174 155440
rect 370866 155428 370872 155440
rect 330168 155400 370872 155428
rect 330168 155388 330174 155400
rect 370866 155388 370872 155400
rect 370924 155388 370930 155440
rect 7926 155320 7932 155372
rect 7984 155360 7990 155372
rect 124674 155360 124680 155372
rect 7984 155332 124680 155360
rect 7984 155320 7990 155332
rect 124674 155320 124680 155332
rect 124732 155320 124738 155372
rect 142522 155320 142528 155372
rect 142580 155360 142586 155372
rect 227806 155360 227812 155372
rect 142580 155332 227812 155360
rect 142580 155320 142586 155332
rect 227806 155320 227812 155332
rect 227864 155320 227870 155372
rect 250162 155320 250168 155372
rect 250220 155360 250226 155372
rect 309870 155360 309876 155372
rect 250220 155332 309876 155360
rect 250220 155320 250226 155332
rect 309870 155320 309876 155332
rect 309928 155320 309934 155372
rect 319990 155320 319996 155372
rect 320048 155360 320054 155372
rect 363230 155360 363236 155372
rect 320048 155332 363236 155360
rect 320048 155320 320054 155332
rect 363230 155320 363236 155332
rect 363288 155320 363294 155372
rect 4522 155252 4528 155304
rect 4580 155292 4586 155304
rect 122006 155292 122012 155304
rect 4580 155264 122012 155292
rect 4580 155252 4586 155264
rect 122006 155252 122012 155264
rect 122064 155252 122070 155304
rect 125778 155252 125784 155304
rect 125836 155292 125842 155304
rect 214834 155292 214840 155304
rect 125836 155264 214840 155292
rect 125836 155252 125842 155264
rect 214834 155252 214840 155264
rect 214892 155252 214898 155304
rect 240042 155252 240048 155304
rect 240100 155292 240106 155304
rect 302326 155292 302332 155304
rect 240100 155264 302332 155292
rect 240100 155252 240106 155264
rect 302326 155252 302332 155264
rect 302384 155252 302390 155304
rect 306558 155252 306564 155304
rect 306616 155292 306622 155304
rect 352466 155292 352472 155304
rect 306616 155264 352472 155292
rect 306616 155252 306622 155264
rect 352466 155252 352472 155264
rect 352524 155252 352530 155304
rect 373810 155252 373816 155304
rect 373868 155292 373874 155304
rect 404078 155292 404084 155304
rect 373868 155264 404084 155292
rect 373868 155252 373874 155264
rect 404078 155252 404084 155264
rect 404136 155252 404142 155304
rect 5350 155184 5356 155236
rect 5408 155224 5414 155236
rect 123018 155224 123024 155236
rect 5408 155196 123024 155224
rect 5408 155184 5414 155196
rect 123018 155184 123024 155196
rect 123076 155184 123082 155236
rect 128998 155184 129004 155236
rect 129056 155224 129062 155236
rect 217410 155224 217416 155236
rect 129056 155196 217416 155224
rect 129056 155184 129062 155196
rect 217410 155184 217416 155196
rect 217468 155184 217474 155236
rect 233326 155184 233332 155236
rect 233384 155224 233390 155236
rect 297082 155224 297088 155236
rect 233384 155196 297088 155224
rect 233384 155184 233390 155196
rect 297082 155184 297088 155196
rect 297140 155184 297146 155236
rect 299750 155184 299756 155236
rect 299808 155224 299814 155236
rect 347866 155224 347872 155236
rect 299808 155196 347872 155224
rect 299808 155184 299814 155196
rect 347866 155184 347872 155196
rect 347924 155184 347930 155236
rect 370406 155184 370412 155236
rect 370464 155224 370470 155236
rect 401686 155224 401692 155236
rect 370464 155196 401692 155224
rect 370464 155184 370470 155196
rect 401686 155184 401692 155196
rect 401744 155184 401750 155236
rect 92014 155116 92020 155168
rect 92072 155156 92078 155168
rect 189166 155156 189172 155168
rect 92072 155128 189172 155156
rect 92072 155116 92078 155128
rect 189166 155116 189172 155128
rect 189224 155116 189230 155168
rect 192846 155116 192852 155168
rect 192904 155156 192910 155168
rect 194318 155156 194324 155168
rect 192904 155128 194324 155156
rect 192904 155116 192910 155128
rect 194318 155116 194324 155128
rect 194376 155116 194382 155168
rect 196342 155116 196348 155168
rect 196400 155156 196406 155168
rect 268838 155156 268844 155168
rect 196400 155128 268844 155156
rect 196400 155116 196406 155128
rect 268838 155116 268844 155128
rect 268896 155116 268902 155168
rect 303154 155116 303160 155168
rect 303212 155156 303218 155168
rect 350350 155156 350356 155168
rect 303212 155128 350356 155156
rect 303212 155116 303218 155128
rect 350350 155116 350356 155128
rect 350408 155116 350414 155168
rect 95418 155048 95424 155100
rect 95476 155088 95482 155100
rect 95476 155060 186452 155088
rect 95476 155048 95482 155060
rect 98730 154980 98736 155032
rect 98788 155020 98794 155032
rect 186314 155020 186320 155032
rect 98788 154992 186320 155020
rect 98788 154980 98794 154992
rect 186314 154980 186320 154992
rect 186372 154980 186378 155032
rect 186424 155020 186452 155060
rect 186774 155048 186780 155100
rect 186832 155088 186838 155100
rect 186832 155060 195974 155088
rect 186832 155048 186838 155060
rect 191742 155020 191748 155032
rect 186424 154992 191748 155020
rect 191742 154980 191748 154992
rect 191800 154980 191806 155032
rect 195946 155020 195974 155060
rect 199654 155048 199660 155100
rect 199712 155088 199718 155100
rect 271414 155088 271420 155100
rect 199712 155060 271420 155088
rect 199712 155048 199718 155060
rect 271414 155048 271420 155060
rect 271472 155048 271478 155100
rect 200114 155020 200120 155032
rect 195946 154992 200120 155020
rect 200114 154980 200120 154992
rect 200172 154980 200178 155032
rect 207014 154980 207020 155032
rect 207072 155020 207078 155032
rect 269482 155020 269488 155032
rect 207072 154992 269488 155020
rect 207072 154980 207078 154992
rect 269482 154980 269488 154992
rect 269540 154980 269546 155032
rect 15470 154912 15476 154964
rect 15528 154952 15534 154964
rect 109034 154952 109040 154964
rect 15528 154924 109040 154952
rect 15528 154912 15534 154924
rect 109034 154912 109040 154924
rect 109092 154912 109098 154964
rect 122282 154912 122288 154964
rect 122340 154952 122346 154964
rect 211246 154952 211252 154964
rect 122340 154924 211252 154952
rect 122340 154912 122346 154924
rect 211246 154912 211252 154924
rect 211304 154912 211310 154964
rect 214558 154912 214564 154964
rect 214616 154952 214622 154964
rect 261386 154952 261392 154964
rect 214616 154924 261392 154952
rect 214616 154912 214622 154924
rect 261386 154912 261392 154924
rect 261444 154912 261450 154964
rect 106366 154844 106372 154896
rect 106424 154884 106430 154896
rect 186406 154884 186412 154896
rect 106424 154856 186412 154884
rect 106424 154844 106430 154856
rect 186406 154844 186412 154856
rect 186464 154844 186470 154896
rect 186682 154844 186688 154896
rect 186740 154884 186746 154896
rect 245838 154884 245844 154896
rect 186740 154856 245844 154884
rect 186740 154844 186746 154856
rect 245838 154844 245844 154856
rect 245896 154844 245902 154896
rect 110506 154776 110512 154828
rect 110564 154816 110570 154828
rect 139302 154816 139308 154828
rect 110564 154788 139308 154816
rect 110564 154776 110570 154788
rect 139302 154776 139308 154788
rect 139360 154776 139366 154828
rect 149238 154776 149244 154828
rect 149296 154816 149302 154828
rect 232866 154816 232872 154828
rect 149296 154788 232872 154816
rect 149296 154776 149302 154788
rect 232866 154776 232872 154788
rect 232924 154776 232930 154828
rect 109218 154708 109224 154760
rect 109276 154748 109282 154760
rect 133046 154748 133052 154760
rect 109276 154720 133052 154748
rect 109276 154708 109282 154720
rect 133046 154708 133052 154720
rect 133104 154708 133110 154760
rect 151906 154708 151912 154760
rect 151964 154748 151970 154760
rect 153102 154748 153108 154760
rect 151964 154720 153108 154748
rect 151964 154708 151970 154720
rect 153102 154708 153108 154720
rect 153160 154708 153166 154760
rect 155954 154708 155960 154760
rect 156012 154748 156018 154760
rect 238018 154748 238024 154760
rect 156012 154720 238024 154748
rect 156012 154708 156018 154720
rect 238018 154708 238024 154720
rect 238076 154708 238082 154760
rect 280264 154720 283788 154748
rect 159358 154640 159364 154692
rect 159416 154680 159422 154692
rect 240594 154680 240600 154692
rect 159416 154652 240600 154680
rect 159416 154640 159422 154652
rect 240594 154640 240600 154652
rect 240652 154640 240658 154692
rect 118602 154572 118608 154624
rect 118660 154612 118666 154624
rect 119982 154612 119988 154624
rect 118660 154584 119988 154612
rect 118660 154572 118666 154584
rect 119982 154572 119988 154584
rect 120040 154572 120046 154624
rect 137094 154572 137100 154624
rect 137152 154612 137158 154624
rect 138014 154612 138020 154624
rect 137152 154584 138020 154612
rect 137152 154572 137158 154584
rect 138014 154572 138020 154584
rect 138072 154572 138078 154624
rect 152642 154612 152648 154624
rect 152384 154584 152648 154612
rect 48314 154504 48320 154556
rect 48372 154544 48378 154556
rect 152384 154544 152412 154584
rect 152642 154572 152648 154584
rect 152700 154572 152706 154624
rect 162670 154572 162676 154624
rect 162728 154612 162734 154624
rect 243078 154612 243084 154624
rect 162728 154584 243084 154612
rect 162728 154572 162734 154584
rect 243078 154572 243084 154584
rect 243136 154572 243142 154624
rect 48372 154516 152412 154544
rect 48372 154504 48378 154516
rect 152458 154504 152464 154556
rect 152516 154544 152522 154556
rect 202690 154544 202696 154556
rect 152516 154516 202696 154544
rect 152516 154504 152522 154516
rect 202690 154504 202696 154516
rect 202748 154504 202754 154556
rect 218330 154504 218336 154556
rect 218388 154544 218394 154556
rect 280264 154544 280292 154720
rect 283650 154544 283656 154556
rect 218388 154516 280292 154544
rect 283024 154516 283656 154544
rect 218388 154504 218394 154516
rect 44174 154436 44180 154488
rect 44232 154476 44238 154488
rect 142890 154476 142896 154488
rect 44232 154448 142896 154476
rect 44232 154436 44238 154448
rect 142890 154436 142896 154448
rect 142948 154436 142954 154488
rect 142982 154436 142988 154488
rect 143040 154476 143046 154488
rect 188246 154476 188252 154488
rect 143040 154448 188252 154476
rect 143040 154436 143046 154448
rect 188246 154436 188252 154448
rect 188304 154436 188310 154488
rect 189810 154476 189816 154488
rect 188356 154448 189816 154476
rect 114462 154368 114468 154420
rect 114520 154408 114526 154420
rect 118602 154408 118608 154420
rect 114520 154380 118608 154408
rect 114520 154368 114526 154380
rect 118602 154368 118608 154380
rect 118660 154368 118666 154420
rect 118694 154368 118700 154420
rect 118752 154408 118758 154420
rect 119890 154408 119896 154420
rect 118752 154380 119896 154408
rect 118752 154368 118758 154380
rect 119890 154368 119896 154380
rect 119948 154368 119954 154420
rect 119982 154368 119988 154420
rect 120040 154408 120046 154420
rect 188356 154408 188384 154448
rect 189810 154436 189816 154448
rect 189868 154436 189874 154488
rect 191006 154436 191012 154488
rect 191064 154476 191070 154488
rect 191064 154448 198412 154476
rect 191064 154436 191070 154448
rect 120040 154380 188384 154408
rect 120040 154368 120046 154380
rect 188430 154368 188436 154420
rect 188488 154408 188494 154420
rect 197538 154408 197544 154420
rect 188488 154380 197544 154408
rect 188488 154368 188494 154380
rect 197538 154368 197544 154380
rect 197596 154368 197602 154420
rect 198384 154408 198412 154448
rect 198458 154436 198464 154488
rect 198516 154476 198522 154488
rect 210418 154476 210424 154488
rect 198516 154448 210424 154476
rect 198516 154436 198522 154448
rect 210418 154436 210424 154448
rect 210476 154436 210482 154488
rect 215294 154436 215300 154488
rect 215352 154476 215358 154488
rect 283024 154476 283052 154516
rect 283650 154504 283656 154516
rect 283708 154504 283714 154556
rect 283760 154544 283788 154720
rect 285582 154544 285588 154556
rect 283760 154516 285588 154544
rect 285582 154504 285588 154516
rect 285640 154504 285646 154556
rect 285674 154504 285680 154556
rect 285732 154544 285738 154556
rect 337470 154544 337476 154556
rect 285732 154516 337476 154544
rect 285732 154504 285738 154516
rect 337470 154504 337476 154516
rect 337528 154504 337534 154556
rect 353662 154504 353668 154556
rect 353720 154544 353726 154556
rect 388898 154544 388904 154556
rect 353720 154516 388904 154544
rect 353720 154504 353726 154516
rect 388898 154504 388904 154516
rect 388956 154504 388962 154556
rect 215352 154448 283052 154476
rect 215352 154436 215358 154448
rect 283282 154436 283288 154488
rect 283340 154476 283346 154488
rect 334894 154476 334900 154488
rect 283340 154448 334900 154476
rect 283340 154436 283346 154448
rect 334894 154436 334900 154448
rect 334952 154436 334958 154488
rect 349522 154436 349528 154488
rect 349580 154476 349586 154488
rect 386230 154476 386236 154488
rect 349580 154448 386236 154476
rect 349580 154436 349586 154448
rect 386230 154436 386236 154448
rect 386288 154436 386294 154488
rect 390646 154436 390652 154488
rect 390704 154476 390710 154488
rect 417142 154476 417148 154488
rect 390704 154448 417148 154476
rect 390704 154436 390710 154448
rect 417142 154436 417148 154448
rect 417200 154436 417206 154488
rect 202046 154408 202052 154420
rect 198384 154380 202052 154408
rect 202046 154368 202052 154380
rect 202104 154368 202110 154420
rect 205082 154368 205088 154420
rect 205140 154408 205146 154420
rect 275830 154408 275836 154420
rect 205140 154380 275836 154408
rect 205140 154368 205146 154380
rect 275830 154368 275836 154380
rect 275888 154368 275894 154420
rect 276198 154368 276204 154420
rect 276256 154408 276262 154420
rect 329926 154408 329932 154420
rect 276256 154380 329932 154408
rect 276256 154368 276262 154380
rect 329926 154368 329932 154380
rect 329984 154368 329990 154420
rect 346394 154368 346400 154420
rect 346452 154408 346458 154420
rect 383746 154408 383752 154420
rect 346452 154380 383752 154408
rect 346452 154368 346458 154380
rect 383746 154368 383752 154380
rect 383804 154368 383810 154420
rect 397362 154368 397368 154420
rect 397420 154408 397426 154420
rect 422294 154408 422300 154420
rect 397420 154380 422300 154408
rect 397420 154368 397426 154380
rect 422294 154368 422300 154380
rect 422352 154368 422358 154420
rect 34514 154300 34520 154352
rect 34572 154340 34578 154352
rect 142614 154340 142620 154352
rect 34572 154312 142620 154340
rect 34572 154300 34578 154312
rect 142614 154300 142620 154312
rect 142672 154300 142678 154352
rect 142706 154300 142712 154352
rect 142764 154340 142770 154352
rect 205266 154340 205272 154352
rect 142764 154312 205272 154340
rect 142764 154300 142770 154312
rect 205266 154300 205272 154312
rect 205324 154300 205330 154352
rect 208394 154300 208400 154352
rect 208452 154340 208458 154352
rect 278406 154340 278412 154352
rect 208452 154312 278412 154340
rect 208452 154300 208458 154312
rect 278406 154300 278412 154312
rect 278464 154300 278470 154352
rect 278866 154300 278872 154352
rect 278924 154340 278930 154352
rect 332410 154340 332416 154352
rect 278924 154312 332416 154340
rect 278924 154300 278930 154312
rect 332410 154300 332416 154312
rect 332468 154300 332474 154352
rect 342806 154300 342812 154352
rect 342864 154340 342870 154352
rect 381170 154340 381176 154352
rect 342864 154312 381176 154340
rect 342864 154300 342870 154312
rect 381170 154300 381176 154312
rect 381228 154300 381234 154352
rect 393314 154300 393320 154352
rect 393372 154340 393378 154352
rect 419718 154340 419724 154352
rect 393372 154312 419724 154340
rect 393372 154300 393378 154312
rect 419718 154300 419724 154312
rect 419776 154300 419782 154352
rect 434714 154300 434720 154352
rect 434772 154340 434778 154352
rect 444282 154340 444288 154352
rect 434772 154312 444288 154340
rect 434772 154300 434778 154312
rect 444282 154300 444288 154312
rect 444340 154300 444346 154352
rect 37918 154232 37924 154284
rect 37976 154272 37982 154284
rect 37976 154244 142660 154272
rect 37976 154232 37982 154244
rect 27246 154164 27252 154216
rect 27304 154204 27310 154216
rect 136910 154204 136916 154216
rect 27304 154176 136916 154204
rect 27304 154164 27310 154176
rect 136910 154164 136916 154176
rect 136968 154164 136974 154216
rect 142632 154204 142660 154244
rect 143074 154232 143080 154284
rect 143132 154272 143138 154284
rect 152458 154272 152464 154284
rect 143132 154244 152464 154272
rect 143132 154232 143138 154244
rect 152458 154232 152464 154244
rect 152516 154232 152522 154284
rect 152642 154232 152648 154284
rect 152700 154272 152706 154284
rect 155770 154272 155776 154284
rect 152700 154244 155776 154272
rect 152700 154232 152706 154244
rect 155770 154232 155776 154244
rect 155828 154232 155834 154284
rect 161474 154232 161480 154284
rect 161532 154272 161538 154284
rect 166074 154272 166080 154284
rect 161532 154244 166080 154272
rect 161532 154232 161538 154244
rect 166074 154232 166080 154244
rect 166132 154232 166138 154284
rect 176654 154232 176660 154284
rect 176712 154272 176718 154284
rect 179690 154272 179696 154284
rect 176712 154244 179696 154272
rect 176712 154232 176718 154244
rect 179690 154232 179696 154244
rect 179748 154232 179754 154284
rect 182174 154232 182180 154284
rect 182232 154272 182238 154284
rect 258534 154272 258540 154284
rect 182232 154244 258540 154272
rect 182232 154232 182238 154244
rect 258534 154232 258540 154244
rect 258592 154232 258598 154284
rect 262214 154232 262220 154284
rect 262272 154272 262278 154284
rect 319530 154272 319536 154284
rect 262272 154244 319536 154272
rect 262272 154232 262278 154244
rect 319530 154232 319536 154244
rect 319588 154232 319594 154284
rect 339494 154232 339500 154284
rect 339552 154272 339558 154284
rect 378594 154272 378600 154284
rect 339552 154244 378600 154272
rect 339552 154232 339558 154244
rect 378594 154232 378600 154244
rect 378652 154232 378658 154284
rect 386506 154232 386512 154284
rect 386564 154272 386570 154284
rect 414566 154272 414572 154284
rect 386564 154244 414572 154272
rect 386564 154232 386570 154244
rect 414566 154232 414572 154244
rect 414624 154232 414630 154284
rect 137112 154176 142568 154204
rect 142632 154176 142752 154204
rect 23474 154096 23480 154148
rect 23532 154136 23538 154148
rect 137002 154136 137008 154148
rect 23532 154108 137008 154136
rect 23532 154096 23538 154108
rect 137002 154096 137008 154108
rect 137060 154096 137066 154148
rect 13814 154028 13820 154080
rect 13872 154068 13878 154080
rect 129274 154068 129280 154080
rect 13872 154040 129280 154068
rect 13872 154028 13878 154040
rect 129274 154028 129280 154040
rect 129332 154028 129338 154080
rect 137112 154068 137140 154176
rect 142430 154136 142436 154148
rect 129476 154040 137140 154068
rect 137204 154108 142436 154136
rect 9674 153960 9680 154012
rect 9732 154000 9738 154012
rect 126882 154000 126888 154012
rect 9732 153972 126888 154000
rect 9732 153960 9738 153972
rect 126882 153960 126888 153972
rect 126940 153960 126946 154012
rect 127618 153960 127624 154012
rect 127676 154000 127682 154012
rect 129366 154000 129372 154012
rect 127676 153972 129372 154000
rect 127676 153960 127682 153972
rect 129366 153960 129372 153972
rect 129424 153960 129430 154012
rect 7098 153892 7104 153944
rect 7156 153932 7162 153944
rect 124306 153932 124312 153944
rect 7156 153904 124312 153932
rect 7156 153892 7162 153904
rect 124306 153892 124312 153904
rect 124364 153892 124370 153944
rect 125502 153892 125508 153944
rect 125560 153932 125566 153944
rect 129476 153932 129504 154040
rect 129642 153960 129648 154012
rect 129700 154000 129706 154012
rect 137204 154000 137232 154108
rect 142430 154096 142436 154108
rect 142488 154096 142494 154148
rect 142540 154136 142568 154176
rect 142724 154136 142752 154176
rect 142890 154164 142896 154216
rect 142948 154204 142954 154216
rect 142948 154176 151952 154204
rect 142948 154164 142954 154176
rect 148134 154136 148140 154148
rect 142540 154108 142660 154136
rect 142724 154108 148140 154136
rect 137278 154028 137284 154080
rect 137336 154068 137342 154080
rect 139762 154068 139768 154080
rect 137336 154040 139768 154068
rect 137336 154028 137342 154040
rect 139762 154028 139768 154040
rect 139820 154028 139826 154080
rect 139854 154028 139860 154080
rect 139912 154068 139918 154080
rect 142522 154068 142528 154080
rect 139912 154040 142528 154068
rect 139912 154028 139918 154040
rect 142522 154028 142528 154040
rect 142580 154028 142586 154080
rect 142632 154068 142660 154108
rect 148134 154096 148140 154108
rect 148192 154096 148198 154148
rect 148318 154096 148324 154148
rect 148376 154136 148382 154148
rect 151924 154136 151952 154176
rect 152274 154164 152280 154216
rect 152332 154204 152338 154216
rect 163498 154204 163504 154216
rect 152332 154176 163504 154204
rect 152332 154164 152338 154176
rect 163498 154164 163504 154176
rect 163556 154164 163562 154216
rect 172514 154164 172520 154216
rect 172572 154204 172578 154216
rect 250806 154204 250812 154216
rect 172572 154176 250812 154204
rect 172572 154164 172578 154176
rect 250806 154164 250812 154176
rect 250864 154164 250870 154216
rect 255314 154164 255320 154216
rect 255372 154204 255378 154216
rect 314378 154204 314384 154216
rect 255372 154176 314384 154204
rect 255372 154164 255378 154176
rect 314378 154164 314384 154176
rect 314436 154164 314442 154216
rect 336826 154164 336832 154216
rect 336884 154204 336890 154216
rect 376018 154204 376024 154216
rect 336884 154176 376024 154204
rect 336884 154164 336890 154176
rect 376018 154164 376024 154176
rect 376076 154164 376082 154216
rect 383654 154164 383660 154216
rect 383712 154204 383718 154216
rect 411990 154204 411996 154216
rect 383712 154176 411996 154204
rect 383712 154164 383718 154176
rect 411990 154164 411996 154176
rect 412048 154164 412054 154216
rect 153194 154136 153200 154148
rect 148376 154108 150756 154136
rect 151924 154108 153200 154136
rect 148376 154096 148382 154108
rect 142982 154068 142988 154080
rect 142632 154040 142988 154068
rect 142982 154028 142988 154040
rect 143040 154028 143046 154080
rect 143092 154040 143304 154068
rect 143092 154000 143120 154040
rect 129700 153972 137232 154000
rect 137940 153972 143120 154000
rect 143276 154000 143304 154040
rect 143534 154028 143540 154080
rect 143592 154068 143598 154080
rect 150618 154068 150624 154080
rect 143592 154040 150624 154068
rect 143592 154028 143598 154040
rect 150618 154028 150624 154040
rect 150676 154028 150682 154080
rect 150728 154068 150756 154108
rect 153194 154096 153200 154108
rect 153252 154096 153258 154148
rect 153286 154096 153292 154148
rect 153344 154136 153350 154148
rect 158438 154136 158444 154148
rect 153344 154108 158444 154136
rect 153344 154096 153350 154108
rect 158438 154096 158444 154108
rect 158496 154096 158502 154148
rect 160186 154096 160192 154148
rect 160244 154136 160250 154148
rect 160244 154108 162900 154136
rect 160244 154096 160250 154108
rect 152182 154068 152188 154080
rect 150728 154040 152188 154068
rect 152182 154028 152188 154040
rect 152240 154028 152246 154080
rect 152366 154028 152372 154080
rect 152424 154068 152430 154080
rect 161566 154068 161572 154080
rect 152424 154040 161572 154068
rect 152424 154028 152430 154040
rect 161566 154028 161572 154040
rect 161624 154028 161630 154080
rect 162872 154068 162900 154108
rect 165614 154096 165620 154148
rect 165672 154136 165678 154148
rect 245654 154136 245660 154148
rect 165672 154108 245660 154136
rect 165672 154096 165678 154108
rect 245654 154096 245660 154108
rect 245712 154096 245718 154148
rect 245930 154096 245936 154148
rect 245988 154136 245994 154148
rect 306650 154136 306656 154148
rect 245988 154108 306656 154136
rect 245988 154096 245994 154108
rect 306650 154096 306656 154108
rect 306708 154096 306714 154148
rect 326706 154096 326712 154148
rect 326764 154136 326770 154148
rect 368290 154136 368296 154148
rect 326764 154108 368296 154136
rect 326764 154096 326770 154108
rect 368290 154096 368296 154108
rect 368348 154096 368354 154148
rect 376846 154096 376852 154148
rect 376904 154136 376910 154148
rect 406838 154136 406844 154148
rect 376904 154108 406844 154136
rect 376904 154096 376910 154108
rect 406838 154096 406844 154108
rect 406896 154096 406902 154148
rect 241238 154068 241244 154080
rect 162872 154040 241244 154068
rect 241238 154028 241244 154040
rect 241296 154028 241302 154080
rect 248598 154028 248604 154080
rect 248656 154068 248662 154080
rect 309226 154068 309232 154080
rect 248656 154040 309232 154068
rect 248656 154028 248662 154040
rect 309226 154028 309232 154040
rect 309284 154028 309290 154080
rect 323302 154028 323308 154080
rect 323360 154068 323366 154080
rect 365806 154068 365812 154080
rect 323360 154040 365812 154068
rect 323360 154028 323366 154040
rect 365806 154028 365812 154040
rect 365864 154028 365870 154080
rect 380158 154028 380164 154080
rect 380216 154068 380222 154080
rect 409414 154068 409420 154080
rect 380216 154040 409420 154068
rect 380216 154028 380222 154040
rect 409414 154028 409420 154040
rect 409472 154028 409478 154080
rect 219894 154000 219900 154012
rect 143276 153972 219900 154000
rect 129700 153960 129706 153972
rect 125560 153904 129504 153932
rect 125560 153892 125566 153904
rect 132402 153892 132408 153944
rect 132460 153932 132466 153944
rect 137940 153932 137968 153972
rect 219894 153960 219900 153972
rect 219952 153960 219958 154012
rect 222378 153960 222384 154012
rect 222436 154000 222442 154012
rect 288710 154000 288716 154012
rect 222436 153972 288716 154000
rect 222436 153960 222442 153972
rect 288710 153960 288716 153972
rect 288768 153960 288774 154012
rect 313274 153960 313280 154012
rect 313332 154000 313338 154012
rect 357894 154000 357900 154012
rect 313332 153972 357900 154000
rect 313332 153960 313338 153972
rect 357894 153960 357900 153972
rect 357952 153960 357958 154012
rect 367094 153960 367100 154012
rect 367152 154000 367158 154012
rect 399110 154000 399116 154012
rect 367152 153972 399116 154000
rect 367152 153960 367158 153972
rect 399110 153960 399116 153972
rect 399168 153960 399174 154012
rect 132460 153904 137968 153932
rect 132460 153892 132466 153904
rect 138014 153892 138020 153944
rect 138072 153932 138078 153944
rect 143074 153932 143080 153944
rect 138072 153904 143080 153932
rect 138072 153892 138078 153904
rect 143074 153892 143080 153904
rect 143132 153892 143138 153944
rect 143258 153892 143264 153944
rect 143316 153932 143322 153944
rect 145558 153932 145564 153944
rect 143316 153904 145564 153932
rect 143316 153892 143322 153904
rect 145558 153892 145564 153904
rect 145616 153892 145622 153944
rect 223206 153932 223212 153944
rect 145668 153904 223212 153932
rect 474 153824 480 153876
rect 532 153864 538 153876
rect 119798 153864 119804 153876
rect 532 153836 119804 153864
rect 532 153824 538 153836
rect 119798 153824 119804 153836
rect 119856 153824 119862 153876
rect 119890 153824 119896 153876
rect 119948 153864 119954 153876
rect 142798 153864 142804 153876
rect 119948 153836 142804 153864
rect 119948 153824 119954 153836
rect 142798 153824 142804 153836
rect 142856 153824 142862 153876
rect 143350 153824 143356 153876
rect 143408 153864 143414 153876
rect 145668 153864 145696 153904
rect 223206 153892 223212 153904
rect 223264 153892 223270 153944
rect 225230 153892 225236 153944
rect 225288 153932 225294 153944
rect 291286 153932 291292 153944
rect 225288 153904 291292 153932
rect 225288 153892 225294 153904
rect 291286 153892 291292 153904
rect 291344 153892 291350 153944
rect 316034 153892 316040 153944
rect 316092 153932 316098 153944
rect 360654 153932 360660 153944
rect 316092 153904 360660 153932
rect 316092 153892 316098 153904
rect 360654 153892 360660 153904
rect 360712 153892 360718 153944
rect 363046 153892 363052 153944
rect 363104 153932 363110 153944
rect 396534 153932 396540 153944
rect 363104 153904 396540 153932
rect 363104 153892 363110 153904
rect 396534 153892 396540 153904
rect 396592 153892 396598 153944
rect 401594 153892 401600 153944
rect 401652 153932 401658 153944
rect 425514 153932 425520 153944
rect 401652 153904 425520 153932
rect 401652 153892 401658 153904
rect 425514 153892 425520 153904
rect 425572 153892 425578 153944
rect 143408 153836 145696 153864
rect 143408 153824 143414 153836
rect 147398 153824 147404 153876
rect 147456 153864 147462 153876
rect 152366 153864 152372 153876
rect 147456 153836 152372 153864
rect 147456 153824 147462 153836
rect 152366 153824 152372 153836
rect 152424 153824 152430 153876
rect 158346 153864 158352 153876
rect 152476 153836 158352 153864
rect 51074 153756 51080 153808
rect 51132 153796 51138 153808
rect 152476 153796 152504 153836
rect 158346 153824 158352 153836
rect 158404 153824 158410 153876
rect 158438 153824 158444 153876
rect 158496 153864 158502 153876
rect 235442 153864 235448 153876
rect 158496 153836 235448 153864
rect 158496 153824 158502 153836
rect 235442 153824 235448 153836
rect 235500 153824 235506 153876
rect 241882 153824 241888 153876
rect 241940 153864 241946 153876
rect 304074 153864 304080 153876
rect 241940 153836 304080 153864
rect 241940 153824 241946 153836
rect 304074 153824 304080 153836
rect 304132 153824 304138 153876
rect 309134 153824 309140 153876
rect 309192 153864 309198 153876
rect 355502 153864 355508 153876
rect 309192 153836 355508 153864
rect 309192 153824 309198 153836
rect 355502 153824 355508 153836
rect 355560 153824 355566 153876
rect 356238 153824 356244 153876
rect 356296 153864 356302 153876
rect 391474 153864 391480 153876
rect 356296 153836 391480 153864
rect 356296 153824 356302 153836
rect 391474 153824 391480 153836
rect 391532 153824 391538 153876
rect 397454 153824 397460 153876
rect 397512 153864 397518 153876
rect 422846 153864 422852 153876
rect 397512 153836 422852 153864
rect 397512 153824 397518 153836
rect 422846 153824 422852 153836
rect 422904 153824 422910 153876
rect 51132 153768 152504 153796
rect 51132 153756 51138 153768
rect 152642 153756 152648 153808
rect 152700 153796 152706 153808
rect 212902 153796 212908 153808
rect 152700 153768 212908 153796
rect 152700 153756 152706 153768
rect 212902 153756 212908 153768
rect 212960 153756 212966 153808
rect 231854 153756 231860 153808
rect 231912 153796 231918 153808
rect 296438 153796 296444 153808
rect 231912 153768 296444 153796
rect 231912 153756 231918 153768
rect 296438 153756 296444 153768
rect 296496 153756 296502 153808
rect 360378 153756 360384 153808
rect 360436 153796 360442 153808
rect 394050 153796 394056 153808
rect 360436 153768 394056 153796
rect 360436 153756 360442 153768
rect 394050 153756 394056 153768
rect 394108 153756 394114 153808
rect 61102 153688 61108 153740
rect 61160 153728 61166 153740
rect 161474 153728 161480 153740
rect 61160 153700 152596 153728
rect 61160 153688 61166 153700
rect 57974 153620 57980 153672
rect 58032 153660 58038 153672
rect 152274 153660 152280 153672
rect 58032 153632 152280 153660
rect 58032 153620 58038 153632
rect 152274 153620 152280 153632
rect 152332 153620 152338 153672
rect 152568 153660 152596 153700
rect 152752 153700 161480 153728
rect 152752 153660 152780 153700
rect 161474 153688 161480 153700
rect 161532 153688 161538 153740
rect 161566 153688 161572 153740
rect 161624 153728 161630 153740
rect 198458 153728 198464 153740
rect 161624 153700 198464 153728
rect 161624 153688 161630 153700
rect 198458 153688 198464 153700
rect 198516 153688 198522 153740
rect 198550 153688 198556 153740
rect 198608 153728 198614 153740
rect 209774 153728 209780 153740
rect 198608 153700 209780 153728
rect 198608 153688 198614 153700
rect 209774 153688 209780 153700
rect 209832 153688 209838 153740
rect 229094 153688 229100 153740
rect 229152 153728 229158 153740
rect 293862 153728 293868 153740
rect 229152 153700 293868 153728
rect 229152 153688 229158 153700
rect 293862 153688 293868 153700
rect 293920 153688 293926 153740
rect 152568 153632 152780 153660
rect 154482 153620 154488 153672
rect 154540 153660 154546 153672
rect 218054 153660 218060 153672
rect 154540 153632 218060 153660
rect 154540 153620 154546 153632
rect 218054 153620 218060 153632
rect 218112 153620 218118 153672
rect 235074 153620 235080 153672
rect 235132 153660 235138 153672
rect 299014 153660 299020 153672
rect 235132 153632 299020 153660
rect 235132 153620 235138 153632
rect 299014 153620 299020 153632
rect 299072 153620 299078 153672
rect 78674 153552 78680 153604
rect 78732 153592 78738 153604
rect 179598 153592 179604 153604
rect 78732 153564 179604 153592
rect 78732 153552 78738 153564
rect 179598 153552 179604 153564
rect 179656 153552 179662 153604
rect 179690 153552 179696 153604
rect 179748 153592 179754 153604
rect 230934 153592 230940 153604
rect 179748 153564 230940 153592
rect 179748 153552 179754 153564
rect 230934 153552 230940 153564
rect 230992 153552 230998 153604
rect 238846 153552 238852 153604
rect 238904 153592 238910 153604
rect 301590 153592 301596 153604
rect 238904 153564 301596 153592
rect 238904 153552 238910 153564
rect 301590 153552 301596 153564
rect 301648 153552 301654 153604
rect 102134 153484 102140 153536
rect 102192 153524 102198 153536
rect 196894 153524 196900 153536
rect 102192 153496 196900 153524
rect 102192 153484 102198 153496
rect 196894 153484 196900 153496
rect 196952 153484 196958 153536
rect 197262 153484 197268 153536
rect 197320 153524 197326 153536
rect 198642 153524 198648 153536
rect 197320 153496 198648 153524
rect 197320 153484 197326 153496
rect 198642 153484 198648 153496
rect 198700 153484 198706 153536
rect 198918 153484 198924 153536
rect 198976 153524 198982 153536
rect 248874 153524 248880 153536
rect 198976 153496 248880 153524
rect 198976 153484 198982 153496
rect 248874 153484 248880 153496
rect 248932 153484 248938 153536
rect 252646 153484 252652 153536
rect 252704 153524 252710 153536
rect 311802 153524 311808 153536
rect 252704 153496 311808 153524
rect 252704 153484 252710 153496
rect 311802 153484 311808 153496
rect 311860 153484 311866 153536
rect 104894 153416 104900 153468
rect 104952 153456 104958 153468
rect 199470 153456 199476 153468
rect 104952 153428 199476 153456
rect 104952 153416 104958 153428
rect 199470 153416 199476 153428
rect 199528 153416 199534 153468
rect 207842 153456 207848 153468
rect 200316 153428 207848 153456
rect 108298 153348 108304 153400
rect 108356 153388 108362 153400
rect 191006 153388 191012 153400
rect 108356 153360 191012 153388
rect 108356 153348 108362 153360
rect 191006 153348 191012 153360
rect 191064 153348 191070 153400
rect 191650 153348 191656 153400
rect 191708 153388 191714 153400
rect 200206 153388 200212 153400
rect 191708 153360 200212 153388
rect 191708 153348 191714 153360
rect 200206 153348 200212 153360
rect 200264 153348 200270 153400
rect 115934 153280 115940 153332
rect 115992 153320 115998 153332
rect 200316 153320 200344 153428
rect 207842 153416 207848 153428
rect 207900 153416 207906 153468
rect 207934 153416 207940 153468
rect 207992 153456 207998 153468
rect 259178 153456 259184 153468
rect 207992 153428 259184 153456
rect 207992 153416 207998 153428
rect 259178 153416 259184 153428
rect 259236 153416 259242 153468
rect 265434 153416 265440 153468
rect 265492 153456 265498 153468
rect 322198 153456 322204 153468
rect 265492 153428 322204 153456
rect 265492 153416 265498 153428
rect 322198 153416 322204 153428
rect 322256 153416 322262 153468
rect 243722 153388 243728 153400
rect 115992 153292 200344 153320
rect 200500 153360 243728 153388
rect 115992 153280 115998 153292
rect 41598 153212 41604 153264
rect 41656 153252 41662 153264
rect 138382 153252 138388 153264
rect 41656 153224 138388 153252
rect 41656 153212 41662 153224
rect 138382 153212 138388 153224
rect 138440 153212 138446 153264
rect 142798 153212 142804 153264
rect 142856 153252 142862 153264
rect 198550 153252 198556 153264
rect 142856 153224 198556 153252
rect 142856 153212 142862 153224
rect 198550 153212 198556 153224
rect 198608 153212 198614 153264
rect 198642 153212 198648 153264
rect 198700 153252 198706 153264
rect 200500 153252 200528 153360
rect 243722 153348 243728 153360
rect 243780 153348 243786 153400
rect 259454 153348 259460 153400
rect 259512 153388 259518 153400
rect 316954 153388 316960 153400
rect 259512 153360 316960 153388
rect 259512 153348 259518 153360
rect 316954 153348 316960 153360
rect 317012 153348 317018 153400
rect 200574 153280 200580 153332
rect 200632 153320 200638 153332
rect 238662 153320 238668 153332
rect 200632 153292 238668 153320
rect 200632 153280 200638 153292
rect 238662 153280 238668 153292
rect 238720 153280 238726 153332
rect 269206 153280 269212 153332
rect 269264 153320 269270 153332
rect 324682 153320 324688 153332
rect 269264 153292 324688 153320
rect 269264 153280 269270 153292
rect 324682 153280 324688 153292
rect 324740 153280 324746 153332
rect 198700 153224 200528 153252
rect 198700 153212 198706 153224
rect 201402 153212 201408 153264
rect 201460 153252 201466 153264
rect 207934 153252 207940 153264
rect 201460 153224 207940 153252
rect 201460 153212 201466 153224
rect 207934 153212 207940 153224
rect 207992 153212 207998 153264
rect 272886 153212 272892 153264
rect 272944 153252 272950 153264
rect 327258 153252 327264 153264
rect 272944 153224 327264 153252
rect 272944 153212 272950 153224
rect 327258 153212 327264 153224
rect 327316 153212 327322 153264
rect 113174 153144 113180 153196
rect 113232 153184 113238 153196
rect 205910 153184 205916 153196
rect 113232 153156 205916 153184
rect 113232 153144 113238 153156
rect 205910 153144 205916 153156
rect 205968 153144 205974 153196
rect 215386 153144 215392 153196
rect 215444 153184 215450 153196
rect 279694 153184 279700 153196
rect 215444 153156 279700 153184
rect 215444 153144 215450 153156
rect 279694 153144 279700 153156
rect 279752 153144 279758 153196
rect 285490 153144 285496 153196
rect 285548 153184 285554 153196
rect 336826 153184 336832 153196
rect 285548 153156 336832 153184
rect 285548 153144 285554 153156
rect 336826 153144 336832 153156
rect 336884 153144 336890 153196
rect 339678 153144 339684 153196
rect 339736 153184 339742 153196
rect 377306 153184 377312 153196
rect 339736 153156 377312 153184
rect 339736 153144 339742 153156
rect 377306 153144 377312 153156
rect 377364 153144 377370 153196
rect 378226 153144 378232 153196
rect 378284 153184 378290 153196
rect 379882 153184 379888 153196
rect 378284 153156 379888 153184
rect 378284 153144 378290 153156
rect 379882 153144 379888 153156
rect 379940 153144 379946 153196
rect 385034 153144 385040 153196
rect 385092 153184 385098 153196
rect 399754 153184 399760 153196
rect 385092 153156 399760 153184
rect 385092 153144 385098 153156
rect 399754 153144 399760 153156
rect 399812 153144 399818 153196
rect 402422 153144 402428 153196
rect 402480 153184 402486 153196
rect 423490 153184 423496 153196
rect 402480 153156 423496 153184
rect 402480 153144 402486 153156
rect 423490 153144 423496 153156
rect 423548 153144 423554 153196
rect 423582 153144 423588 153196
rect 423640 153184 423646 153196
rect 423640 153156 429608 153184
rect 423640 153144 423646 153156
rect 80054 153076 80060 153128
rect 80112 153116 80118 153128
rect 175090 153116 175096 153128
rect 80112 153088 175096 153116
rect 80112 153076 80118 153088
rect 175090 153076 175096 153088
rect 175148 153076 175154 153128
rect 180794 153076 180800 153128
rect 180852 153116 180858 153128
rect 257246 153116 257252 153128
rect 180852 153088 257252 153116
rect 180852 153076 180858 153088
rect 257246 153076 257252 153088
rect 257304 153076 257310 153128
rect 264974 153076 264980 153128
rect 265032 153116 265038 153128
rect 321462 153116 321468 153128
rect 265032 153088 321468 153116
rect 265032 153076 265038 153088
rect 321462 153076 321468 153088
rect 321520 153076 321526 153128
rect 324314 153076 324320 153128
rect 324372 153116 324378 153128
rect 367002 153116 367008 153128
rect 324372 153088 367008 153116
rect 324372 153076 324378 153088
rect 367002 153076 367008 153088
rect 367060 153076 367066 153128
rect 367186 153076 367192 153128
rect 367244 153116 367250 153128
rect 368934 153116 368940 153128
rect 367244 153088 368940 153116
rect 367244 153076 367250 153088
rect 368934 153076 368940 153088
rect 368992 153076 368998 153128
rect 380986 153076 380992 153128
rect 381044 153116 381050 153128
rect 410058 153116 410064 153128
rect 381044 153088 410064 153116
rect 381044 153076 381050 153088
rect 410058 153076 410064 153088
rect 410116 153076 410122 153128
rect 410702 153076 410708 153128
rect 410760 153116 410766 153128
rect 421006 153116 421012 153128
rect 410760 153088 421012 153116
rect 410760 153076 410766 153088
rect 421006 153076 421012 153088
rect 421064 153076 421070 153128
rect 422570 153076 422576 153128
rect 422628 153116 422634 153128
rect 429470 153116 429476 153128
rect 422628 153088 429476 153116
rect 422628 153076 422634 153088
rect 429470 153076 429476 153088
rect 429528 153076 429534 153128
rect 429580 153116 429608 153156
rect 430206 153144 430212 153196
rect 430264 153184 430270 153196
rect 447318 153184 447324 153196
rect 430264 153156 447324 153184
rect 430264 153144 430270 153156
rect 447318 153144 447324 153156
rect 447376 153144 447382 153196
rect 456794 153144 456800 153196
rect 456852 153184 456858 153196
rect 459462 153184 459468 153196
rect 456852 153156 459468 153184
rect 456852 153144 456858 153156
rect 459462 153144 459468 153156
rect 459520 153144 459526 153196
rect 461670 153144 461676 153196
rect 461728 153184 461734 153196
rect 465902 153184 465908 153196
rect 461728 153156 465908 153184
rect 461728 153144 461734 153156
rect 465902 153144 465908 153156
rect 465960 153144 465966 153196
rect 466454 153144 466460 153196
rect 466512 153184 466518 153196
rect 470410 153184 470416 153196
rect 466512 153156 470416 153184
rect 466512 153144 466518 153156
rect 470410 153144 470416 153156
rect 470468 153144 470474 153196
rect 471790 153144 471796 153196
rect 471848 153184 471854 153196
rect 472986 153184 472992 153196
rect 471848 153156 472992 153184
rect 471848 153144 471854 153156
rect 472986 153144 472992 153156
rect 473044 153144 473050 153196
rect 473354 153144 473360 153196
rect 473412 153184 473418 153196
rect 475562 153184 475568 153196
rect 473412 153156 475568 153184
rect 473412 153144 473418 153156
rect 475562 153144 475568 153156
rect 475620 153144 475626 153196
rect 476114 153144 476120 153196
rect 476172 153184 476178 153196
rect 478138 153184 478144 153196
rect 476172 153156 478144 153184
rect 476172 153144 476178 153156
rect 478138 153144 478144 153156
rect 478196 153144 478202 153196
rect 484026 153144 484032 153196
rect 484084 153184 484090 153196
rect 488442 153184 488448 153196
rect 484084 153156 488448 153184
rect 484084 153144 484090 153156
rect 488442 153144 488448 153156
rect 488500 153144 488506 153196
rect 489914 153144 489920 153196
rect 489972 153184 489978 153196
rect 492858 153184 492864 153196
rect 489972 153156 492864 153184
rect 489972 153144 489978 153156
rect 492858 153144 492864 153156
rect 492916 153144 492922 153196
rect 494054 153144 494060 153196
rect 494112 153184 494118 153196
rect 496078 153184 496084 153196
rect 494112 153156 496084 153184
rect 494112 153144 494118 153156
rect 496078 153144 496084 153156
rect 496136 153144 496142 153196
rect 496630 153144 496636 153196
rect 496688 153184 496694 153196
rect 498010 153184 498016 153196
rect 496688 153156 498016 153184
rect 496688 153144 496694 153156
rect 498010 153144 498016 153156
rect 498068 153144 498074 153196
rect 510982 153144 510988 153196
rect 511040 153184 511046 153196
rect 513466 153184 513472 153196
rect 511040 153156 513472 153184
rect 511040 153144 511046 153156
rect 513466 153144 513472 153156
rect 513524 153144 513530 153196
rect 514202 153144 514208 153196
rect 514260 153184 514266 153196
rect 517422 153184 517428 153196
rect 514260 153156 517428 153184
rect 514260 153144 514266 153156
rect 517422 153144 517428 153156
rect 517480 153144 517486 153196
rect 431862 153116 431868 153128
rect 429580 153088 431868 153116
rect 431862 153076 431868 153088
rect 431920 153076 431926 153128
rect 431954 153076 431960 153128
rect 432012 153116 432018 153128
rect 441982 153116 441988 153128
rect 432012 153088 441988 153116
rect 432012 153076 432018 153088
rect 441982 153076 441988 153088
rect 442040 153076 442046 153128
rect 442166 153116 442172 153128
rect 442092 153088 442172 153116
rect 103514 153008 103520 153060
rect 103572 153048 103578 153060
rect 198182 153048 198188 153060
rect 103572 153020 198188 153048
rect 103572 153008 103578 153020
rect 198182 153008 198188 153020
rect 198240 153008 198246 153060
rect 204162 153008 204168 153060
rect 204220 153048 204226 153060
rect 267550 153048 267556 153060
rect 204220 153020 267556 153048
rect 204220 153008 204226 153020
rect 267550 153008 267556 153020
rect 267608 153008 267614 153060
rect 272150 153008 272156 153060
rect 272208 153048 272214 153060
rect 326614 153048 326620 153060
rect 272208 153020 326620 153048
rect 272208 153008 272214 153020
rect 326614 153008 326620 153020
rect 326672 153008 326678 153060
rect 330938 153008 330944 153060
rect 330996 153048 331002 153060
rect 371510 153048 371516 153060
rect 330996 153020 371516 153048
rect 330996 153008 331002 153020
rect 371510 153008 371516 153020
rect 371568 153008 371574 153060
rect 375466 153008 375472 153060
rect 375524 153048 375530 153060
rect 398098 153048 398104 153060
rect 375524 153020 398104 153048
rect 375524 153008 375530 153020
rect 398098 153008 398104 153020
rect 398156 153008 398162 153060
rect 405826 153008 405832 153060
rect 405884 153048 405890 153060
rect 408770 153048 408776 153060
rect 405884 153020 408776 153048
rect 405884 153008 405890 153020
rect 408770 153008 408776 153020
rect 408828 153008 408834 153060
rect 413370 153008 413376 153060
rect 413428 153048 413434 153060
rect 416498 153048 416504 153060
rect 413428 153020 416504 153048
rect 413428 153008 413434 153020
rect 416498 153008 416504 153020
rect 416556 153008 416562 153060
rect 419258 153008 419264 153060
rect 419316 153048 419322 153060
rect 434622 153048 434628 153060
rect 419316 153020 434628 153048
rect 419316 153008 419322 153020
rect 434622 153008 434628 153020
rect 434680 153008 434686 153060
rect 436094 153008 436100 153060
rect 436152 153048 436158 153060
rect 437750 153048 437756 153060
rect 436152 153020 437756 153048
rect 436152 153008 436158 153020
rect 437750 153008 437756 153020
rect 437808 153008 437814 153060
rect 437842 153008 437848 153060
rect 437900 153048 437906 153060
rect 442092 153048 442120 153088
rect 442166 153076 442172 153088
rect 442224 153076 442230 153128
rect 449894 153116 449900 153128
rect 442276 153088 449900 153116
rect 437900 153020 442120 153048
rect 437900 153008 437906 153020
rect 92474 152940 92480 152992
rect 92532 152980 92538 152992
rect 187878 152980 187884 152992
rect 92532 152952 187884 152980
rect 92532 152940 92538 152952
rect 187878 152940 187884 152952
rect 187936 152940 187942 152992
rect 195422 152940 195428 152992
rect 195480 152980 195486 152992
rect 218698 152980 218704 152992
rect 195480 152952 218704 152980
rect 195480 152940 195486 152952
rect 218698 152940 218704 152952
rect 218756 152940 218762 152992
rect 220354 152940 220360 152992
rect 220412 152980 220418 152992
rect 284846 152980 284852 152992
rect 220412 152952 284852 152980
rect 220412 152940 220418 152952
rect 284846 152940 284852 152952
rect 284904 152940 284910 152992
rect 288158 152940 288164 152992
rect 288216 152980 288222 152992
rect 289998 152980 290004 152992
rect 288216 152952 290004 152980
rect 288216 152940 288222 152952
rect 289998 152940 290004 152952
rect 290056 152940 290062 152992
rect 291378 152940 291384 152992
rect 291436 152980 291442 152992
rect 341334 152980 341340 152992
rect 291436 152952 341340 152980
rect 291436 152940 291442 152952
rect 341334 152940 341340 152952
rect 341392 152940 341398 152992
rect 342254 152940 342260 152992
rect 342312 152980 342318 152992
rect 343910 152980 343916 152992
rect 342312 152952 343916 152980
rect 342312 152940 342318 152952
rect 343910 152940 343916 152952
rect 343968 152940 343974 152992
rect 345290 152940 345296 152992
rect 345348 152980 345354 152992
rect 382458 152980 382464 152992
rect 345348 152952 382464 152980
rect 345348 152940 345354 152952
rect 382458 152940 382464 152952
rect 382516 152940 382522 152992
rect 382550 152940 382556 152992
rect 382608 152980 382614 152992
rect 386966 152980 386972 152992
rect 382608 152952 386972 152980
rect 382608 152940 382614 152952
rect 386966 152940 386972 152952
rect 387024 152940 387030 152992
rect 390370 152940 390376 152992
rect 390428 152980 390434 152992
rect 415210 152980 415216 152992
rect 390428 152952 415216 152980
rect 390428 152940 390434 152952
rect 415210 152940 415216 152952
rect 415268 152940 415274 152992
rect 415394 152940 415400 152992
rect 415452 152980 415458 152992
rect 436370 152980 436376 152992
rect 415452 152952 436376 152980
rect 415452 152940 415458 152952
rect 436370 152940 436376 152952
rect 436428 152940 436434 152992
rect 437474 152940 437480 152992
rect 437532 152980 437538 152992
rect 441890 152980 441896 152992
rect 437532 152952 441896 152980
rect 437532 152940 437538 152952
rect 441890 152940 441896 152952
rect 441948 152940 441954 152992
rect 96614 152872 96620 152924
rect 96672 152912 96678 152924
rect 193030 152912 193036 152924
rect 96672 152884 193036 152912
rect 96672 152872 96678 152884
rect 193030 152872 193036 152884
rect 193088 152872 193094 152924
rect 212442 152872 212448 152924
rect 212500 152912 212506 152924
rect 277762 152912 277768 152924
rect 212500 152884 277768 152912
rect 212500 152872 212506 152884
rect 277762 152872 277768 152884
rect 277820 152872 277826 152924
rect 278774 152872 278780 152924
rect 278832 152912 278838 152924
rect 331766 152912 331772 152924
rect 278832 152884 331772 152912
rect 278832 152872 278838 152884
rect 331766 152872 331772 152884
rect 331824 152872 331830 152924
rect 335354 152872 335360 152924
rect 335412 152912 335418 152924
rect 375374 152912 375380 152924
rect 335412 152884 375380 152912
rect 335412 152872 335418 152884
rect 375374 152872 375380 152884
rect 375432 152872 375438 152924
rect 382182 152872 382188 152924
rect 382240 152912 382246 152924
rect 410702 152912 410708 152924
rect 382240 152884 410708 152912
rect 382240 152872 382246 152884
rect 410702 152872 410708 152884
rect 410760 152872 410766 152924
rect 411254 152872 411260 152924
rect 411312 152912 411318 152924
rect 433150 152912 433156 152924
rect 411312 152884 433156 152912
rect 411312 152872 411318 152884
rect 433150 152872 433156 152884
rect 433208 152872 433214 152924
rect 433518 152872 433524 152924
rect 433576 152912 433582 152924
rect 442276 152912 442304 153088
rect 449894 153076 449900 153088
rect 449952 153076 449958 153128
rect 463602 153076 463608 153128
rect 463660 153116 463666 153128
rect 466546 153116 466552 153128
rect 463660 153088 466552 153116
rect 463660 153076 463666 153088
rect 466546 153076 466552 153088
rect 466604 153076 466610 153128
rect 466638 153076 466644 153128
rect 466696 153116 466702 153128
rect 469766 153116 469772 153128
rect 466696 153088 469772 153116
rect 466696 153076 466702 153088
rect 469766 153076 469772 153088
rect 469824 153076 469830 153128
rect 471422 153076 471428 153128
rect 471480 153116 471486 153128
rect 473630 153116 473636 153128
rect 471480 153088 473636 153116
rect 471480 153076 471486 153088
rect 473630 153076 473636 153088
rect 473688 153076 473694 153128
rect 474826 153076 474832 153128
rect 474884 153116 474890 153128
rect 476850 153116 476856 153128
rect 474884 153088 476856 153116
rect 474884 153076 474890 153088
rect 476850 153076 476856 153088
rect 476908 153076 476914 153128
rect 484946 153076 484952 153128
rect 485004 153116 485010 153128
rect 489638 153116 489644 153128
rect 485004 153088 489644 153116
rect 485004 153076 485010 153088
rect 489638 153076 489644 153088
rect 489696 153076 489702 153128
rect 491662 153076 491668 153128
rect 491720 153116 491726 153128
rect 494790 153116 494796 153128
rect 491720 153088 494796 153116
rect 491720 153076 491726 153088
rect 494790 153076 494796 153088
rect 494848 153076 494854 153128
rect 494974 153076 494980 153128
rect 495032 153116 495038 153128
rect 496722 153116 496728 153128
rect 495032 153088 496728 153116
rect 495032 153076 495038 153088
rect 496722 153076 496728 153088
rect 496780 153076 496786 153128
rect 496814 153076 496820 153128
rect 496872 153116 496878 153128
rect 498654 153116 498660 153128
rect 496872 153088 498660 153116
rect 496872 153076 496878 153088
rect 498654 153076 498660 153088
rect 498712 153076 498718 153128
rect 512914 153076 512920 153128
rect 512972 153116 512978 153128
rect 515214 153116 515220 153128
rect 512972 153088 515220 153116
rect 512972 153076 512978 153088
rect 515214 153076 515220 153088
rect 515272 153076 515278 153128
rect 455046 153048 455052 153060
rect 433576 152884 442304 152912
rect 442368 153020 455052 153048
rect 433576 152872 433582 152884
rect 33134 152804 33140 152856
rect 33192 152844 33198 152856
rect 138014 152844 138020 152856
rect 33192 152816 138020 152844
rect 33192 152804 33198 152816
rect 138014 152804 138020 152816
rect 138072 152804 138078 152856
rect 138106 152804 138112 152856
rect 138164 152844 138170 152856
rect 141694 152844 141700 152856
rect 138164 152816 141700 152844
rect 138164 152804 138170 152816
rect 141694 152804 141700 152816
rect 141752 152804 141758 152856
rect 146478 152804 146484 152856
rect 146536 152844 146542 152856
rect 167362 152844 167368 152856
rect 146536 152816 167368 152844
rect 146536 152804 146542 152816
rect 167362 152804 167368 152816
rect 167420 152804 167426 152856
rect 173894 152804 173900 152856
rect 173952 152844 173958 152856
rect 252094 152844 252100 152856
rect 173952 152816 252100 152844
rect 173952 152804 173958 152816
rect 252094 152804 252100 152816
rect 252152 152804 252158 152856
rect 255406 152804 255412 152856
rect 255464 152844 255470 152856
rect 313090 152844 313096 152856
rect 255464 152816 313096 152844
rect 255464 152804 255470 152816
rect 313090 152804 313096 152816
rect 313148 152804 313154 152856
rect 313182 152804 313188 152856
rect 313240 152844 313246 152856
rect 356146 152844 356152 152856
rect 313240 152816 356152 152844
rect 313240 152804 313246 152816
rect 356146 152804 356152 152816
rect 356204 152804 356210 152856
rect 357434 152804 357440 152856
rect 357492 152844 357498 152856
rect 359366 152844 359372 152856
rect 357492 152816 359372 152844
rect 357492 152804 357498 152816
rect 359366 152804 359372 152816
rect 359424 152804 359430 152856
rect 361574 152804 361580 152856
rect 361632 152844 361638 152856
rect 395246 152844 395252 152856
rect 361632 152816 395252 152844
rect 361632 152804 361638 152816
rect 395246 152804 395252 152816
rect 395304 152804 395310 152856
rect 395522 152804 395528 152856
rect 395580 152844 395586 152856
rect 397822 152844 397828 152856
rect 395580 152816 397828 152844
rect 395580 152804 395586 152816
rect 397822 152804 397828 152816
rect 397880 152804 397886 152856
rect 399202 152804 399208 152856
rect 399260 152844 399266 152856
rect 424226 152844 424232 152856
rect 399260 152816 424232 152844
rect 399260 152804 399266 152816
rect 424226 152804 424232 152816
rect 424284 152804 424290 152856
rect 426158 152844 426164 152856
rect 425164 152816 426164 152844
rect 26418 152736 26424 152788
rect 26476 152776 26482 152788
rect 139118 152776 139124 152788
rect 26476 152748 139124 152776
rect 26476 152736 26482 152748
rect 139118 152736 139124 152748
rect 139176 152736 139182 152788
rect 140774 152736 140780 152788
rect 140832 152776 140838 152788
rect 144270 152776 144276 152788
rect 140832 152748 144276 152776
rect 140832 152736 140838 152748
rect 144270 152736 144276 152748
rect 144328 152736 144334 152788
rect 144362 152736 144368 152788
rect 144420 152776 144426 152788
rect 162210 152776 162216 152788
rect 144420 152748 162216 152776
rect 144420 152736 144426 152748
rect 162210 152736 162216 152748
rect 162268 152736 162274 152788
rect 164418 152736 164424 152788
rect 164476 152776 164482 152788
rect 244366 152776 244372 152788
rect 164476 152748 244372 152776
rect 164476 152736 164482 152748
rect 244366 152736 244372 152748
rect 244424 152736 244430 152788
rect 257706 152736 257712 152788
rect 257764 152776 257770 152788
rect 315666 152776 315672 152788
rect 257764 152748 315672 152776
rect 257764 152736 257770 152748
rect 315666 152736 315672 152748
rect 315724 152736 315730 152788
rect 317046 152736 317052 152788
rect 317104 152776 317110 152788
rect 318242 152776 318248 152788
rect 317104 152748 318248 152776
rect 317104 152736 317110 152748
rect 318242 152736 318248 152748
rect 318300 152736 318306 152788
rect 320266 152736 320272 152788
rect 320324 152776 320330 152788
rect 323118 152776 323124 152788
rect 320324 152748 323124 152776
rect 320324 152736 320330 152748
rect 323118 152736 323124 152748
rect 323176 152736 323182 152788
rect 324222 152736 324228 152788
rect 324280 152776 324286 152788
rect 366358 152776 366364 152788
rect 324280 152748 366364 152776
rect 324280 152736 324286 152748
rect 366358 152736 366364 152748
rect 366416 152736 366422 152788
rect 372614 152736 372620 152788
rect 372672 152776 372678 152788
rect 403618 152776 403624 152788
rect 372672 152748 403624 152776
rect 372672 152736 372678 152748
rect 403618 152736 403624 152748
rect 403676 152736 403682 152788
rect 406654 152736 406660 152788
rect 406712 152776 406718 152788
rect 422938 152776 422944 152788
rect 406712 152748 422944 152776
rect 406712 152736 406718 152748
rect 422938 152736 422944 152748
rect 422996 152736 423002 152788
rect 423490 152736 423496 152788
rect 423548 152776 423554 152788
rect 425164 152776 425192 152816
rect 426158 152804 426164 152816
rect 426216 152804 426222 152856
rect 426434 152804 426440 152856
rect 426492 152844 426498 152856
rect 440142 152844 440148 152856
rect 426492 152816 440148 152844
rect 426492 152804 426498 152816
rect 440142 152804 440148 152816
rect 440200 152804 440206 152856
rect 440234 152804 440240 152856
rect 440292 152844 440298 152856
rect 442368 152844 442396 153020
rect 455046 153008 455052 153020
rect 455104 153008 455110 153060
rect 463142 153008 463148 153060
rect 463200 153048 463206 153060
rect 467190 153048 467196 153060
rect 463200 153020 467196 153048
rect 463200 153008 463206 153020
rect 467190 153008 467196 153020
rect 467248 153008 467254 153060
rect 472158 153008 472164 153060
rect 472216 153048 472222 153060
rect 474274 153048 474280 153060
rect 472216 153020 474280 153048
rect 472216 153008 472222 153020
rect 474274 153008 474280 153020
rect 474332 153008 474338 153060
rect 484394 153008 484400 153060
rect 484452 153048 484458 153060
rect 488994 153048 489000 153060
rect 484452 153020 489000 153048
rect 484452 153008 484458 153020
rect 488994 153008 489000 153020
rect 489052 153008 489058 153060
rect 492674 153008 492680 153060
rect 492732 153048 492738 153060
rect 495434 153048 495440 153060
rect 492732 153020 495440 153048
rect 492732 153008 492738 153020
rect 495434 153008 495440 153020
rect 495492 153008 495498 153060
rect 495526 153008 495532 153060
rect 495584 153048 495590 153060
rect 497366 153048 497372 153060
rect 495584 153020 497372 153048
rect 495584 153008 495590 153020
rect 497366 153008 497372 153020
rect 497424 153008 497430 153060
rect 442534 152940 442540 152992
rect 442592 152980 442598 152992
rect 453114 152980 453120 152992
rect 442592 152952 453120 152980
rect 442592 152940 442598 152952
rect 453114 152940 453120 152952
rect 453172 152940 453178 152992
rect 464522 152940 464528 152992
rect 464580 152980 464586 152992
rect 468386 152980 468392 152992
rect 464580 152952 468392 152980
rect 464580 152940 464586 152952
rect 468386 152940 468392 152952
rect 468444 152940 468450 152992
rect 472342 152940 472348 152992
rect 472400 152980 472406 152992
rect 474918 152980 474924 152992
rect 472400 152952 474924 152980
rect 472400 152940 472406 152952
rect 474918 152940 474924 152952
rect 474976 152940 474982 152992
rect 483106 152940 483112 152992
rect 483164 152980 483170 152992
rect 487798 152980 487804 152992
rect 483164 152952 487804 152980
rect 483164 152940 483170 152952
rect 487798 152940 487804 152952
rect 487856 152940 487862 152992
rect 491294 152940 491300 152992
rect 491352 152980 491358 152992
rect 494146 152980 494152 152992
rect 491352 152952 494152 152980
rect 491352 152940 491358 152952
rect 494146 152940 494152 152952
rect 494204 152940 494210 152992
rect 512270 152940 512276 152992
rect 512328 152980 512334 152992
rect 514754 152980 514760 152992
rect 512328 152952 514760 152980
rect 512328 152940 512334 152952
rect 514754 152940 514760 152952
rect 514812 152940 514818 152992
rect 442994 152872 443000 152924
rect 443052 152912 443058 152924
rect 451182 152912 451188 152924
rect 443052 152884 451188 152912
rect 443052 152872 443058 152884
rect 451182 152872 451188 152884
rect 451240 152872 451246 152924
rect 465074 152872 465080 152924
rect 465132 152912 465138 152924
rect 469122 152912 469128 152924
rect 465132 152884 469128 152912
rect 465132 152872 465138 152884
rect 469122 152872 469128 152884
rect 469180 152872 469186 152924
rect 490006 152872 490012 152924
rect 490064 152912 490070 152924
rect 493502 152912 493508 152924
rect 490064 152884 493508 152912
rect 490064 152872 490070 152884
rect 493502 152872 493508 152884
rect 493560 152872 493566 152924
rect 440292 152816 442396 152844
rect 440292 152804 440298 152816
rect 442442 152804 442448 152856
rect 442500 152844 442506 152856
rect 444374 152844 444380 152856
rect 442500 152816 444380 152844
rect 442500 152804 442506 152816
rect 444374 152804 444380 152816
rect 444432 152804 444438 152856
rect 446306 152804 446312 152856
rect 446364 152844 446370 152856
rect 460014 152844 460020 152856
rect 446364 152816 460020 152844
rect 446364 152804 446370 152816
rect 460014 152804 460020 152816
rect 460072 152804 460078 152856
rect 510338 152804 510344 152856
rect 510396 152844 510402 152856
rect 511994 152844 512000 152856
rect 510396 152816 512000 152844
rect 510396 152804 510402 152816
rect 511994 152804 512000 152816
rect 512052 152804 512058 152856
rect 423548 152748 425192 152776
rect 423548 152736 423554 152748
rect 425238 152736 425244 152788
rect 425296 152776 425302 152788
rect 434254 152776 434260 152788
rect 425296 152748 434260 152776
rect 425296 152736 425302 152748
rect 434254 152736 434260 152748
rect 434312 152736 434318 152788
rect 434346 152736 434352 152788
rect 434404 152776 434410 152788
rect 450538 152776 450544 152788
rect 434404 152748 450544 152776
rect 434404 152736 434410 152748
rect 450538 152736 450544 152748
rect 450596 152736 450602 152788
rect 28166 152668 28172 152720
rect 28224 152708 28230 152720
rect 141050 152708 141056 152720
rect 28224 152680 141056 152708
rect 28224 152668 28230 152680
rect 141050 152668 141056 152680
rect 141108 152668 141114 152720
rect 142798 152668 142804 152720
rect 142856 152708 142862 152720
rect 149422 152708 149428 152720
rect 142856 152680 149428 152708
rect 142856 152668 142862 152680
rect 149422 152668 149428 152680
rect 149480 152668 149486 152720
rect 149514 152668 149520 152720
rect 149572 152708 149578 152720
rect 231578 152708 231584 152720
rect 149572 152680 231584 152708
rect 149572 152668 149578 152680
rect 231578 152668 231584 152680
rect 231636 152668 231642 152720
rect 240318 152668 240324 152720
rect 240376 152708 240382 152720
rect 241882 152708 241888 152720
rect 240376 152680 241888 152708
rect 240376 152668 240382 152680
rect 241882 152668 241888 152680
rect 241940 152668 241946 152720
rect 247034 152668 247040 152720
rect 247092 152708 247098 152720
rect 307938 152708 307944 152720
rect 247092 152680 307944 152708
rect 247092 152668 247098 152680
rect 307938 152668 307944 152680
rect 307996 152668 308002 152720
rect 318334 152668 318340 152720
rect 318392 152708 318398 152720
rect 361942 152708 361948 152720
rect 318392 152680 361948 152708
rect 318392 152668 318398 152680
rect 361942 152668 361948 152680
rect 362000 152668 362006 152720
rect 368474 152668 368480 152720
rect 368532 152708 368538 152720
rect 400398 152708 400404 152720
rect 368532 152680 400404 152708
rect 368532 152668 368538 152680
rect 400398 152668 400404 152680
rect 400456 152668 400462 152720
rect 404354 152668 404360 152720
rect 404412 152708 404418 152720
rect 427998 152708 428004 152720
rect 404412 152680 428004 152708
rect 404412 152668 404418 152680
rect 427998 152668 428004 152680
rect 428056 152668 428062 152720
rect 430574 152668 430580 152720
rect 430632 152708 430638 152720
rect 447962 152708 447968 152720
rect 430632 152680 447968 152708
rect 430632 152668 430638 152680
rect 447962 152668 447968 152680
rect 448020 152668 448026 152720
rect 22186 152600 22192 152652
rect 22244 152640 22250 152652
rect 135898 152640 135904 152652
rect 22244 152612 135904 152640
rect 22244 152600 22250 152612
rect 135898 152600 135904 152612
rect 135956 152600 135962 152652
rect 151906 152640 151912 152652
rect 137986 152612 151912 152640
rect 19334 152532 19340 152584
rect 19392 152572 19398 152584
rect 133966 152572 133972 152584
rect 19392 152544 133972 152572
rect 19392 152532 19398 152544
rect 133966 152532 133972 152544
rect 134024 152532 134030 152584
rect 136818 152532 136824 152584
rect 136876 152572 136882 152584
rect 137986 152572 138014 152612
rect 151906 152600 151912 152612
rect 151964 152600 151970 152652
rect 153562 152600 153568 152652
rect 153620 152640 153626 152652
rect 236730 152640 236736 152652
rect 153620 152612 236736 152640
rect 153620 152600 153626 152612
rect 236730 152600 236736 152612
rect 236788 152600 236794 152652
rect 244458 152600 244464 152652
rect 244516 152640 244522 152652
rect 306006 152640 306012 152652
rect 244516 152612 306012 152640
rect 244516 152600 244522 152612
rect 306006 152600 306012 152612
rect 306064 152600 306070 152652
rect 311526 152600 311532 152652
rect 311584 152640 311590 152652
rect 356790 152640 356796 152652
rect 311584 152612 356796 152640
rect 311584 152600 311590 152612
rect 356790 152600 356796 152612
rect 356848 152600 356854 152652
rect 358814 152600 358820 152652
rect 358872 152640 358878 152652
rect 393406 152640 393412 152652
rect 358872 152612 393412 152640
rect 358872 152600 358878 152612
rect 393406 152600 393412 152612
rect 393464 152600 393470 152652
rect 394878 152600 394884 152652
rect 394936 152640 394942 152652
rect 420362 152640 420368 152652
rect 394936 152612 420368 152640
rect 394936 152600 394942 152612
rect 420362 152600 420368 152612
rect 420420 152600 420426 152652
rect 421374 152600 421380 152652
rect 421432 152640 421438 152652
rect 421432 152612 434208 152640
rect 421432 152600 421438 152612
rect 136876 152544 138014 152572
rect 136876 152532 136882 152544
rect 138106 152532 138112 152584
rect 138164 152572 138170 152584
rect 144270 152572 144276 152584
rect 138164 152544 144276 152572
rect 138164 152532 138170 152544
rect 144270 152532 144276 152544
rect 144328 152532 144334 152584
rect 144362 152532 144368 152584
rect 144420 152572 144426 152584
rect 226426 152572 226432 152584
rect 144420 152544 226432 152572
rect 144420 152532 144426 152544
rect 226426 152532 226432 152544
rect 226484 152532 226490 152584
rect 234154 152532 234160 152584
rect 234212 152572 234218 152584
rect 297726 152572 297732 152584
rect 234212 152544 297732 152572
rect 234212 152532 234218 152544
rect 297726 152532 297732 152544
rect 297784 152532 297790 152584
rect 304810 152532 304816 152584
rect 304868 152572 304874 152584
rect 351638 152572 351644 152584
rect 304868 152544 351644 152572
rect 304868 152532 304874 152544
rect 351638 152532 351644 152544
rect 351696 152532 351702 152584
rect 352006 152532 352012 152584
rect 352064 152572 352070 152584
rect 388254 152572 388260 152584
rect 352064 152544 388260 152572
rect 352064 152532 352070 152544
rect 388254 152532 388260 152544
rect 388312 152532 388318 152584
rect 388346 152532 388352 152584
rect 388404 152572 388410 152584
rect 392210 152572 392216 152584
rect 388404 152544 392216 152572
rect 388404 152532 388410 152544
rect 392210 152532 392216 152544
rect 392268 152532 392274 152584
rect 393130 152532 393136 152584
rect 393188 152572 393194 152584
rect 419074 152572 419080 152584
rect 393188 152544 419080 152572
rect 393188 152532 393194 152544
rect 419074 152532 419080 152544
rect 419132 152532 419138 152584
rect 419534 152532 419540 152584
rect 419592 152572 419598 152584
rect 419810 152572 419816 152584
rect 419592 152544 419816 152572
rect 419592 152532 419598 152544
rect 419810 152532 419816 152544
rect 419868 152532 419874 152584
rect 421006 152532 421012 152584
rect 421064 152572 421070 152584
rect 423306 152572 423312 152584
rect 421064 152544 423312 152572
rect 421064 152532 421070 152544
rect 423306 152532 423312 152544
rect 423364 152532 423370 152584
rect 423398 152532 423404 152584
rect 423456 152572 423462 152584
rect 434180 152572 434208 152612
rect 434254 152600 434260 152652
rect 434312 152640 434318 152652
rect 436922 152640 436928 152652
rect 434312 152612 436928 152640
rect 434312 152600 434318 152612
rect 436922 152600 436928 152612
rect 436980 152600 436986 152652
rect 437014 152600 437020 152652
rect 437072 152640 437078 152652
rect 438946 152640 438952 152652
rect 437072 152612 438952 152640
rect 437072 152600 437078 152612
rect 438946 152600 438952 152612
rect 439004 152600 439010 152652
rect 440326 152600 440332 152652
rect 440384 152640 440390 152652
rect 455690 152640 455696 152652
rect 440384 152612 455696 152640
rect 440384 152600 440390 152612
rect 455690 152600 455696 152612
rect 455748 152600 455754 152652
rect 440878 152572 440884 152584
rect 423456 152544 434024 152572
rect 434180 152544 440884 152572
rect 423456 152532 423462 152544
rect 2866 152464 2872 152516
rect 2924 152504 2930 152516
rect 121086 152504 121092 152516
rect 2924 152476 121092 152504
rect 2924 152464 2930 152476
rect 121086 152464 121092 152476
rect 121144 152464 121150 152516
rect 126974 152464 126980 152516
rect 127032 152504 127038 152516
rect 216122 152504 216128 152516
rect 127032 152476 216128 152504
rect 127032 152464 127038 152476
rect 216122 152464 216128 152476
rect 216180 152464 216186 152516
rect 227714 152464 227720 152516
rect 227772 152504 227778 152516
rect 293218 152504 293224 152516
rect 227772 152476 293224 152504
rect 227772 152464 227778 152476
rect 293218 152464 293224 152476
rect 293276 152464 293282 152516
rect 298646 152464 298652 152516
rect 298704 152504 298710 152516
rect 347130 152504 347136 152516
rect 298704 152476 347136 152504
rect 298704 152464 298710 152476
rect 347130 152464 347136 152476
rect 347188 152464 347194 152516
rect 347958 152464 347964 152516
rect 348016 152504 348022 152516
rect 385034 152504 385040 152516
rect 348016 152476 385040 152504
rect 348016 152464 348022 152476
rect 385034 152464 385040 152476
rect 385092 152464 385098 152516
rect 386414 152464 386420 152516
rect 386472 152504 386478 152516
rect 413922 152504 413928 152516
rect 386472 152476 413928 152504
rect 386472 152464 386478 152476
rect 413922 152464 413928 152476
rect 413980 152464 413986 152516
rect 414382 152464 414388 152516
rect 414440 152504 414446 152516
rect 414440 152476 433932 152504
rect 414440 152464 414446 152476
rect 67082 152396 67088 152448
rect 67140 152436 67146 152448
rect 159634 152436 159640 152448
rect 67140 152408 159640 152436
rect 67140 152396 67146 152408
rect 159634 152396 159640 152408
rect 159692 152396 159698 152448
rect 173250 152396 173256 152448
rect 173308 152436 173314 152448
rect 249518 152436 249524 152448
rect 173308 152408 249524 152436
rect 173308 152396 173314 152408
rect 249518 152396 249524 152408
rect 249576 152396 249582 152448
rect 251174 152396 251180 152448
rect 251232 152436 251238 152448
rect 311158 152436 311164 152448
rect 251232 152408 311164 152436
rect 251232 152396 251238 152408
rect 311158 152396 311164 152408
rect 311216 152396 311222 152448
rect 317414 152396 317420 152448
rect 317472 152436 317478 152448
rect 361298 152436 361304 152448
rect 317472 152408 361304 152436
rect 317472 152396 317478 152408
rect 361298 152396 361304 152408
rect 361356 152396 361362 152448
rect 365714 152396 365720 152448
rect 365772 152436 365778 152448
rect 398466 152436 398472 152448
rect 365772 152408 398472 152436
rect 365772 152396 365778 152408
rect 398466 152396 398472 152408
rect 398524 152396 398530 152448
rect 398558 152396 398564 152448
rect 398616 152436 398622 152448
rect 408126 152436 408132 152448
rect 398616 152408 408132 152436
rect 398616 152396 398622 152408
rect 408126 152396 408132 152408
rect 408184 152396 408190 152448
rect 412818 152396 412824 152448
rect 412876 152436 412882 152448
rect 412876 152408 432184 152436
rect 412876 152396 412882 152408
rect 120074 152328 120080 152380
rect 120132 152368 120138 152380
rect 211062 152368 211068 152380
rect 120132 152340 211068 152368
rect 120132 152328 120138 152340
rect 211062 152328 211068 152340
rect 211120 152328 211126 152380
rect 224586 152328 224592 152380
rect 224644 152368 224650 152380
rect 288066 152368 288072 152380
rect 224644 152340 288072 152368
rect 224644 152328 224650 152340
rect 288066 152328 288072 152340
rect 288124 152328 288130 152380
rect 292206 152328 292212 152380
rect 292264 152368 292270 152380
rect 341978 152368 341984 152380
rect 292264 152340 341984 152368
rect 292264 152328 292270 152340
rect 341978 152328 341984 152340
rect 342036 152328 342042 152380
rect 343634 152328 343640 152380
rect 343692 152368 343698 152380
rect 349798 152368 349804 152380
rect 343692 152340 349804 152368
rect 343692 152328 343698 152340
rect 349798 152328 349804 152340
rect 349856 152328 349862 152380
rect 349890 152328 349896 152380
rect 349948 152368 349954 152380
rect 385678 152368 385684 152380
rect 349948 152340 385684 152368
rect 349948 152328 349954 152340
rect 385678 152328 385684 152340
rect 385736 152328 385742 152380
rect 385770 152328 385776 152380
rect 385828 152368 385834 152380
rect 387610 152368 387616 152380
rect 385828 152340 387616 152368
rect 385828 152328 385834 152340
rect 387610 152328 387616 152340
rect 387668 152328 387674 152380
rect 389174 152328 389180 152380
rect 389232 152368 389238 152380
rect 412634 152368 412640 152380
rect 389232 152340 412640 152368
rect 389232 152328 389238 152340
rect 412634 152328 412640 152340
rect 412692 152328 412698 152380
rect 415854 152328 415860 152380
rect 415912 152368 415918 152380
rect 426802 152368 426808 152380
rect 415912 152340 426808 152368
rect 415912 152328 415918 152340
rect 426802 152328 426808 152340
rect 426860 152328 426866 152380
rect 426894 152328 426900 152380
rect 426952 152368 426958 152380
rect 432046 152368 432052 152380
rect 426952 152340 432052 152368
rect 426952 152328 426958 152340
rect 432046 152328 432052 152340
rect 432104 152328 432110 152380
rect 432156 152368 432184 152408
rect 433794 152368 433800 152380
rect 432156 152340 433800 152368
rect 433794 152328 433800 152340
rect 433852 152328 433858 152380
rect 433904 152368 433932 152476
rect 433996 152436 434024 152544
rect 440878 152532 440884 152544
rect 440936 152532 440942 152584
rect 442074 152532 442080 152584
rect 442132 152572 442138 152584
rect 456978 152572 456984 152584
rect 442132 152544 456984 152572
rect 442132 152532 442138 152544
rect 456978 152532 456984 152544
rect 457036 152532 457042 152584
rect 459554 152532 459560 152584
rect 459612 152572 459618 152584
rect 464614 152572 464620 152584
rect 459612 152544 464620 152572
rect 459612 152532 459618 152544
rect 464614 152532 464620 152544
rect 464672 152532 464678 152584
rect 454402 152504 454408 152516
rect 444116 152476 454408 152504
rect 442166 152436 442172 152448
rect 433996 152408 442172 152436
rect 442166 152396 442172 152408
rect 442224 152396 442230 152448
rect 434530 152368 434536 152380
rect 433904 152340 434536 152368
rect 434530 152328 434536 152340
rect 434588 152328 434594 152380
rect 434622 152328 434628 152380
rect 434680 152368 434686 152380
rect 437014 152368 437020 152380
rect 434680 152340 437020 152368
rect 434680 152328 434686 152340
rect 437014 152328 437020 152340
rect 437072 152328 437078 152380
rect 437750 152328 437756 152380
rect 437808 152368 437814 152380
rect 437808 152340 438532 152368
rect 437808 152328 437814 152340
rect 91094 152260 91100 152312
rect 91152 152300 91158 152312
rect 180242 152300 180248 152312
rect 91152 152272 180248 152300
rect 91152 152260 91158 152272
rect 180242 152260 180248 152272
rect 180300 152260 180306 152312
rect 187970 152260 187976 152312
rect 188028 152300 188034 152312
rect 262398 152300 262404 152312
rect 188028 152272 262404 152300
rect 188028 152260 188034 152272
rect 262398 152260 262404 152272
rect 262456 152260 262462 152312
rect 266354 152260 266360 152312
rect 266412 152300 266418 152312
rect 320818 152300 320824 152312
rect 266412 152272 320824 152300
rect 266412 152260 266418 152272
rect 320818 152260 320824 152272
rect 320876 152260 320882 152312
rect 325878 152260 325884 152312
rect 325936 152300 325942 152312
rect 367646 152300 367652 152312
rect 325936 152272 367652 152300
rect 325936 152260 325942 152272
rect 367646 152260 367652 152272
rect 367704 152260 367710 152312
rect 371326 152260 371332 152312
rect 371384 152300 371390 152312
rect 402330 152300 402336 152312
rect 371384 152272 402336 152300
rect 371384 152260 371390 152272
rect 402330 152260 402336 152272
rect 402388 152260 402394 152312
rect 404262 152260 404268 152312
rect 404320 152300 404326 152312
rect 405090 152300 405096 152312
rect 404320 152272 405096 152300
rect 404320 152260 404326 152272
rect 405090 152260 405096 152272
rect 405148 152260 405154 152312
rect 409230 152260 409236 152312
rect 409288 152300 409294 152312
rect 417878 152300 417884 152312
rect 409288 152272 417884 152300
rect 409288 152260 409294 152272
rect 417878 152260 417884 152272
rect 417936 152260 417942 152312
rect 419902 152260 419908 152312
rect 419960 152300 419966 152312
rect 428642 152300 428648 152312
rect 419960 152272 428648 152300
rect 419960 152260 419966 152272
rect 428642 152260 428648 152272
rect 428700 152260 428706 152312
rect 429286 152260 429292 152312
rect 429344 152300 429350 152312
rect 438394 152300 438400 152312
rect 429344 152272 438400 152300
rect 429344 152260 429350 152272
rect 438394 152260 438400 152272
rect 438452 152260 438458 152312
rect 109034 152192 109040 152244
rect 109092 152232 109098 152244
rect 130746 152232 130752 152244
rect 109092 152204 130752 152232
rect 109092 152192 109098 152204
rect 130746 152192 130752 152204
rect 130804 152192 130810 152244
rect 134058 152192 134064 152244
rect 134116 152232 134122 152244
rect 221274 152232 221280 152244
rect 134116 152204 221280 152232
rect 134116 152192 134122 152204
rect 221274 152192 221280 152204
rect 221332 152192 221338 152244
rect 221458 152192 221464 152244
rect 221516 152232 221522 152244
rect 282914 152232 282920 152244
rect 221516 152204 282920 152232
rect 221516 152192 221522 152204
rect 282914 152192 282920 152204
rect 282972 152192 282978 152244
rect 285766 152192 285772 152244
rect 285824 152232 285830 152244
rect 336182 152232 336188 152244
rect 285824 152204 336188 152232
rect 285824 152192 285830 152204
rect 336182 152192 336188 152204
rect 336240 152192 336246 152244
rect 342438 152192 342444 152244
rect 342496 152232 342502 152244
rect 344554 152232 344560 152244
rect 342496 152204 344560 152232
rect 342496 152192 342502 152204
rect 344554 152192 344560 152204
rect 344612 152192 344618 152244
rect 349154 152192 349160 152244
rect 349212 152232 349218 152244
rect 349890 152232 349896 152244
rect 349212 152204 349896 152232
rect 349212 152192 349218 152204
rect 349890 152192 349896 152204
rect 349948 152192 349954 152244
rect 354490 152192 354496 152244
rect 354548 152232 354554 152244
rect 389542 152232 389548 152244
rect 354548 152204 389548 152232
rect 354548 152192 354554 152204
rect 389542 152192 389548 152204
rect 389600 152192 389606 152244
rect 394602 152192 394608 152244
rect 394660 152232 394666 152244
rect 417786 152232 417792 152244
rect 394660 152204 417792 152232
rect 394660 152192 394666 152204
rect 417786 152192 417792 152204
rect 417844 152192 417850 152244
rect 419810 152192 419816 152244
rect 419868 152232 419874 152244
rect 421742 152232 421748 152244
rect 419868 152204 421748 152232
rect 419868 152192 419874 152204
rect 421742 152192 421748 152204
rect 421800 152192 421806 152244
rect 422938 152192 422944 152244
rect 422996 152232 423002 152244
rect 429378 152232 429384 152244
rect 422996 152204 429384 152232
rect 422996 152192 423002 152204
rect 429378 152192 429384 152204
rect 429436 152192 429442 152244
rect 429470 152192 429476 152244
rect 429528 152232 429534 152244
rect 431954 152232 431960 152244
rect 429528 152204 431960 152232
rect 429528 152192 429534 152204
rect 431954 152192 431960 152204
rect 432012 152192 432018 152244
rect 432046 152192 432052 152244
rect 432104 152232 432110 152244
rect 438302 152232 438308 152244
rect 432104 152204 438308 152232
rect 432104 152192 432110 152204
rect 438302 152192 438308 152204
rect 438360 152192 438366 152244
rect 438504 152232 438532 152340
rect 438854 152328 438860 152380
rect 438912 152368 438918 152380
rect 444116 152368 444144 152476
rect 454402 152464 454408 152476
rect 454460 152464 454466 152516
rect 452470 152436 452476 152448
rect 444300 152408 452476 152436
rect 438912 152340 444144 152368
rect 438912 152328 438918 152340
rect 444190 152328 444196 152380
rect 444248 152368 444254 152380
rect 444300 152368 444328 152408
rect 452470 152396 452476 152408
rect 452528 152396 452534 152448
rect 444248 152340 444328 152368
rect 444248 152328 444254 152340
rect 444374 152328 444380 152380
rect 444432 152368 444438 152380
rect 453758 152368 453764 152380
rect 444432 152340 453764 152368
rect 444432 152328 444438 152340
rect 453758 152328 453764 152340
rect 453816 152328 453822 152380
rect 511626 152328 511632 152380
rect 511684 152368 511690 152380
rect 513558 152368 513564 152380
rect 511684 152340 513564 152368
rect 511684 152328 511690 152340
rect 513558 152328 513564 152340
rect 513616 152328 513622 152380
rect 438578 152260 438584 152312
rect 438636 152300 438642 152312
rect 446674 152300 446680 152312
rect 438636 152272 446680 152300
rect 438636 152260 438642 152272
rect 446674 152260 446680 152272
rect 446732 152260 446738 152312
rect 441430 152232 441436 152244
rect 438504 152204 441436 152232
rect 441430 152192 441436 152204
rect 441488 152192 441494 152244
rect 441614 152192 441620 152244
rect 441672 152232 441678 152244
rect 456334 152232 456340 152244
rect 441672 152204 456340 152232
rect 441672 152192 441678 152204
rect 456334 152192 456340 152204
rect 456392 152192 456398 152244
rect 513558 152192 513564 152244
rect 513616 152232 513622 152244
rect 516134 152232 516140 152244
rect 513616 152204 516140 152232
rect 513616 152192 513622 152204
rect 516134 152192 516140 152204
rect 516192 152192 516198 152244
rect 82814 152124 82820 152176
rect 82872 152164 82878 152176
rect 169938 152164 169944 152176
rect 82872 152136 169944 152164
rect 82872 152124 82878 152136
rect 169938 152124 169944 152136
rect 169996 152124 170002 152176
rect 172146 152124 172152 152176
rect 172204 152164 172210 152176
rect 190454 152164 190460 152176
rect 172204 152136 190460 152164
rect 172204 152124 172210 152136
rect 190454 152124 190460 152136
rect 190512 152124 190518 152176
rect 194134 152124 194140 152176
rect 194192 152164 194198 152176
rect 213546 152164 213552 152176
rect 194192 152136 213552 152164
rect 194192 152124 194198 152136
rect 213546 152124 213552 152136
rect 213604 152124 213610 152176
rect 274542 152164 274548 152176
rect 219406 152136 274548 152164
rect 79318 152056 79324 152108
rect 79376 152096 79382 152108
rect 164786 152096 164792 152108
rect 79376 152068 164792 152096
rect 79376 152056 79382 152068
rect 164786 152056 164792 152068
rect 164844 152056 164850 152108
rect 166994 152056 167000 152108
rect 167052 152096 167058 152108
rect 182726 152096 182732 152108
rect 167052 152068 182732 152096
rect 167052 152056 167058 152068
rect 182726 152056 182732 152068
rect 182784 152056 182790 152108
rect 183462 152056 183468 152108
rect 183520 152096 183526 152108
rect 200758 152096 200764 152108
rect 183520 152068 200764 152096
rect 183520 152056 183526 152068
rect 200758 152056 200764 152068
rect 200816 152056 200822 152108
rect 212718 152056 212724 152108
rect 212776 152096 212782 152108
rect 219406 152096 219434 152136
rect 274542 152124 274548 152136
rect 274600 152124 274606 152176
rect 277394 152124 277400 152176
rect 277452 152164 277458 152176
rect 331122 152164 331128 152176
rect 277452 152136 331128 152164
rect 277452 152124 277458 152136
rect 331122 152124 331128 152136
rect 331180 152124 331186 152176
rect 332594 152124 332600 152176
rect 332652 152164 332658 152176
rect 372798 152164 372804 152176
rect 332652 152136 372804 152164
rect 332652 152124 332658 152136
rect 372798 152124 372804 152136
rect 372856 152124 372862 152176
rect 384942 152124 384948 152176
rect 385000 152164 385006 152176
rect 392118 152164 392124 152176
rect 385000 152136 392124 152164
rect 385000 152124 385006 152136
rect 392118 152124 392124 152136
rect 392176 152124 392182 152176
rect 392210 152124 392216 152176
rect 392268 152164 392274 152176
rect 407482 152164 407488 152176
rect 392268 152136 407488 152164
rect 392268 152124 392274 152136
rect 407482 152124 407488 152136
rect 407540 152124 407546 152176
rect 408494 152124 408500 152176
rect 408552 152164 408558 152176
rect 423582 152164 423588 152176
rect 408552 152136 423588 152164
rect 408552 152124 408558 152136
rect 423582 152124 423588 152136
rect 423640 152124 423646 152176
rect 423674 152124 423680 152176
rect 423732 152164 423738 152176
rect 427078 152164 427084 152176
rect 423732 152136 427084 152164
rect 423732 152124 423738 152136
rect 427078 152124 427084 152136
rect 427136 152124 427142 152176
rect 427814 152124 427820 152176
rect 427872 152164 427878 152176
rect 427872 152136 436784 152164
rect 427872 152124 427878 152136
rect 212776 152068 219434 152096
rect 212776 152056 212782 152068
rect 225322 152056 225328 152108
rect 225380 152096 225386 152108
rect 229002 152096 229008 152108
rect 225380 152068 229008 152096
rect 225380 152056 225386 152068
rect 229002 152056 229008 152068
rect 229060 152056 229066 152108
rect 243354 152056 243360 152108
rect 243412 152096 243418 152108
rect 302878 152096 302884 152108
rect 243412 152068 302884 152096
rect 243412 152056 243418 152068
rect 302878 152056 302884 152068
rect 302936 152056 302942 152108
rect 303706 152056 303712 152108
rect 303764 152096 303770 152108
rect 350994 152096 351000 152108
rect 303764 152068 351000 152096
rect 303764 152056 303770 152068
rect 350994 152056 351000 152068
rect 351052 152056 351058 152108
rect 354674 152056 354680 152108
rect 354732 152096 354738 152108
rect 390186 152096 390192 152108
rect 354732 152068 390192 152096
rect 354732 152056 354738 152068
rect 390186 152056 390192 152068
rect 390244 152056 390250 152108
rect 398834 152056 398840 152108
rect 398892 152096 398898 152108
rect 398892 152068 405044 152096
rect 398892 152056 398898 152068
rect 68830 151988 68836 152040
rect 68888 152028 68894 152040
rect 142798 152028 142804 152040
rect 68888 152000 142804 152028
rect 68888 151988 68894 152000
rect 142798 151988 142804 152000
rect 142856 151988 142862 152040
rect 143442 151988 143448 152040
rect 143500 152028 143506 152040
rect 146938 152028 146944 152040
rect 143500 152000 146944 152028
rect 143500 151988 143506 152000
rect 146938 151988 146944 152000
rect 146996 151988 147002 152040
rect 156322 151988 156328 152040
rect 156380 152028 156386 152040
rect 172514 152028 172520 152040
rect 156380 152000 172520 152028
rect 156380 151988 156386 152000
rect 172514 151988 172520 152000
rect 172572 151988 172578 152040
rect 191466 151988 191472 152040
rect 191524 152028 191530 152040
rect 208486 152028 208492 152040
rect 191524 152000 208492 152028
rect 191524 151988 191530 152000
rect 208486 151988 208492 152000
rect 208544 151988 208550 152040
rect 242434 151988 242440 152040
rect 242492 152028 242498 152040
rect 300946 152028 300952 152040
rect 242492 152000 300952 152028
rect 242492 151988 242498 152000
rect 300946 151988 300952 152000
rect 301004 151988 301010 152040
rect 307386 151988 307392 152040
rect 307444 152028 307450 152040
rect 352282 152028 352288 152040
rect 307444 152000 352288 152028
rect 307444 151988 307450 152000
rect 352282 151988 352288 152000
rect 352340 151988 352346 152040
rect 364518 151988 364524 152040
rect 364576 152028 364582 152040
rect 397178 152028 397184 152040
rect 364576 152000 397184 152028
rect 364576 151988 364582 152000
rect 397178 151988 397184 152000
rect 397236 151988 397242 152040
rect 75454 151920 75460 151972
rect 75512 151960 75518 151972
rect 154482 151960 154488 151972
rect 75512 151932 154488 151960
rect 75512 151920 75518 151932
rect 154482 151920 154488 151932
rect 154540 151920 154546 151972
rect 162486 151920 162492 151972
rect 162544 151960 162550 151972
rect 177666 151960 177672 151972
rect 162544 151932 177672 151960
rect 162544 151920 162550 151932
rect 177666 151920 177672 151932
rect 177724 151920 177730 151972
rect 184382 151920 184388 151972
rect 184440 151960 184446 151972
rect 195606 151960 195612 151972
rect 184440 151932 195612 151960
rect 184440 151920 184446 151932
rect 195606 151920 195612 151932
rect 195664 151920 195670 151972
rect 213730 151920 213736 151972
rect 213788 151960 213794 151972
rect 272702 151960 272708 151972
rect 213788 151932 272708 151960
rect 213788 151920 213794 151932
rect 272702 151920 272708 151932
rect 272760 151920 272766 151972
rect 272794 151920 272800 151972
rect 272852 151960 272858 151972
rect 325970 151960 325976 151972
rect 272852 151932 325976 151960
rect 272852 151920 272858 151932
rect 325970 151920 325976 151932
rect 326028 151920 326034 151972
rect 331214 151920 331220 151972
rect 331272 151960 331278 151972
rect 372154 151960 372160 151972
rect 331272 151932 372160 151960
rect 331272 151920 331278 151932
rect 372154 151920 372160 151932
rect 372212 151920 372218 151972
rect 378778 151920 378784 151972
rect 378836 151960 378842 151972
rect 384390 151960 384396 151972
rect 378836 151932 384396 151960
rect 378836 151920 378842 151932
rect 384390 151920 384396 151932
rect 384448 151920 384454 151972
rect 388438 151920 388444 151972
rect 388496 151960 388502 151972
rect 404906 151960 404912 151972
rect 388496 151932 404912 151960
rect 388496 151920 388502 151932
rect 404906 151920 404912 151932
rect 404964 151920 404970 151972
rect 405016 151960 405044 152068
rect 405642 152056 405648 152108
rect 405700 152096 405706 152108
rect 421006 152096 421012 152108
rect 405700 152068 421012 152096
rect 405700 152056 405706 152068
rect 421006 152056 421012 152068
rect 421064 152056 421070 152108
rect 434438 152096 434444 152108
rect 421116 152068 434444 152096
rect 405090 151988 405096 152040
rect 405148 152028 405154 152040
rect 418430 152028 418436 152040
rect 405148 152000 418436 152028
rect 405148 151988 405154 152000
rect 418430 151988 418436 152000
rect 418488 151988 418494 152040
rect 419626 151988 419632 152040
rect 419684 152028 419690 152040
rect 421116 152028 421144 152068
rect 434438 152056 434444 152068
rect 434496 152056 434502 152108
rect 434714 152056 434720 152108
rect 434772 152096 434778 152108
rect 435726 152096 435732 152108
rect 434772 152068 435732 152096
rect 434772 152056 434778 152068
rect 435726 152056 435732 152068
rect 435784 152056 435790 152108
rect 436756 152096 436784 152136
rect 436830 152124 436836 152176
rect 436888 152164 436894 152176
rect 443454 152164 443460 152176
rect 436888 152136 443460 152164
rect 436888 152124 436894 152136
rect 443454 152124 443460 152136
rect 443512 152124 443518 152176
rect 445202 152164 445208 152176
rect 444300 152136 445208 152164
rect 444300 152096 444328 152136
rect 445202 152124 445208 152136
rect 445260 152124 445266 152176
rect 445294 152124 445300 152176
rect 445352 152164 445358 152176
rect 458818 152164 458824 152176
rect 445352 152136 458824 152164
rect 445352 152124 445358 152136
rect 458818 152124 458824 152136
rect 458876 152124 458882 152176
rect 436756 152068 444328 152096
rect 444374 152056 444380 152108
rect 444432 152096 444438 152108
rect 449250 152096 449256 152108
rect 444432 152068 449256 152096
rect 444432 152056 444438 152068
rect 449250 152056 449256 152068
rect 449308 152056 449314 152108
rect 419684 152000 421144 152028
rect 419684 151988 419690 152000
rect 425054 151988 425060 152040
rect 425112 152028 425118 152040
rect 436830 152028 436836 152040
rect 425112 152000 436836 152028
rect 425112 151988 425118 152000
rect 436830 151988 436836 152000
rect 436888 151988 436894 152040
rect 436922 151988 436928 152040
rect 436980 152028 436986 152040
rect 444098 152028 444104 152040
rect 436980 152000 444104 152028
rect 436980 151988 436986 152000
rect 444098 151988 444104 152000
rect 444156 151988 444162 152040
rect 444466 151988 444472 152040
rect 444524 152028 444530 152040
rect 458174 152028 458180 152040
rect 444524 152000 458180 152028
rect 444524 151988 444530 152000
rect 458174 151988 458180 152000
rect 458232 151988 458238 152040
rect 467834 151988 467840 152040
rect 467892 152028 467898 152040
rect 471698 152028 471704 152040
rect 467892 152000 471704 152028
rect 467892 151988 467898 152000
rect 471698 151988 471704 152000
rect 471756 151988 471762 152040
rect 485774 151988 485780 152040
rect 485832 152028 485838 152040
rect 490282 152028 490288 152040
rect 485832 152000 490288 152028
rect 485832 151988 485838 152000
rect 490282 151988 490288 152000
rect 490340 151988 490346 152040
rect 516686 151988 516692 152040
rect 516744 152028 516750 152040
rect 520274 152028 520280 152040
rect 516744 152000 520280 152028
rect 516744 151988 516750 152000
rect 520274 151988 520280 152000
rect 520332 151988 520338 152040
rect 413278 151960 413284 151972
rect 405016 151932 413284 151960
rect 413278 151920 413284 151932
rect 413336 151920 413342 151972
rect 417234 151920 417240 151972
rect 417292 151960 417298 151972
rect 431770 151960 431776 151972
rect 417292 151932 431776 151960
rect 417292 151920 417298 151932
rect 431770 151920 431776 151932
rect 431828 151920 431834 151972
rect 431862 151920 431868 151972
rect 431920 151960 431926 151972
rect 439590 151960 439596 151972
rect 431920 151932 439596 151960
rect 431920 151920 431926 151932
rect 439590 151920 439596 151932
rect 439648 151920 439654 151972
rect 440142 151920 440148 151972
rect 440200 151960 440206 151972
rect 440200 151932 444144 151960
rect 440200 151920 440206 151932
rect 26694 151852 26700 151904
rect 26752 151892 26758 151904
rect 71682 151892 71688 151904
rect 26752 151864 71688 151892
rect 26752 151852 26758 151864
rect 71682 151852 71688 151864
rect 71740 151852 71746 151904
rect 109126 151852 109132 151904
rect 109184 151892 109190 151904
rect 109184 151864 110460 151892
rect 109184 151852 109190 151864
rect 33594 151784 33600 151836
rect 33652 151824 33658 151836
rect 82814 151824 82820 151836
rect 33652 151796 82820 151824
rect 33652 151784 33658 151796
rect 82814 151784 82820 151796
rect 82872 151784 82878 151836
rect 105814 151784 105820 151836
rect 105872 151824 105878 151836
rect 110322 151824 110328 151836
rect 105872 151796 110328 151824
rect 105872 151784 105878 151796
rect 110322 151784 110328 151796
rect 110380 151784 110386 151836
rect 110432 151824 110460 151864
rect 110506 151852 110512 151904
rect 110564 151892 110570 151904
rect 138474 151892 138480 151904
rect 110564 151864 138480 151892
rect 110564 151852 110570 151864
rect 138474 151852 138480 151864
rect 138532 151852 138538 151904
rect 139302 151852 139308 151904
rect 139360 151892 139366 151904
rect 203334 151892 203340 151904
rect 139360 151864 203340 151892
rect 139360 151852 139366 151864
rect 203334 151852 203340 151864
rect 203392 151852 203398 151904
rect 260926 151852 260932 151904
rect 260984 151892 260990 151904
rect 316310 151892 316316 151904
rect 260984 151864 316316 151892
rect 260984 151852 260990 151864
rect 316310 151852 316316 151864
rect 316368 151852 316374 151904
rect 321554 151852 321560 151904
rect 321612 151892 321618 151904
rect 362586 151892 362592 151904
rect 321612 151864 362592 151892
rect 321612 151852 321618 151864
rect 362586 151852 362592 151864
rect 362644 151852 362650 151904
rect 363138 151852 363144 151904
rect 363196 151892 363202 151904
rect 364518 151892 364524 151904
rect 363196 151864 364524 151892
rect 363196 151852 363202 151864
rect 364518 151852 364524 151864
rect 364576 151852 364582 151904
rect 386322 151852 386328 151904
rect 386380 151892 386386 151904
rect 394694 151892 394700 151904
rect 386380 151864 394700 151892
rect 386380 151852 386386 151864
rect 394694 151852 394700 151864
rect 394752 151852 394758 151904
rect 396166 151852 396172 151904
rect 396224 151892 396230 151904
rect 402974 151892 402980 151904
rect 396224 151864 402980 151892
rect 396224 151852 396230 151864
rect 402974 151852 402980 151864
rect 403032 151852 403038 151904
rect 404170 151852 404176 151904
rect 404228 151892 404234 151904
rect 404228 151864 408494 151892
rect 404228 151852 404234 151864
rect 128170 151824 128176 151836
rect 110432 151796 128176 151824
rect 128170 151784 128176 151796
rect 128228 151784 128234 151836
rect 129734 151784 129740 151836
rect 129792 151824 129798 151836
rect 146846 151824 146852 151836
rect 129792 151796 146852 151824
rect 129792 151784 129798 151796
rect 146846 151784 146852 151796
rect 146904 151784 146910 151836
rect 146938 151784 146944 151836
rect 146996 151824 147002 151836
rect 157058 151824 157064 151836
rect 146996 151796 157064 151824
rect 146996 151784 147002 151796
rect 157058 151784 157064 151796
rect 157116 151784 157122 151836
rect 169754 151784 169760 151836
rect 169812 151824 169818 151836
rect 185302 151824 185308 151836
rect 169812 151796 185308 151824
rect 169812 151784 169818 151796
rect 185302 151784 185308 151796
rect 185360 151784 185366 151836
rect 283190 151784 283196 151836
rect 283248 151824 283254 151836
rect 287422 151824 287428 151836
rect 283248 151796 287428 151824
rect 283248 151784 283254 151796
rect 287422 151784 287428 151796
rect 287480 151784 287486 151836
rect 299566 151784 299572 151836
rect 299624 151824 299630 151836
rect 346486 151824 346492 151836
rect 299624 151796 342852 151824
rect 299624 151784 299630 151796
rect 342824 151756 342852 151796
rect 344020 151796 346492 151824
rect 344020 151756 344048 151796
rect 346486 151784 346492 151796
rect 346544 151784 346550 151836
rect 349798 151784 349804 151836
rect 349856 151824 349862 151836
rect 380526 151824 380532 151836
rect 349856 151796 380532 151824
rect 349856 151784 349862 151796
rect 380526 151784 380532 151796
rect 380584 151784 380590 151836
rect 398098 151784 398104 151836
rect 398156 151824 398162 151836
rect 405550 151824 405556 151836
rect 398156 151796 405556 151824
rect 398156 151784 398162 151796
rect 405550 151784 405556 151796
rect 405608 151784 405614 151836
rect 408466 151824 408494 151864
rect 413186 151852 413192 151904
rect 413244 151892 413250 151904
rect 413244 151864 415992 151892
rect 413244 151852 413250 151864
rect 415854 151824 415860 151836
rect 408466 151796 415860 151824
rect 415854 151784 415860 151796
rect 415912 151784 415918 151836
rect 415964 151824 415992 151864
rect 418522 151852 418528 151904
rect 418580 151892 418586 151904
rect 426894 151892 426900 151904
rect 418580 151864 426900 151892
rect 418580 151852 418586 151864
rect 426894 151852 426900 151864
rect 426952 151852 426958 151904
rect 437014 151892 437020 151904
rect 427004 151864 437020 151892
rect 421650 151824 421656 151836
rect 415964 151796 421656 151824
rect 421650 151784 421656 151796
rect 421708 151784 421714 151836
rect 421742 151784 421748 151836
rect 421800 151824 421806 151836
rect 427004 151824 427032 151864
rect 437014 151852 437020 151864
rect 437072 151852 437078 151904
rect 437106 151852 437112 151904
rect 437164 151892 437170 151904
rect 443822 151892 443828 151904
rect 437164 151864 443828 151892
rect 437164 151852 437170 151864
rect 443822 151852 443828 151864
rect 443880 151852 443886 151904
rect 444116 151892 444144 151932
rect 444282 151920 444288 151972
rect 444340 151960 444346 151972
rect 451090 151960 451096 151972
rect 444340 151932 451096 151960
rect 444340 151920 444346 151932
rect 451090 151920 451096 151932
rect 451148 151920 451154 151972
rect 451182 151920 451188 151972
rect 451240 151960 451246 151972
rect 457622 151960 457628 151972
rect 451240 151932 457628 151960
rect 451240 151920 451246 151932
rect 457622 151920 457628 151932
rect 457680 151920 457686 151972
rect 469214 151920 469220 151972
rect 469272 151960 469278 151972
rect 472342 151960 472348 151972
rect 469272 151932 472348 151960
rect 469272 151920 469278 151932
rect 472342 151920 472348 151932
rect 472400 151920 472406 151972
rect 487338 151920 487344 151972
rect 487396 151960 487402 151972
rect 490926 151960 490932 151972
rect 487396 151932 490932 151960
rect 487396 151920 487402 151932
rect 490926 151920 490932 151932
rect 490984 151920 490990 151972
rect 509050 151920 509056 151972
rect 509108 151960 509114 151972
rect 510890 151960 510896 151972
rect 509108 151932 510896 151960
rect 509108 151920 509114 151932
rect 510890 151920 510896 151932
rect 510948 151920 510954 151972
rect 515490 151920 515496 151972
rect 515548 151960 515554 151972
rect 518894 151960 518900 151972
rect 515548 151932 518900 151960
rect 515548 151920 515554 151932
rect 518894 151920 518900 151932
rect 518952 151920 518958 151972
rect 444466 151892 444472 151904
rect 444116 151864 444472 151892
rect 444466 151852 444472 151864
rect 444524 151852 444530 151904
rect 451826 151892 451832 151904
rect 444668 151864 451832 151892
rect 421800 151796 427032 151824
rect 421800 151784 421806 151796
rect 427078 151784 427084 151836
rect 427136 151824 427142 151836
rect 431218 151824 431224 151836
rect 427136 151796 431224 151824
rect 427136 151784 427142 151796
rect 431218 151784 431224 151796
rect 431276 151784 431282 151836
rect 431954 151784 431960 151836
rect 432012 151824 432018 151836
rect 441522 151824 441528 151836
rect 432012 151796 441528 151824
rect 432012 151784 432018 151796
rect 441522 151784 441528 151796
rect 441580 151784 441586 151836
rect 441982 151784 441988 151836
rect 442040 151824 442046 151836
rect 444374 151824 444380 151836
rect 442040 151796 444380 151824
rect 442040 151784 442046 151796
rect 444374 151784 444380 151796
rect 444432 151784 444438 151836
rect 342824 151728 344048 151756
rect 441430 151648 441436 151700
rect 441488 151688 441494 151700
rect 444668 151688 444696 151864
rect 451826 151852 451832 151864
rect 451884 151852 451890 151904
rect 464338 151852 464344 151904
rect 464396 151892 464402 151904
rect 467834 151892 467840 151904
rect 464396 151864 467840 151892
rect 464396 151852 464402 151864
rect 467834 151852 467840 151864
rect 467892 151852 467898 151904
rect 467926 151852 467932 151904
rect 467984 151892 467990 151904
rect 471054 151892 471060 151904
rect 467984 151864 471060 151892
rect 467984 151852 467990 151864
rect 471054 151852 471060 151864
rect 471112 151852 471118 151904
rect 488534 151852 488540 151904
rect 488592 151892 488598 151904
rect 492214 151892 492220 151904
rect 488592 151864 492220 151892
rect 488592 151852 488598 151864
rect 492214 151852 492220 151864
rect 492272 151852 492278 151904
rect 507762 151852 507768 151904
rect 507820 151892 507826 151904
rect 509510 151892 509516 151904
rect 507820 151864 509516 151892
rect 507820 151852 507826 151864
rect 509510 151852 509516 151864
rect 509568 151852 509574 151904
rect 516042 151852 516048 151904
rect 516100 151892 516106 151904
rect 519446 151892 519452 151904
rect 516100 151864 519452 151892
rect 516100 151852 516106 151864
rect 519446 151852 519452 151864
rect 519504 151852 519510 151904
rect 445202 151784 445208 151836
rect 445260 151824 445266 151836
rect 446030 151824 446036 151836
rect 445260 151796 446036 151824
rect 445260 151784 445266 151796
rect 446030 151784 446036 151796
rect 446088 151784 446094 151836
rect 488166 151784 488172 151836
rect 488224 151824 488230 151836
rect 491570 151824 491576 151836
rect 488224 151796 491576 151824
rect 488224 151784 488230 151796
rect 491570 151784 491576 151796
rect 491628 151784 491634 151836
rect 499114 151784 499120 151836
rect 499172 151824 499178 151836
rect 499942 151824 499948 151836
rect 499172 151796 499948 151824
rect 499172 151784 499178 151796
rect 499942 151784 499948 151796
rect 500000 151784 500006 151836
rect 517422 151784 517428 151836
rect 517480 151824 517486 151836
rect 521562 151824 521568 151836
rect 517480 151796 521568 151824
rect 517480 151784 517486 151796
rect 521562 151784 521568 151796
rect 521620 151784 521626 151836
rect 441488 151660 444696 151688
rect 441488 151648 441494 151660
rect 82814 151376 82820 151428
rect 82872 151416 82878 151428
rect 117222 151416 117228 151428
rect 82872 151388 117228 151416
rect 82872 151376 82878 151388
rect 117222 151376 117228 151388
rect 117280 151376 117286 151428
rect 68002 151308 68008 151360
rect 68060 151348 68066 151360
rect 112714 151348 112720 151360
rect 68060 151320 112720 151348
rect 68060 151308 68066 151320
rect 112714 151308 112720 151320
rect 112772 151308 112778 151360
rect 71682 151240 71688 151292
rect 71740 151280 71746 151292
rect 117038 151280 117044 151292
rect 71740 151252 117044 151280
rect 71740 151240 71746 151252
rect 117038 151240 117044 151252
rect 117096 151240 117102 151292
rect 64506 151172 64512 151224
rect 64564 151212 64570 151224
rect 112622 151212 112628 151224
rect 64564 151184 112628 151212
rect 64564 151172 64570 151184
rect 112622 151172 112628 151184
rect 112680 151172 112686 151224
rect 61102 151104 61108 151156
rect 61160 151144 61166 151156
rect 112530 151144 112536 151156
rect 61160 151116 112536 151144
rect 61160 151104 61166 151116
rect 112530 151104 112536 151116
rect 112588 151104 112594 151156
rect 57698 151036 57704 151088
rect 57756 151076 57762 151088
rect 111702 151076 111708 151088
rect 57756 151048 111708 151076
rect 57756 151036 57762 151048
rect 111702 151036 111708 151048
rect 111760 151036 111766 151088
rect 54202 150968 54208 151020
rect 54260 151008 54266 151020
rect 112438 151008 112444 151020
rect 54260 150980 112444 151008
rect 54260 150968 54266 150980
rect 112438 150968 112444 150980
rect 112496 150968 112502 151020
rect 50798 150900 50804 150952
rect 50856 150940 50862 150952
rect 111610 150940 111616 150952
rect 50856 150912 111616 150940
rect 50856 150900 50862 150912
rect 111610 150900 111616 150912
rect 111668 150900 111674 150952
rect 47302 150832 47308 150884
rect 47360 150872 47366 150884
rect 111518 150872 111524 150884
rect 47360 150844 111524 150872
rect 47360 150832 47366 150844
rect 111518 150832 111524 150844
rect 111576 150832 111582 150884
rect 43898 150764 43904 150816
rect 43956 150804 43962 150816
rect 111426 150804 111432 150816
rect 43956 150776 111432 150804
rect 43956 150764 43962 150776
rect 111426 150764 111432 150776
rect 111484 150764 111490 150816
rect 40494 150696 40500 150748
rect 40552 150736 40558 150748
rect 111334 150736 111340 150748
rect 40552 150708 111340 150736
rect 40552 150696 40558 150708
rect 111334 150696 111340 150708
rect 111392 150696 111398 150748
rect 36998 150628 37004 150680
rect 37056 150668 37062 150680
rect 111242 150668 111248 150680
rect 37056 150640 111248 150668
rect 37056 150628 37062 150640
rect 111242 150628 111248 150640
rect 111300 150628 111306 150680
rect 23290 150560 23296 150612
rect 23348 150600 23354 150612
rect 116946 150600 116952 150612
rect 23348 150572 116952 150600
rect 23348 150560 23354 150572
rect 116946 150560 116952 150572
rect 117004 150560 117010 150612
rect 12986 150492 12992 150544
rect 13044 150532 13050 150544
rect 116670 150532 116676 150544
rect 13044 150504 116676 150532
rect 13044 150492 13050 150504
rect 116670 150492 116676 150504
rect 116728 150492 116734 150544
rect 2682 150424 2688 150476
rect 2740 150464 2746 150476
rect 111058 150464 111064 150476
rect 2740 150436 111064 150464
rect 2740 150424 2746 150436
rect 111058 150424 111064 150436
rect 111116 150424 111122 150476
rect 263686 150288 263692 150340
rect 263744 150328 263750 150340
rect 263744 150300 264422 150328
rect 263744 150288 263750 150300
rect 264394 150204 264422 150300
rect 122834 150152 122840 150204
rect 122892 150192 122898 150204
rect 123708 150192 123714 150204
rect 122892 150164 123714 150192
rect 122892 150152 122898 150164
rect 123708 150152 123714 150164
rect 123766 150152 123772 150204
rect 146386 150152 146392 150204
rect 146444 150192 146450 150204
rect 147536 150192 147542 150204
rect 146444 150164 147542 150192
rect 146444 150152 146450 150164
rect 147536 150152 147542 150164
rect 147594 150152 147600 150204
rect 164326 150152 164332 150204
rect 164384 150192 164390 150204
rect 165476 150192 165482 150204
rect 164384 150164 165482 150192
rect 164384 150152 164390 150164
rect 165476 150152 165482 150164
rect 165534 150152 165540 150204
rect 168374 150152 168380 150204
rect 168432 150192 168438 150204
rect 169340 150192 169346 150204
rect 168432 150164 169346 150192
rect 168432 150152 168438 150164
rect 169340 150152 169346 150164
rect 169398 150152 169404 150204
rect 171134 150152 171140 150204
rect 171192 150192 171198 150204
rect 171916 150192 171922 150204
rect 171192 150164 171922 150192
rect 171192 150152 171198 150164
rect 171916 150152 171922 150164
rect 171974 150152 171980 150204
rect 172698 150152 172704 150204
rect 172756 150192 172762 150204
rect 173848 150192 173854 150204
rect 172756 150164 173854 150192
rect 172756 150152 172762 150164
rect 173848 150152 173854 150164
rect 173906 150152 173912 150204
rect 182266 150152 182272 150204
rect 182324 150192 182330 150204
rect 183416 150192 183422 150204
rect 182324 150164 183422 150192
rect 182324 150152 182330 150164
rect 183416 150152 183422 150164
rect 183474 150152 183480 150204
rect 211246 150152 211252 150204
rect 211304 150192 211310 150204
rect 212304 150192 212310 150204
rect 211304 150164 212310 150192
rect 211304 150152 211310 150164
rect 212304 150152 212310 150164
rect 212362 150152 212368 150204
rect 225046 150152 225052 150204
rect 225104 150192 225110 150204
rect 225828 150192 225834 150204
rect 225104 150164 225834 150192
rect 225104 150152 225110 150164
rect 225828 150152 225834 150164
rect 225886 150152 225892 150204
rect 229186 150152 229192 150204
rect 229244 150192 229250 150204
rect 230336 150192 230342 150204
rect 229244 150164 230342 150192
rect 229244 150152 229250 150164
rect 230336 150152 230342 150164
rect 230394 150152 230400 150204
rect 233234 150152 233240 150204
rect 233292 150192 233298 150204
rect 234200 150192 234206 150204
rect 233292 150164 234206 150192
rect 233292 150152 233298 150164
rect 234200 150152 234206 150164
rect 234258 150152 234264 150204
rect 238938 150152 238944 150204
rect 238996 150192 239002 150204
rect 239996 150192 240002 150204
rect 238996 150164 240002 150192
rect 238996 150152 239002 150164
rect 239996 150152 240002 150164
rect 240054 150152 240060 150204
rect 253934 150152 253940 150204
rect 253992 150192 253998 150204
rect 254716 150192 254722 150204
rect 253992 150164 254722 150192
rect 253992 150152 253998 150164
rect 254716 150152 254722 150164
rect 254774 150152 254780 150204
rect 256786 150152 256792 150204
rect 256844 150192 256850 150204
rect 257936 150192 257942 150204
rect 256844 150164 257942 150192
rect 256844 150152 256850 150164
rect 257936 150152 257942 150164
rect 257994 150152 258000 150204
rect 264376 150152 264382 150204
rect 264434 150152 264440 150204
rect 269114 150152 269120 150204
rect 269172 150192 269178 150204
rect 270172 150192 270178 150204
rect 269172 150164 270178 150192
rect 269172 150152 269178 150164
rect 270172 150152 270178 150164
rect 270230 150152 270236 150204
rect 281534 150152 281540 150204
rect 281592 150192 281598 150204
rect 282316 150192 282322 150204
rect 281592 150164 282322 150192
rect 281592 150152 281598 150164
rect 282316 150152 282322 150164
rect 282374 150152 282380 150204
rect 283098 150152 283104 150204
rect 283156 150192 283162 150204
rect 284248 150192 284254 150204
rect 283156 150164 284254 150192
rect 283156 150152 283162 150164
rect 284248 150152 284254 150164
rect 284306 150152 284312 150204
rect 284386 150152 284392 150204
rect 284444 150192 284450 150204
rect 285536 150192 285542 150204
rect 284444 150164 285542 150192
rect 284444 150152 284450 150164
rect 285536 150152 285542 150164
rect 285594 150152 285600 150204
rect 299474 150152 299480 150204
rect 299532 150192 299538 150204
rect 300348 150192 300354 150204
rect 299532 150164 300354 150192
rect 299532 150152 299538 150164
rect 300348 150152 300354 150164
rect 300406 150152 300412 150204
rect 321738 150152 321744 150204
rect 321796 150192 321802 150204
rect 322796 150192 322802 150204
rect 321796 150164 322802 150192
rect 321796 150152 321802 150164
rect 322796 150152 322802 150164
rect 322854 150152 322860 150204
rect 328454 150152 328460 150204
rect 328512 150192 328518 150204
rect 329236 150192 329242 150204
rect 328512 150164 329242 150192
rect 328512 150152 328518 150164
rect 329236 150152 329242 150164
rect 329294 150152 329300 150204
rect 332686 150152 332692 150204
rect 332744 150192 332750 150204
rect 333744 150192 333750 150204
rect 332744 150164 333750 150192
rect 332744 150152 332750 150164
rect 333744 150152 333750 150164
rect 333802 150152 333808 150204
rect 338390 150152 338396 150204
rect 338448 150192 338454 150204
rect 339448 150192 339454 150204
rect 338448 150164 339454 150192
rect 338448 150152 338454 150164
rect 339448 150152 339454 150164
rect 339506 150152 339512 150204
rect 345106 150152 345112 150204
rect 345164 150192 345170 150204
rect 345888 150192 345894 150204
rect 345164 150164 345894 150192
rect 345164 150152 345170 150164
rect 345888 150152 345894 150164
rect 345946 150152 345952 150204
rect 358906 150152 358912 150204
rect 358964 150192 358970 150204
rect 360056 150192 360062 150204
rect 358964 150164 360062 150192
rect 358964 150152 358970 150164
rect 360056 150152 360062 150164
rect 360114 150152 360120 150204
rect 362954 150152 362960 150204
rect 363012 150192 363018 150204
rect 363920 150192 363926 150204
rect 363012 150164 363926 150192
rect 363012 150152 363018 150164
rect 363920 150152 363926 150164
rect 363978 150152 363984 150204
rect 375558 150152 375564 150204
rect 375616 150192 375622 150204
rect 376708 150192 376714 150204
rect 375616 150164 376714 150192
rect 375616 150152 375622 150164
rect 376708 150152 376714 150164
rect 376766 150152 376772 150204
rect 378134 150152 378140 150204
rect 378192 150192 378198 150204
rect 379284 150192 379290 150204
rect 378192 150164 379290 150192
rect 378192 150152 378198 150164
rect 379284 150152 379290 150164
rect 379342 150152 379348 150204
rect 394970 150152 394976 150204
rect 395028 150192 395034 150204
rect 396028 150192 396034 150204
rect 395028 150164 396034 150192
rect 395028 150152 395034 150164
rect 396028 150152 396034 150164
rect 396086 150152 396092 150204
rect 462314 150152 462320 150204
rect 462372 150192 462378 150204
rect 463372 150192 463378 150204
rect 462372 150164 463378 150192
rect 462372 150152 462378 150164
rect 463372 150152 463378 150164
rect 463430 150152 463436 150204
rect 477678 150152 477684 150204
rect 477736 150192 477742 150204
rect 478828 150192 478834 150204
rect 477736 150164 478834 150192
rect 477736 150152 477742 150164
rect 478828 150152 478834 150164
rect 478886 150152 478892 150204
rect 478966 150152 478972 150204
rect 479024 150192 479030 150204
rect 480116 150192 480122 150204
rect 479024 150164 480122 150192
rect 479024 150152 479030 150164
rect 480116 150152 480122 150164
rect 480174 150152 480180 150204
rect 481634 150152 481640 150204
rect 481692 150192 481698 150204
rect 482692 150192 482698 150204
rect 481692 150164 482698 150192
rect 481692 150152 481698 150164
rect 482692 150152 482698 150164
rect 482750 150152 482756 150204
rect 483198 150152 483204 150204
rect 483256 150192 483262 150204
rect 483980 150192 483986 150204
rect 483256 150164 483986 150192
rect 483256 150152 483262 150164
rect 483980 150152 483986 150164
rect 484038 150152 484044 150204
rect 518020 150152 518026 150204
rect 518078 150192 518084 150204
rect 518802 150192 518808 150204
rect 518078 150164 518808 150192
rect 518078 150152 518084 150164
rect 518802 150152 518808 150164
rect 518860 150152 518866 150204
rect 102594 150016 102600 150068
rect 102652 150056 102658 150068
rect 116210 150056 116216 150068
rect 102652 150028 116216 150056
rect 102652 150016 102658 150028
rect 116210 150016 116216 150028
rect 116268 150016 116274 150068
rect 20162 149948 20168 150000
rect 20220 149988 20226 150000
rect 116854 149988 116860 150000
rect 20220 149960 116860 149988
rect 20220 149948 20226 149960
rect 116854 149948 116860 149960
rect 116912 149948 116918 150000
rect 16482 149880 16488 149932
rect 16540 149920 16546 149932
rect 116762 149920 116768 149932
rect 16540 149892 116768 149920
rect 16540 149880 16546 149892
rect 116762 149880 116768 149892
rect 116820 149880 116826 149932
rect 9582 149812 9588 149864
rect 9640 149852 9646 149864
rect 116578 149852 116584 149864
rect 9640 149824 116584 149852
rect 9640 149812 9646 149824
rect 116578 149812 116584 149824
rect 116636 149812 116642 149864
rect 6362 149744 6368 149796
rect 6420 149784 6426 149796
rect 111150 149784 111156 149796
rect 6420 149756 111156 149784
rect 6420 149744 6426 149756
rect 111150 149744 111156 149756
rect 111208 149744 111214 149796
rect 85482 149676 85488 149728
rect 85540 149716 85546 149728
rect 112346 149716 112352 149728
rect 85540 149688 112352 149716
rect 85540 149676 85546 149688
rect 112346 149676 112352 149688
rect 112404 149676 112410 149728
rect 81986 149608 81992 149660
rect 82044 149648 82050 149660
rect 113082 149648 113088 149660
rect 82044 149620 113088 149648
rect 82044 149608 82050 149620
rect 113082 149608 113088 149620
rect 113140 149608 113146 149660
rect 78582 149540 78588 149592
rect 78640 149580 78646 149592
rect 112990 149580 112996 149592
rect 78640 149552 112996 149580
rect 78640 149540 78646 149552
rect 112990 149540 112996 149552
rect 113048 149540 113054 149592
rect 75178 149472 75184 149524
rect 75236 149512 75242 149524
rect 112898 149512 112904 149524
rect 75236 149484 112904 149512
rect 75236 149472 75242 149484
rect 112898 149472 112904 149484
rect 112956 149472 112962 149524
rect 71682 149404 71688 149456
rect 71740 149444 71746 149456
rect 112806 149444 112812 149456
rect 71740 149416 112812 149444
rect 71740 149404 71746 149416
rect 112806 149404 112812 149416
rect 112864 149404 112870 149456
rect 30282 149336 30288 149388
rect 30340 149376 30346 149388
rect 117130 149376 117136 149388
rect 30340 149348 117136 149376
rect 30340 149336 30346 149348
rect 117130 149336 117136 149348
rect 117188 149336 117194 149388
rect 88978 149268 88984 149320
rect 89036 149308 89042 149320
rect 89036 149280 93854 149308
rect 89036 149268 89042 149280
rect 92014 149200 92020 149252
rect 92072 149200 92078 149252
rect 92032 149104 92060 149200
rect 93826 149172 93854 149280
rect 95786 149268 95792 149320
rect 95844 149268 95850 149320
rect 99282 149268 99288 149320
rect 99340 149308 99346 149320
rect 116026 149308 116032 149320
rect 99340 149280 116032 149308
rect 99340 149268 99346 149280
rect 116026 149268 116032 149280
rect 116084 149268 116090 149320
rect 95804 149240 95832 149268
rect 116394 149240 116400 149252
rect 95804 149212 116400 149240
rect 116394 149200 116400 149212
rect 116452 149200 116458 149252
rect 116486 149172 116492 149184
rect 93826 149144 116492 149172
rect 116486 149132 116492 149144
rect 116544 149132 116550 149184
rect 112254 149104 112260 149116
rect 92032 149076 112260 149104
rect 112254 149064 112260 149076
rect 112312 149064 112318 149116
rect 109586 148996 109592 149048
rect 109644 149036 109650 149048
rect 116118 149036 116124 149048
rect 109644 149008 116124 149036
rect 109644 148996 109650 149008
rect 116118 148996 116124 149008
rect 116176 148996 116182 149048
rect 110322 147568 110328 147620
rect 110380 147608 110386 147620
rect 116118 147608 116124 147620
rect 110380 147580 116124 147608
rect 110380 147568 110386 147580
rect 116118 147568 116124 147580
rect 116176 147568 116182 147620
rect 112254 140700 112260 140752
rect 112312 140740 112318 140752
rect 116118 140740 116124 140752
rect 112312 140712 116124 140740
rect 112312 140700 112318 140712
rect 116118 140700 116124 140712
rect 116176 140700 116182 140752
rect 112346 136552 112352 136604
rect 112404 136592 112410 136604
rect 116118 136592 116124 136604
rect 112404 136564 116124 136592
rect 112404 136552 112410 136564
rect 116118 136552 116124 136564
rect 116176 136552 116182 136604
rect 113082 133832 113088 133884
rect 113140 133872 113146 133884
rect 116026 133872 116032 133884
rect 113140 133844 116032 133872
rect 113140 133832 113146 133844
rect 116026 133832 116032 133844
rect 116084 133832 116090 133884
rect 114186 132608 114192 132660
rect 114244 132648 114250 132660
rect 115198 132648 115204 132660
rect 114244 132620 115204 132648
rect 114244 132608 114250 132620
rect 115198 132608 115204 132620
rect 115256 132608 115262 132660
rect 112990 132404 112996 132456
rect 113048 132444 113054 132456
rect 116118 132444 116124 132456
rect 113048 132416 116124 132444
rect 113048 132404 113054 132416
rect 116118 132404 116124 132416
rect 116176 132404 116182 132456
rect 112898 131044 112904 131096
rect 112956 131084 112962 131096
rect 116118 131084 116124 131096
rect 112956 131056 116124 131084
rect 112956 131044 112962 131056
rect 116118 131044 116124 131056
rect 116176 131044 116182 131096
rect 112806 128256 112812 128308
rect 112864 128296 112870 128308
rect 116118 128296 116124 128308
rect 112864 128268 116124 128296
rect 112864 128256 112870 128268
rect 116118 128256 116124 128268
rect 116176 128256 116182 128308
rect 112714 126896 112720 126948
rect 112772 126936 112778 126948
rect 116026 126936 116032 126948
rect 112772 126908 116032 126936
rect 112772 126896 112778 126908
rect 116026 126896 116032 126908
rect 116084 126896 116090 126948
rect 112622 124108 112628 124160
rect 112680 124148 112686 124160
rect 116118 124148 116124 124160
rect 112680 124120 116124 124148
rect 112680 124108 112686 124120
rect 116118 124108 116124 124120
rect 116176 124108 116182 124160
rect 112530 122748 112536 122800
rect 112588 122788 112594 122800
rect 115934 122788 115940 122800
rect 112588 122760 115940 122788
rect 112588 122748 112594 122760
rect 115934 122748 115940 122760
rect 115992 122748 115998 122800
rect 111702 121388 111708 121440
rect 111760 121428 111766 121440
rect 116118 121428 116124 121440
rect 111760 121400 116124 121428
rect 111760 121388 111766 121400
rect 116118 121388 116124 121400
rect 116176 121388 116182 121440
rect 112438 118600 112444 118652
rect 112496 118640 112502 118652
rect 116118 118640 116124 118652
rect 112496 118612 116124 118640
rect 112496 118600 112502 118612
rect 116118 118600 116124 118612
rect 116176 118600 116182 118652
rect 116486 117988 116492 118040
rect 116544 118028 116550 118040
rect 117222 118028 117228 118040
rect 116544 118000 117228 118028
rect 116544 117988 116550 118000
rect 117222 117988 117228 118000
rect 117280 117988 117286 118040
rect 111610 117240 111616 117292
rect 111668 117280 111674 117292
rect 116118 117280 116124 117292
rect 111668 117252 116124 117280
rect 111668 117240 111674 117252
rect 116118 117240 116124 117252
rect 116176 117240 116182 117292
rect 111518 114452 111524 114504
rect 111576 114492 111582 114504
rect 116118 114492 116124 114504
rect 111576 114464 116124 114492
rect 111576 114452 111582 114464
rect 116118 114452 116124 114464
rect 116176 114452 116182 114504
rect 111426 113092 111432 113144
rect 111484 113132 111490 113144
rect 115934 113132 115940 113144
rect 111484 113104 115940 113132
rect 111484 113092 111490 113104
rect 115934 113092 115940 113104
rect 115992 113092 115998 113144
rect 111334 111732 111340 111784
rect 111392 111772 111398 111784
rect 116118 111772 116124 111784
rect 111392 111744 116124 111772
rect 111392 111732 111398 111744
rect 116118 111732 116124 111744
rect 116176 111732 116182 111784
rect 111242 108944 111248 108996
rect 111300 108984 111306 108996
rect 116118 108984 116124 108996
rect 111300 108956 116124 108984
rect 111300 108944 111306 108956
rect 116118 108944 116124 108956
rect 116176 108944 116182 108996
rect 111150 92420 111156 92472
rect 111208 92460 111214 92472
rect 116118 92460 116124 92472
rect 111208 92432 116124 92460
rect 111208 92420 111214 92432
rect 116118 92420 116124 92432
rect 116176 92420 116182 92472
rect 111058 89632 111064 89684
rect 111116 89672 111122 89684
rect 116118 89672 116124 89684
rect 111116 89644 116124 89672
rect 111116 89632 111122 89644
rect 116118 89632 116124 89644
rect 116176 89632 116182 89684
rect 113818 88272 113824 88324
rect 113876 88312 113882 88324
rect 116026 88312 116032 88324
rect 113876 88284 116032 88312
rect 113876 88272 113882 88284
rect 116026 88272 116032 88284
rect 116084 88272 116090 88324
rect 114462 87184 114468 87236
rect 114520 87224 114526 87236
rect 116486 87224 116492 87236
rect 114520 87196 116492 87224
rect 114520 87184 114526 87196
rect 116486 87184 116492 87196
rect 116544 87184 116550 87236
rect 113910 83920 113916 83972
rect 113968 83960 113974 83972
rect 116578 83960 116584 83972
rect 113968 83932 116584 83960
rect 113968 83920 113974 83932
rect 116578 83920 116584 83932
rect 116636 83920 116642 83972
rect 114002 82764 114008 82816
rect 114060 82804 114066 82816
rect 116210 82804 116216 82816
rect 114060 82776 116216 82804
rect 114060 82764 114066 82776
rect 116210 82764 116216 82776
rect 116268 82764 116274 82816
rect 114094 79976 114100 80028
rect 114152 80016 114158 80028
rect 115934 80016 115940 80028
rect 114152 79988 115940 80016
rect 114152 79976 114158 79988
rect 115934 79976 115940 79988
rect 115992 79976 115998 80028
rect 114186 71748 114192 71800
rect 114244 71788 114250 71800
rect 116578 71788 116584 71800
rect 114244 71760 116584 71788
rect 114244 71748 114250 71760
rect 116578 71748 116584 71760
rect 116636 71748 116642 71800
rect 114094 69028 114100 69080
rect 114152 69068 114158 69080
rect 116302 69068 116308 69080
rect 114152 69040 116308 69068
rect 114152 69028 114158 69040
rect 116302 69028 116308 69040
rect 116360 69028 116366 69080
rect 114002 67600 114008 67652
rect 114060 67640 114066 67652
rect 116118 67640 116124 67652
rect 114060 67612 116124 67640
rect 114060 67600 114066 67612
rect 116118 67600 116124 67612
rect 116176 67600 116182 67652
rect 113910 66240 113916 66292
rect 113968 66280 113974 66292
rect 116578 66280 116584 66292
rect 113968 66252 116584 66280
rect 113968 66240 113974 66252
rect 116578 66240 116584 66252
rect 116636 66240 116642 66292
rect 114462 64540 114468 64592
rect 114520 64580 114526 64592
rect 116578 64580 116584 64592
rect 114520 64552 116584 64580
rect 114520 64540 114526 64552
rect 116578 64540 116584 64552
rect 116636 64540 116642 64592
rect 113818 63520 113824 63572
rect 113876 63560 113882 63572
rect 116210 63560 116216 63572
rect 113876 63532 116216 63560
rect 113876 63520 113882 63532
rect 116210 63520 116216 63532
rect 116268 63520 116274 63572
rect 109678 41420 109684 41472
rect 109736 41460 109742 41472
rect 116118 41460 116124 41472
rect 109736 41432 116124 41460
rect 109736 41420 109742 41432
rect 116118 41420 116124 41432
rect 116176 41420 116182 41472
rect 114094 38632 114100 38684
rect 114152 38672 114158 38684
rect 116394 38672 116400 38684
rect 114152 38644 116400 38672
rect 114152 38632 114158 38644
rect 116394 38632 116400 38644
rect 116452 38632 116458 38684
rect 116210 38496 116216 38548
rect 116268 38536 116274 38548
rect 116394 38536 116400 38548
rect 116268 38508 116400 38536
rect 116268 38496 116274 38508
rect 116394 38496 116400 38508
rect 116452 38496 116458 38548
rect 114186 37272 114192 37324
rect 114244 37312 114250 37324
rect 116210 37312 116216 37324
rect 114244 37284 116216 37312
rect 114244 37272 114250 37284
rect 116210 37272 116216 37284
rect 116268 37272 116274 37324
rect 111058 34484 111064 34536
rect 111116 34524 111122 34536
rect 116118 34524 116124 34536
rect 111116 34496 116124 34524
rect 111116 34484 111122 34496
rect 116118 34484 116124 34496
rect 116176 34484 116182 34536
rect 112438 33124 112444 33176
rect 112496 33164 112502 33176
rect 116118 33164 116124 33176
rect 112496 33136 116124 33164
rect 112496 33124 112502 33136
rect 116118 33124 116124 33136
rect 116176 33124 116182 33176
rect 112530 31764 112536 31816
rect 112588 31804 112594 31816
rect 116118 31804 116124 31816
rect 112588 31776 116124 31804
rect 112588 31764 112594 31776
rect 116118 31764 116124 31776
rect 116176 31764 116182 31816
rect 112622 28976 112628 29028
rect 112680 29016 112686 29028
rect 116118 29016 116124 29028
rect 112680 28988 116124 29016
rect 112680 28976 112686 28988
rect 116118 28976 116124 28988
rect 116176 28976 116182 29028
rect 112714 27616 112720 27668
rect 112772 27656 112778 27668
rect 116118 27656 116124 27668
rect 112772 27628 116124 27656
rect 112772 27616 112778 27628
rect 116118 27616 116124 27628
rect 116176 27616 116182 27668
rect 112806 24828 112812 24880
rect 112864 24868 112870 24880
rect 116118 24868 116124 24880
rect 112864 24840 116124 24868
rect 112864 24828 112870 24840
rect 116118 24828 116124 24840
rect 116176 24828 116182 24880
rect 111150 23468 111156 23520
rect 111208 23508 111214 23520
rect 116118 23508 116124 23520
rect 111208 23480 116124 23508
rect 111208 23468 111214 23480
rect 116118 23468 116124 23480
rect 116176 23468 116182 23520
rect 111242 22108 111248 22160
rect 111300 22148 111306 22160
rect 116026 22148 116032 22160
rect 111300 22120 116032 22148
rect 111300 22108 111306 22120
rect 116026 22108 116032 22120
rect 116084 22108 116090 22160
rect 116026 16464 116032 16516
rect 116084 16504 116090 16516
rect 116210 16504 116216 16516
rect 116084 16476 116216 16504
rect 116084 16464 116090 16476
rect 116210 16464 116216 16476
rect 116268 16464 116274 16516
rect 116210 11840 116216 11892
rect 116268 11840 116274 11892
rect 116228 11676 116256 11840
rect 116302 11676 116308 11688
rect 116228 11648 116308 11676
rect 116302 11636 116308 11648
rect 116360 11636 116366 11688
rect 116946 11364 116952 11416
rect 117004 11404 117010 11416
rect 117314 11404 117320 11416
rect 117004 11376 117320 11404
rect 117004 11364 117010 11376
rect 117314 11364 117320 11376
rect 117372 11364 117378 11416
rect 116946 5448 116952 5500
rect 117004 5488 117010 5500
rect 117130 5488 117136 5500
rect 117004 5460 117136 5488
rect 117004 5448 117010 5460
rect 117130 5448 117136 5460
rect 117188 5448 117194 5500
rect 116302 5312 116308 5364
rect 116360 5352 116366 5364
rect 116946 5352 116952 5364
rect 116360 5324 116952 5352
rect 116360 5312 116366 5324
rect 116946 5312 116952 5324
rect 117004 5312 117010 5364
rect 115934 5176 115940 5228
rect 115992 5216 115998 5228
rect 116302 5216 116308 5228
rect 115992 5188 116308 5216
rect 115992 5176 115998 5188
rect 116302 5176 116308 5188
rect 116360 5176 116366 5228
rect 115934 5040 115940 5092
rect 115992 5080 115998 5092
rect 116118 5080 116124 5092
rect 115992 5052 116124 5080
rect 115992 5040 115998 5052
rect 116118 5040 116124 5052
rect 116176 5040 116182 5092
rect 109770 4156 109776 4208
rect 109828 4196 109834 4208
rect 116118 4196 116124 4208
rect 109828 4168 116124 4196
rect 109828 4156 109834 4168
rect 116118 4156 116124 4168
rect 116176 4156 116182 4208
rect 111058 3924 111064 3936
rect 63466 3896 77524 3924
rect 39408 3624 58848 3652
rect 27586 3148 35894 3176
rect 27586 3040 27614 3148
rect 26206 3012 27614 3040
rect 26206 2904 26234 3012
rect 2516 2876 26234 2904
rect 2516 2644 2544 2876
rect 2498 2592 2504 2644
rect 2556 2592 2562 2644
rect 35866 2564 35894 3148
rect 39408 2644 39436 3624
rect 44146 3556 52316 3584
rect 44146 3380 44174 3556
rect 39776 3352 44174 3380
rect 39776 2644 39804 3352
rect 43088 3284 51764 3312
rect 39390 2592 39396 2644
rect 39448 2592 39454 2644
rect 39758 2592 39764 2644
rect 39816 2592 39822 2644
rect 42978 2592 42984 2644
rect 43036 2632 43042 2644
rect 43088 2632 43116 3284
rect 43548 3216 47072 3244
rect 43548 2644 43576 3216
rect 47044 3176 47072 3216
rect 46124 3148 46934 3176
rect 47044 3148 47164 3176
rect 46124 2644 46152 3148
rect 43036 2604 43116 2632
rect 43036 2592 43042 2604
rect 43530 2592 43536 2644
rect 43588 2592 43594 2644
rect 46106 2592 46112 2644
rect 46164 2592 46170 2644
rect 46906 2632 46934 3148
rect 47136 2768 47164 3148
rect 51736 2972 51764 3284
rect 52288 3108 52316 3556
rect 52426 3148 58756 3176
rect 52426 3108 52454 3148
rect 52288 3080 52454 3108
rect 51736 2944 52592 2972
rect 52564 2768 52592 2944
rect 47136 2740 52454 2768
rect 52564 2740 53788 2768
rect 50614 2632 50620 2644
rect 46906 2604 50620 2632
rect 50614 2592 50620 2604
rect 50672 2592 50678 2644
rect 52426 2632 52454 2740
rect 53650 2632 53656 2644
rect 52426 2604 53656 2632
rect 53650 2592 53656 2604
rect 53708 2592 53714 2644
rect 53760 2564 53788 2740
rect 58728 2644 58756 3148
rect 58820 2644 58848 3624
rect 63466 3584 63494 3896
rect 77496 3856 77524 3896
rect 78600 3896 111064 3924
rect 78600 3856 78628 3896
rect 111058 3884 111064 3896
rect 111116 3884 111122 3936
rect 112438 3856 112444 3868
rect 77496 3828 77984 3856
rect 77956 3788 77984 3828
rect 78048 3828 78628 3856
rect 79244 3828 112444 3856
rect 78048 3788 78076 3828
rect 77956 3760 78076 3788
rect 79244 3584 79272 3828
rect 112438 3816 112444 3828
rect 112496 3816 112502 3868
rect 112530 3788 112536 3800
rect 62868 3556 63494 3584
rect 77266 3556 79272 3584
rect 81544 3760 112536 3788
rect 62868 2644 62896 3556
rect 62960 3284 75914 3312
rect 58710 2592 58716 2644
rect 58768 2592 58774 2644
rect 58802 2592 58808 2644
rect 58860 2592 58866 2644
rect 62850 2592 62856 2644
rect 62908 2592 62914 2644
rect 58618 2564 58624 2576
rect 35866 2536 46934 2564
rect 53760 2536 58624 2564
rect 32766 2456 32772 2508
rect 32824 2496 32830 2508
rect 43530 2496 43536 2508
rect 32824 2468 43536 2496
rect 32824 2456 32830 2468
rect 43530 2456 43536 2468
rect 43588 2456 43594 2508
rect 46906 2496 46934 2536
rect 58618 2524 58624 2536
rect 58676 2524 58682 2576
rect 59722 2524 59728 2576
rect 59780 2564 59786 2576
rect 62960 2564 62988 3284
rect 75886 3244 75914 3284
rect 77266 3244 77294 3556
rect 71700 3216 74534 3244
rect 75886 3216 77294 3244
rect 71700 2972 71728 3216
rect 74506 3176 74534 3216
rect 74506 3148 77294 3176
rect 77266 3108 77294 3148
rect 77266 3080 79456 3108
rect 63328 2944 71728 2972
rect 79428 2972 79456 3080
rect 79428 2944 80468 2972
rect 63328 2644 63356 2944
rect 76944 2876 77294 2904
rect 76944 2836 76972 2876
rect 63512 2808 76972 2836
rect 77266 2836 77294 2876
rect 77266 2808 80376 2836
rect 63512 2644 63540 2808
rect 67008 2672 80284 2700
rect 67008 2644 67036 2672
rect 80256 2644 80284 2672
rect 80348 2644 80376 2808
rect 80440 2644 80468 2944
rect 81544 2644 81572 3760
rect 112530 3748 112536 3760
rect 112588 3748 112594 3800
rect 112622 3720 112628 3732
rect 81636 3692 112628 3720
rect 81636 2644 81664 3692
rect 112622 3680 112628 3692
rect 112680 3680 112686 3732
rect 112714 3652 112720 3664
rect 81820 3624 112720 3652
rect 81820 2644 81848 3624
rect 112714 3612 112720 3624
rect 112772 3612 112778 3664
rect 112806 3584 112812 3596
rect 81912 3556 112812 3584
rect 81912 2644 81940 3556
rect 112806 3544 112812 3556
rect 112864 3544 112870 3596
rect 111150 3516 111156 3528
rect 82004 3488 111156 3516
rect 82004 2644 82032 3488
rect 111150 3476 111156 3488
rect 111208 3476 111214 3528
rect 111242 3448 111248 3460
rect 82648 3420 111248 3448
rect 63310 2592 63316 2644
rect 63368 2592 63374 2644
rect 63494 2592 63500 2644
rect 63552 2592 63558 2644
rect 66990 2592 66996 2644
rect 67048 2592 67054 2644
rect 68002 2592 68008 2644
rect 68060 2632 68066 2644
rect 80146 2632 80152 2644
rect 68060 2604 80152 2632
rect 68060 2592 68066 2604
rect 80146 2592 80152 2604
rect 80204 2592 80210 2644
rect 80238 2592 80244 2644
rect 80296 2592 80302 2644
rect 80330 2592 80336 2644
rect 80388 2592 80394 2644
rect 80422 2592 80428 2644
rect 80480 2592 80486 2644
rect 81526 2592 81532 2644
rect 81584 2592 81590 2644
rect 81618 2592 81624 2644
rect 81676 2592 81682 2644
rect 81802 2592 81808 2644
rect 81860 2592 81866 2644
rect 81894 2592 81900 2644
rect 81952 2592 81958 2644
rect 81986 2592 81992 2644
rect 82044 2592 82050 2644
rect 82446 2592 82452 2644
rect 82504 2632 82510 2644
rect 82648 2632 82676 3420
rect 111242 3408 111248 3420
rect 111300 3408 111306 3460
rect 114186 3380 114192 3392
rect 82740 3352 114192 3380
rect 82740 2644 82768 3352
rect 114186 3340 114192 3352
rect 114244 3340 114250 3392
rect 114094 3312 114100 3324
rect 86926 3284 89714 3312
rect 86926 3040 86954 3284
rect 89686 3244 89714 3284
rect 91066 3284 114100 3312
rect 91066 3244 91094 3284
rect 114094 3272 114100 3284
rect 114152 3272 114158 3324
rect 112438 3244 112444 3256
rect 89686 3216 91094 3244
rect 107626 3216 112444 3244
rect 107626 3176 107654 3216
rect 112438 3204 112444 3216
rect 112496 3204 112502 3256
rect 99346 3148 107654 3176
rect 99346 3108 99374 3148
rect 82924 3012 86954 3040
rect 89686 3080 99374 3108
rect 82504 2604 82676 2632
rect 82504 2592 82510 2604
rect 82722 2592 82728 2644
rect 82780 2592 82786 2644
rect 59780 2536 62988 2564
rect 59780 2524 59786 2536
rect 73246 2524 73252 2576
rect 73304 2564 73310 2576
rect 82354 2564 82360 2576
rect 73304 2536 82360 2564
rect 73304 2524 73310 2536
rect 82354 2524 82360 2536
rect 82412 2524 82418 2576
rect 73062 2496 73068 2508
rect 46906 2468 73068 2496
rect 73062 2456 73068 2468
rect 73120 2456 73126 2508
rect 73338 2456 73344 2508
rect 73396 2496 73402 2508
rect 82262 2496 82268 2508
rect 73396 2468 82268 2496
rect 73396 2456 73402 2468
rect 82262 2456 82268 2468
rect 82320 2456 82326 2508
rect 36354 2388 36360 2440
rect 36412 2428 36418 2440
rect 39758 2428 39764 2440
rect 36412 2400 39764 2428
rect 36412 2388 36418 2400
rect 39758 2388 39764 2400
rect 39816 2388 39822 2440
rect 50614 2388 50620 2440
rect 50672 2428 50678 2440
rect 56134 2428 56140 2440
rect 50672 2400 56140 2428
rect 50672 2388 50678 2400
rect 56134 2388 56140 2400
rect 56192 2388 56198 2440
rect 58618 2388 58624 2440
rect 58676 2428 58682 2440
rect 68002 2428 68008 2440
rect 58676 2400 68008 2428
rect 58676 2388 58682 2400
rect 68002 2388 68008 2400
rect 68060 2388 68066 2440
rect 80146 2388 80152 2440
rect 80204 2428 80210 2440
rect 81894 2428 81900 2440
rect 80204 2400 81900 2428
rect 80204 2388 80210 2400
rect 81894 2388 81900 2400
rect 81952 2388 81958 2440
rect 82924 2428 82952 3012
rect 89686 2972 89714 3080
rect 117958 3040 117964 3052
rect 83016 2944 89714 2972
rect 100588 3012 107654 3040
rect 83016 2644 83044 2944
rect 83108 2876 98040 2904
rect 83108 2644 83136 2876
rect 86926 2808 96614 2836
rect 82998 2592 83004 2644
rect 83056 2592 83062 2644
rect 83090 2592 83096 2644
rect 83148 2592 83154 2644
rect 82096 2400 82952 2428
rect 52914 2320 52920 2372
rect 52972 2360 52978 2372
rect 66990 2360 66996 2372
rect 52972 2332 66996 2360
rect 52972 2320 52978 2332
rect 66990 2320 66996 2332
rect 67048 2320 67054 2372
rect 69658 2320 69664 2372
rect 69716 2360 69722 2372
rect 82096 2360 82124 2400
rect 69716 2332 82124 2360
rect 69716 2320 69722 2332
rect 82262 2320 82268 2372
rect 82320 2360 82326 2372
rect 86926 2360 86954 2808
rect 96586 2564 96614 2808
rect 98012 2632 98040 2876
rect 100588 2774 100616 3012
rect 107626 2972 107654 3012
rect 109144 3012 117964 3040
rect 109144 2972 109172 3012
rect 117958 3000 117964 3012
rect 118016 3000 118022 3052
rect 107626 2944 109172 2972
rect 112438 2932 112444 2984
rect 112496 2972 112502 2984
rect 117682 2972 117688 2984
rect 112496 2944 117688 2972
rect 112496 2932 112502 2944
rect 117682 2932 117688 2944
rect 117740 2932 117746 2984
rect 116118 2904 116124 2916
rect 105280 2876 116124 2904
rect 100588 2746 100708 2774
rect 100680 2700 100708 2746
rect 98472 2672 100708 2700
rect 98472 2644 98500 2672
rect 98362 2632 98368 2644
rect 98012 2604 98368 2632
rect 98362 2592 98368 2604
rect 98420 2592 98426 2644
rect 98454 2592 98460 2644
rect 98512 2592 98518 2644
rect 100018 2592 100024 2644
rect 100076 2632 100082 2644
rect 105280 2632 105308 2876
rect 116118 2864 116124 2876
rect 116176 2864 116182 2916
rect 100076 2604 105308 2632
rect 105372 2808 293954 2836
rect 100076 2592 100082 2604
rect 105372 2564 105400 2808
rect 96586 2536 105400 2564
rect 98362 2456 98368 2508
rect 98420 2496 98426 2508
rect 100018 2496 100024 2508
rect 98420 2468 100024 2496
rect 98420 2456 98426 2468
rect 100018 2456 100024 2468
rect 100076 2456 100082 2508
rect 109586 2456 109592 2508
rect 109644 2496 109650 2508
rect 116578 2496 116584 2508
rect 109644 2468 116584 2496
rect 109644 2456 109650 2468
rect 116578 2456 116584 2468
rect 116636 2456 116642 2508
rect 293926 2496 293954 2808
rect 425808 2808 443684 2836
rect 425808 2508 425836 2808
rect 443656 2508 443684 2808
rect 294782 2496 294788 2508
rect 293926 2468 294788 2496
rect 294782 2456 294788 2468
rect 294840 2456 294846 2508
rect 425790 2456 425796 2508
rect 425848 2456 425854 2508
rect 443638 2456 443644 2508
rect 443696 2456 443702 2508
rect 106182 2388 106188 2440
rect 106240 2428 106246 2440
rect 116670 2428 116676 2440
rect 106240 2400 116676 2428
rect 106240 2388 106246 2400
rect 116670 2388 116676 2400
rect 116728 2388 116734 2440
rect 82320 2332 86954 2360
rect 82320 2320 82326 2332
rect 102962 2320 102968 2372
rect 103020 2360 103026 2372
rect 116762 2360 116768 2372
rect 103020 2332 116768 2360
rect 103020 2320 103026 2332
rect 116762 2320 116768 2332
rect 116820 2320 116826 2372
rect 49602 2252 49608 2304
rect 49660 2292 49666 2304
rect 49660 2264 52454 2292
rect 49660 2252 49666 2264
rect 52426 2156 52454 2264
rect 58802 2252 58808 2304
rect 58860 2292 58866 2304
rect 81986 2292 81992 2304
rect 58860 2264 81992 2292
rect 58860 2252 58866 2264
rect 81986 2252 81992 2264
rect 82044 2252 82050 2304
rect 99650 2252 99656 2304
rect 99708 2292 99714 2304
rect 116854 2292 116860 2304
rect 99708 2264 116860 2292
rect 99708 2252 99714 2264
rect 116854 2252 116860 2264
rect 116912 2252 116918 2304
rect 56226 2184 56232 2236
rect 56284 2224 56290 2236
rect 73062 2224 73068 2236
rect 56284 2196 73068 2224
rect 56284 2184 56290 2196
rect 73062 2184 73068 2196
rect 73120 2184 73126 2236
rect 80238 2184 80244 2236
rect 80296 2224 80302 2236
rect 81526 2224 81532 2236
rect 80296 2196 81532 2224
rect 80296 2184 80302 2196
rect 81526 2184 81532 2196
rect 81584 2184 81590 2236
rect 82078 2184 82084 2236
rect 82136 2224 82142 2236
rect 82446 2224 82452 2236
rect 82136 2196 82452 2224
rect 82136 2184 82142 2196
rect 82446 2184 82452 2196
rect 82504 2184 82510 2236
rect 96338 2184 96344 2236
rect 96396 2224 96402 2236
rect 117038 2224 117044 2236
rect 96396 2196 117044 2224
rect 96396 2184 96402 2196
rect 117038 2184 117044 2196
rect 117096 2184 117102 2236
rect 63310 2156 63316 2168
rect 52426 2128 63316 2156
rect 63310 2116 63316 2128
rect 63368 2116 63374 2168
rect 80330 2116 80336 2168
rect 80388 2156 80394 2168
rect 81802 2156 81808 2168
rect 80388 2128 81808 2156
rect 80388 2116 80394 2128
rect 81802 2116 81808 2128
rect 81860 2116 81866 2168
rect 93026 2116 93032 2168
rect 93084 2156 93090 2168
rect 117222 2156 117228 2168
rect 93084 2128 117228 2156
rect 93084 2116 93090 2128
rect 117222 2116 117228 2128
rect 117280 2116 117286 2168
rect 80422 2048 80428 2100
rect 80480 2088 80486 2100
rect 81618 2088 81624 2100
rect 80480 2060 81624 2088
rect 80480 2048 80486 2060
rect 81618 2048 81624 2060
rect 81676 2048 81682 2100
rect 89622 2048 89628 2100
rect 89680 2088 89686 2100
rect 117314 2088 117320 2100
rect 89680 2060 117320 2088
rect 89680 2048 89686 2060
rect 117314 2048 117320 2060
rect 117372 2048 117378 2100
rect 86402 1980 86408 2032
rect 86460 2020 86466 2032
rect 117130 2020 117136 2032
rect 86460 1992 117136 2020
rect 86460 1980 86466 1992
rect 117130 1980 117136 1992
rect 117188 1980 117194 2032
rect 82630 1912 82636 1964
rect 82688 1952 82694 1964
rect 116486 1952 116492 1964
rect 82688 1924 116492 1952
rect 82688 1912 82694 1924
rect 116486 1912 116492 1924
rect 116544 1912 116550 1964
rect 79318 1844 79324 1896
rect 79376 1884 79382 1896
rect 116394 1884 116400 1896
rect 79376 1856 116400 1884
rect 79376 1844 79382 1856
rect 116394 1844 116400 1856
rect 116452 1844 116458 1896
rect 72694 1776 72700 1828
rect 72752 1816 72758 1828
rect 109678 1816 109684 1828
rect 72752 1788 109684 1816
rect 72752 1776 72758 1788
rect 109678 1776 109684 1788
rect 109736 1776 109742 1828
rect 76006 1708 76012 1760
rect 76064 1748 76070 1760
rect 116210 1748 116216 1760
rect 76064 1720 116216 1748
rect 76064 1708 76070 1720
rect 116210 1708 116216 1720
rect 116268 1708 116274 1760
rect 32674 1640 32680 1692
rect 32732 1680 32738 1692
rect 116026 1680 116032 1692
rect 32732 1652 116032 1680
rect 32732 1640 32738 1652
rect 116026 1640 116032 1652
rect 116084 1640 116090 1692
rect 29270 1572 29276 1624
rect 29328 1612 29334 1624
rect 115934 1612 115940 1624
rect 29328 1584 115940 1612
rect 29328 1572 29334 1584
rect 115934 1572 115940 1584
rect 115992 1572 115998 1624
rect 25958 1504 25964 1556
rect 26016 1544 26022 1556
rect 116946 1544 116952 1556
rect 26016 1516 116952 1544
rect 26016 1504 26022 1516
rect 116946 1504 116952 1516
rect 117004 1504 117010 1556
rect 22646 1436 22652 1488
rect 22704 1476 22710 1488
rect 116302 1476 116308 1488
rect 22704 1448 116308 1476
rect 22704 1436 22710 1448
rect 116302 1436 116308 1448
rect 116360 1436 116366 1488
rect 117682 1436 117688 1488
rect 117740 1476 117746 1488
rect 143626 1476 143632 1488
rect 117740 1448 143632 1476
rect 117740 1436 117746 1448
rect 143626 1436 143632 1448
rect 143684 1436 143690 1488
rect 5994 1368 6000 1420
rect 6052 1408 6058 1420
rect 109770 1408 109776 1420
rect 6052 1380 109776 1408
rect 6052 1368 6058 1380
rect 109770 1368 109776 1380
rect 109828 1368 109834 1420
rect 117958 1368 117964 1420
rect 118016 1408 118022 1420
rect 193582 1408 193588 1420
rect 118016 1380 193588 1408
rect 118016 1368 118022 1380
rect 193582 1368 193588 1380
rect 193640 1368 193646 1420
rect 294782 1368 294788 1420
rect 294840 1408 294846 1420
rect 343634 1408 343640 1420
rect 294840 1380 343640 1408
rect 294840 1368 294846 1380
rect 343634 1368 343640 1380
rect 343692 1368 343698 1420
rect 491294 1368 491300 1420
rect 491352 1408 491358 1420
rect 493594 1408 493600 1420
rect 491352 1380 493600 1408
rect 491352 1368 491358 1380
rect 493594 1368 493600 1380
rect 493652 1368 493658 1420
<< via1 >>
rect 168564 160284 168616 160336
rect 173348 160284 173400 160336
rect 63408 160012 63460 160064
rect 146484 160012 146536 160064
rect 146944 160012 146996 160064
rect 154488 160012 154540 160064
rect 156788 160012 156840 160064
rect 191656 160012 191708 160064
rect 197176 160012 197228 160064
rect 207020 160012 207072 160064
rect 211436 160012 211488 160064
rect 280344 160012 280396 160064
rect 281264 160012 281316 160064
rect 332692 160012 332744 160064
rect 334256 160012 334308 160064
rect 374092 160012 374144 160064
rect 378876 160012 378928 160064
rect 391388 160012 391440 160064
rect 391480 160012 391532 160064
rect 394608 160012 394660 160064
rect 400772 160012 400824 160064
rect 424876 160012 424928 160064
rect 25596 159944 25648 159996
rect 110328 159944 110380 159996
rect 117228 159944 117280 159996
rect 191472 159944 191524 159996
rect 198004 159944 198056 159996
rect 269120 159944 269172 159996
rect 271236 159944 271288 159996
rect 272800 159944 272852 159996
rect 275376 159944 275428 159996
rect 328460 159944 328512 159996
rect 329196 159944 329248 159996
rect 369952 159944 370004 159996
rect 372160 159944 372212 159996
rect 396172 159944 396224 159996
rect 403256 159944 403308 159996
rect 415860 159944 415912 159996
rect 76932 159876 76984 159928
rect 162492 159876 162544 159928
rect 166908 159876 166960 159928
rect 186412 159876 186464 159928
rect 191288 159876 191340 159928
rect 264888 159876 264940 159928
rect 268660 159876 268712 159928
rect 324044 159876 324096 159928
rect 328368 159876 328420 159928
rect 369492 159876 369544 159928
rect 379704 159876 379756 159928
rect 405832 159876 405884 159928
rect 457076 159876 457128 159928
rect 464344 159876 464396 159928
rect 480628 159876 480680 159928
rect 485964 159876 486016 159928
rect 70124 159808 70176 159860
rect 156328 159808 156380 159860
rect 56692 159740 56744 159792
rect 137284 159740 137336 159792
rect 137376 159740 137428 159792
rect 139400 159740 139452 159792
rect 139952 159740 140004 159792
rect 147036 159740 147088 159792
rect 147128 159740 147180 159792
rect 148324 159740 148376 159792
rect 153476 159740 153528 159792
rect 156604 159740 156656 159792
rect 18880 159672 18932 159724
rect 109224 159672 109276 159724
rect 113088 159672 113140 159724
rect 126428 159672 126480 159724
rect 126520 159672 126572 159724
rect 156512 159672 156564 159724
rect 160100 159808 160152 159860
rect 156788 159740 156840 159792
rect 179420 159808 179472 159860
rect 184572 159808 184624 159860
rect 259552 159808 259604 159860
rect 261116 159808 261168 159860
rect 317052 159808 317104 159860
rect 320824 159808 320876 159860
rect 362960 159808 363012 159860
rect 376300 159808 376352 159860
rect 406200 159808 406252 159860
rect 409972 159808 410024 159860
rect 417240 159808 417292 159860
rect 446128 159808 446180 159860
rect 456800 159808 456852 159860
rect 458732 159808 458784 159860
rect 465080 159808 465132 159860
rect 472256 159808 472308 159860
rect 479432 159808 479484 159860
rect 171140 159740 171192 159792
rect 173256 159740 173308 159792
rect 177856 159740 177908 159792
rect 253940 159740 253992 159792
rect 261944 159740 261996 159792
rect 318892 159740 318944 159792
rect 322480 159740 322532 159792
rect 365168 159740 365220 159792
rect 365444 159740 365496 159792
rect 395528 159740 395580 159792
rect 396540 159740 396592 159792
rect 413192 159740 413244 159792
rect 413376 159740 413428 159792
rect 419632 159740 419684 159792
rect 420920 159740 420972 159792
rect 440424 159740 440476 159792
rect 448704 159740 448756 159792
rect 460940 159740 460992 159792
rect 469680 159740 469732 159792
rect 477408 159740 477460 159792
rect 478972 159740 479024 159792
rect 484676 159740 484728 159792
rect 49976 159604 50028 159656
rect 143264 159604 143316 159656
rect 143356 159604 143408 159656
rect 43260 159536 43312 159588
rect 136824 159536 136876 159588
rect 137284 159536 137336 159588
rect 144000 159536 144052 159588
rect 144092 159536 144144 159588
rect 146852 159536 146904 159588
rect 147220 159536 147272 159588
rect 163780 159672 163832 159724
rect 167736 159672 167788 159724
rect 246948 159672 247000 159724
rect 255228 159672 255280 159724
rect 313372 159672 313424 159724
rect 314108 159672 314160 159724
rect 357992 159672 358044 159724
rect 369584 159672 369636 159724
rect 401048 159672 401100 159724
rect 407488 159672 407540 159724
rect 429936 159672 429988 159724
rect 451188 159672 451240 159724
rect 462320 159672 462372 159724
rect 468024 159672 468076 159724
rect 476028 159672 476080 159724
rect 479800 159672 479852 159724
rect 485228 159672 485280 159724
rect 161020 159604 161072 159656
rect 240324 159604 240376 159656
rect 241796 159604 241848 159656
rect 302240 159604 302292 159656
rect 302332 159604 302384 159656
rect 349252 159604 349304 159656
rect 351920 159604 351972 159656
rect 385776 159604 385828 159656
rect 388076 159604 388128 159656
rect 389088 159604 389140 159656
rect 389824 159604 389876 159656
rect 413376 159604 413428 159656
rect 417516 159604 417568 159656
rect 437664 159604 437716 159656
rect 453764 159604 453816 159656
rect 465264 159604 465316 159656
rect 157616 159536 157668 159588
rect 239312 159536 239364 159588
rect 250996 159536 251048 159588
rect 310612 159536 310664 159588
rect 315764 159536 315816 159588
rect 358912 159536 358964 159588
rect 362868 159536 362920 159588
rect 394976 159536 395028 159588
rect 399024 159536 399076 159588
rect 408500 159536 408552 159588
rect 410800 159536 410852 159588
rect 432512 159536 432564 159588
rect 452016 159536 452068 159588
rect 463976 159536 464028 159588
rect 467196 159536 467248 159588
rect 473360 159536 473412 159588
rect 36544 159468 36596 159520
rect 126336 159468 126388 159520
rect 126428 159468 126480 159520
rect 127624 159468 127676 159520
rect 129924 159468 129976 159520
rect 146944 159468 146996 159520
rect 32312 159400 32364 159452
rect 126612 159400 126664 159452
rect 130752 159400 130804 159452
rect 137192 159400 137244 159452
rect 6276 159332 6328 159384
rect 122840 159332 122892 159384
rect 123116 159332 123168 159384
rect 144092 159400 144144 159452
rect 144184 159400 144236 159452
rect 225328 159468 225380 159520
rect 231676 159468 231728 159520
rect 295524 159468 295576 159520
rect 295616 159468 295668 159520
rect 342444 159468 342496 159520
rect 347688 159468 347740 159520
rect 354220 159468 354272 159520
rect 356152 159468 356204 159520
rect 390560 159468 390612 159520
rect 391388 159468 391440 159520
rect 398564 159468 398616 159520
rect 424324 159468 424376 159520
rect 442816 159468 442868 159520
rect 447876 159468 447928 159520
rect 460112 159468 460164 159520
rect 461308 159468 461360 159520
rect 467932 159468 467984 159520
rect 481456 159468 481508 159520
rect 486516 159468 486568 159520
rect 518808 159468 518860 159520
rect 522672 159468 522724 159520
rect 147588 159400 147640 159452
rect 149520 159400 149572 159452
rect 150900 159400 150952 159452
rect 233240 159400 233292 159452
rect 234988 159400 235040 159452
rect 298008 159400 298060 159452
rect 301504 159400 301556 159452
rect 349068 159400 349120 159452
rect 349804 159400 349856 159452
rect 354864 159400 354916 159452
rect 358636 159400 358688 159452
rect 392768 159400 392820 159452
rect 404084 159400 404136 159452
rect 427360 159400 427412 159452
rect 427636 159400 427688 159452
rect 445392 159400 445444 159452
rect 449532 159400 449584 159452
rect 461492 159400 461544 159452
rect 468852 159400 468904 159452
rect 474832 159400 474884 159452
rect 477316 159400 477368 159452
rect 483296 159400 483348 159452
rect 137468 159332 137520 159384
rect 223580 159332 223632 159384
rect 224960 159332 225012 159384
rect 290648 159332 290700 159384
rect 294788 159332 294840 159384
rect 342260 159332 342312 159384
rect 342720 159332 342772 159384
rect 343640 159332 343692 159384
rect 346032 159332 346084 159384
rect 382832 159332 382884 159384
rect 414204 159332 414256 159384
rect 435088 159332 435140 159384
rect 450360 159332 450412 159384
rect 462688 159332 462740 159384
rect 470508 159332 470560 159384
rect 476120 159332 476172 159384
rect 478144 159332 478196 159384
rect 483204 159332 483256 159384
rect 518716 159332 518768 159384
rect 523500 159332 523552 159384
rect 73528 159264 73580 159316
rect 80060 159264 80112 159316
rect 83648 159264 83700 159316
rect 167000 159264 167052 159316
rect 170220 159264 170272 159316
rect 198924 159264 198976 159316
rect 201408 159264 201460 159316
rect 213736 159264 213788 159316
rect 214012 159264 214064 159316
rect 281540 159264 281592 159316
rect 282092 159264 282144 159316
rect 334348 159264 334400 159316
rect 335084 159264 335136 159316
rect 374736 159264 374788 159316
rect 378048 159264 378100 159316
rect 388352 159264 388404 159316
rect 388996 159264 389048 159316
rect 395160 159264 395212 159316
rect 462136 159264 462188 159316
rect 467840 159264 467892 159316
rect 80244 159196 80296 159248
rect 91100 159196 91152 159248
rect 100484 159196 100536 159248
rect 184388 159196 184440 159248
rect 187056 159196 187108 159248
rect 214564 159196 214616 159248
rect 218244 159196 218296 159248
rect 284392 159196 284444 159248
rect 287980 159196 288032 159248
rect 338764 159196 338816 159248
rect 339316 159196 339368 159248
rect 377956 159196 378008 159248
rect 385592 159196 385644 159248
rect 398840 159196 398892 159248
rect 459652 159196 459704 159248
rect 466644 159196 466696 159248
rect 86960 159128 87012 159180
rect 93676 159060 93728 159112
rect 162860 159060 162912 159112
rect 163044 159128 163096 159180
rect 172152 159128 172204 159180
rect 193772 159128 193824 159180
rect 218060 159128 218112 159180
rect 220728 159128 220780 159180
rect 283196 159128 283248 159180
rect 284668 159128 284720 159180
rect 285772 159128 285824 159180
rect 169760 159060 169812 159112
rect 171784 159060 171836 159112
rect 176660 159060 176712 159112
rect 180340 159060 180392 159112
rect 204904 159060 204956 159112
rect 224132 159060 224184 159112
rect 288164 159128 288216 159180
rect 288900 159128 288952 159180
rect 338396 159128 338448 159180
rect 338488 159128 338540 159180
rect 339684 159128 339736 159180
rect 341892 159128 341944 159180
rect 378232 159128 378284 159180
rect 383108 159128 383160 159180
rect 302240 159060 302292 159112
rect 303528 159060 303580 159112
rect 309048 159060 309100 159112
rect 349804 159060 349856 159112
rect 107200 158992 107252 159044
rect 183468 158992 183520 159044
rect 183744 158992 183796 159044
rect 201408 158992 201460 159044
rect 203892 158992 203944 159044
rect 212724 158992 212776 159044
rect 230848 158992 230900 159044
rect 295156 158992 295208 159044
rect 298100 158992 298152 159044
rect 299572 158992 299624 159044
rect 96252 158924 96304 158976
rect 121920 158924 121972 158976
rect 124036 158924 124088 158976
rect 194140 158924 194192 158976
rect 194692 158924 194744 158976
rect 204168 158924 204220 158976
rect 207296 158924 207348 158976
rect 230756 158924 230808 158976
rect 237564 158924 237616 158976
rect 299480 158924 299532 158976
rect 102968 158856 103020 158908
rect 125508 158856 125560 158908
rect 126336 158856 126388 158908
rect 129740 158856 129792 158908
rect 109684 158788 109736 158840
rect 137100 158856 137152 158908
rect 137192 158856 137244 158908
rect 195428 158856 195480 158908
rect 210608 158856 210660 158908
rect 215392 158856 215444 158908
rect 217324 158856 217376 158908
rect 220360 158856 220412 158908
rect 238392 158856 238444 158908
rect 242440 158856 242492 158908
rect 244280 158856 244332 158908
rect 305368 158992 305420 159044
rect 307392 158992 307444 159044
rect 353208 159060 353260 159112
rect 357808 159060 357860 159112
rect 384948 159060 385000 159112
rect 351092 158992 351144 159044
rect 382556 158992 382608 159044
rect 133236 158788 133288 158840
rect 158720 158788 158772 158840
rect 163504 158788 163556 158840
rect 197268 158788 197320 158840
rect 208124 158788 208176 158840
rect 212448 158788 212500 158840
rect 214840 158788 214892 158840
rect 221464 158788 221516 158840
rect 221556 158788 221608 158840
rect 224592 158788 224644 158840
rect 248512 158788 248564 158840
rect 305644 158856 305696 158908
rect 307392 158856 307444 158908
rect 308220 158924 308272 158976
rect 347688 158924 347740 158976
rect 347780 158924 347832 158976
rect 378784 158924 378836 158976
rect 384764 158924 384816 158976
rect 392308 159128 392360 159180
rect 404268 159128 404320 159180
rect 462964 159128 463016 159180
rect 469220 159128 469272 159180
rect 395712 159060 395764 159112
rect 405648 159060 405700 159112
rect 457904 159060 457956 159112
rect 464528 159060 464580 159112
rect 471428 159060 471480 159112
rect 477684 159060 477736 159112
rect 395160 158992 395212 159044
rect 404176 158992 404228 159044
rect 460480 158992 460532 159044
rect 466460 158992 466512 159044
rect 473912 158992 473964 159044
rect 480260 158992 480312 159044
rect 308588 158856 308640 158908
rect 312452 158856 312504 158908
rect 313648 158856 313700 158908
rect 314936 158856 314988 158908
rect 357440 158856 357492 158908
rect 361212 158856 361264 158908
rect 386328 158856 386380 158908
rect 310704 158788 310756 158840
rect 313188 158788 313240 158840
rect 319168 158788 319220 158840
rect 321560 158788 321612 158840
rect 321652 158788 321704 158840
rect 363144 158788 363196 158840
rect 367928 158788 367980 158840
rect 385040 158788 385092 158840
rect 90364 158720 90416 158772
rect 92480 158720 92532 158772
rect 92848 158720 92900 158772
rect 114468 158720 114520 158772
rect 119804 158720 119856 158772
rect 146576 158720 146628 158772
rect 146668 158720 146720 158772
rect 171784 158720 171836 158772
rect 173624 158720 173676 158772
rect 197360 158720 197412 158772
rect 200580 158720 200632 158772
rect 224960 158720 225012 158772
rect 240876 158720 240928 158772
rect 243360 158720 243412 158772
rect 254400 158720 254452 158772
rect 255412 158720 255464 158772
rect 258540 158720 258592 158772
rect 260932 158720 260984 158772
rect 264428 158720 264480 158772
rect 266360 158720 266412 158772
rect 267832 158720 267884 158772
rect 320272 158720 320324 158772
rect 327540 158720 327592 158772
rect 367192 158720 367244 158772
rect 374644 158720 374696 158772
rect 388444 158720 388496 158772
rect 411352 158924 411404 158976
rect 416688 158924 416740 158976
rect 419540 158924 419592 158976
rect 420092 158924 420144 158976
rect 423588 158924 423640 158976
rect 456248 158924 456300 158976
rect 463148 158924 463200 158976
rect 466368 158924 466420 158976
rect 472348 158924 472400 158976
rect 475568 158924 475620 158976
rect 482008 158924 482060 158976
rect 412548 158856 412600 158908
rect 412824 158856 412876 158908
rect 454592 158856 454644 158908
rect 461676 158856 461728 158908
rect 465540 158856 465592 158908
rect 472164 158856 472216 158908
rect 474740 158856 474792 158908
rect 481364 158856 481416 158908
rect 508320 158856 508372 158908
rect 510068 158856 510120 158908
rect 389088 158788 389140 158840
rect 390376 158788 390428 158840
rect 409144 158788 409196 158840
rect 410708 158788 410760 158840
rect 455420 158788 455472 158840
rect 463608 158788 463660 158840
rect 464620 158788 464672 158840
rect 471428 158788 471480 158840
rect 476396 158788 476448 158840
rect 481640 158788 481692 158840
rect 506388 158788 506440 158840
rect 507584 158788 507636 158840
rect 389180 158720 389232 158772
rect 405740 158720 405792 158772
rect 409236 158720 409288 158772
rect 452844 158720 452896 158772
rect 459560 158720 459612 158772
rect 463792 158720 463844 158772
rect 471796 158720 471848 158772
rect 473084 158720 473136 158772
rect 478972 158720 479024 158772
rect 482284 158720 482336 158772
rect 487252 158720 487304 158772
rect 505284 158720 505336 158772
rect 506756 158720 506808 158772
rect 507032 158720 507084 158772
rect 508412 158720 508464 158772
rect 509424 158720 509476 158772
rect 511724 158720 511776 158772
rect 514944 158720 514996 158772
rect 518532 158720 518584 158772
rect 81072 158652 81124 158704
rect 180892 158652 180944 158704
rect 181996 158652 182048 158704
rect 256792 158652 256844 158704
rect 67640 158584 67692 158636
rect 166080 158584 166132 158636
rect 166540 158584 166592 158636
rect 172980 158584 173032 158636
rect 173348 158584 173400 158636
rect 247132 158584 247184 158636
rect 74356 158516 74408 158568
rect 172888 158516 172940 158568
rect 178684 158516 178736 158568
rect 255596 158516 255648 158568
rect 71044 158448 71096 158500
rect 165988 158448 166040 158500
rect 166448 158448 166500 158500
rect 170404 158448 170456 158500
rect 173164 158448 173216 158500
rect 175188 158448 175240 158500
rect 175280 158448 175332 158500
rect 252744 158448 252796 158500
rect 64236 158380 64288 158432
rect 167552 158380 167604 158432
rect 171968 158380 172020 158432
rect 250076 158380 250128 158432
rect 60924 158312 60976 158364
rect 164332 158312 164384 158364
rect 165252 158312 165304 158364
rect 245016 158312 245068 158364
rect 54208 158244 54260 158296
rect 160284 158244 160336 158296
rect 161848 158244 161900 158296
rect 242072 158244 242124 158296
rect 50804 158176 50856 158228
rect 157708 158176 157760 158228
rect 158444 158176 158496 158228
rect 238944 158176 238996 158228
rect 256884 158176 256936 158228
rect 315028 158176 315080 158228
rect 47492 158108 47544 158160
rect 155040 158108 155092 158160
rect 155132 158108 155184 158160
rect 237380 158108 237432 158160
rect 246764 158108 246816 158160
rect 306932 158108 306984 158160
rect 37372 158040 37424 158092
rect 146392 158040 146444 158092
rect 148416 158040 148468 158092
rect 231952 158040 232004 158092
rect 243452 158040 243504 158092
rect 304724 158040 304776 158092
rect 388 157972 440 158024
rect 118884 157972 118936 158024
rect 131580 157972 131632 158024
rect 219348 157972 219400 158024
rect 236736 157972 236788 158024
rect 299664 157972 299716 158024
rect 77760 157904 77812 157956
rect 87788 157836 87840 157888
rect 164884 157836 164936 157888
rect 84476 157768 84528 157820
rect 170036 157768 170088 157820
rect 170220 157904 170272 157956
rect 182272 157904 182324 157956
rect 170496 157836 170548 157888
rect 185124 157836 185176 157888
rect 178040 157768 178092 157820
rect 179420 157768 179472 157820
rect 185308 157904 185360 157956
rect 185400 157904 185452 157956
rect 260472 157904 260524 157956
rect 188804 157836 188856 157888
rect 263048 157836 263100 157888
rect 91192 157700 91244 157752
rect 185308 157700 185360 157752
rect 94596 157632 94648 157684
rect 190644 157768 190696 157820
rect 195520 157768 195572 157820
rect 267740 157768 267792 157820
rect 185676 157700 185728 157752
rect 188528 157700 188580 157752
rect 190460 157700 190512 157752
rect 263692 157700 263744 157752
rect 185584 157632 185636 157684
rect 236092 157632 236144 157684
rect 97908 157564 97960 157616
rect 193220 157564 193272 157616
rect 197360 157564 197412 157616
rect 251456 157564 251508 157616
rect 111340 157496 111392 157548
rect 203984 157496 204036 157548
rect 204904 157496 204956 157548
rect 255872 157496 255924 157548
rect 114744 157428 114796 157480
rect 206560 157428 206612 157480
rect 141700 157360 141752 157412
rect 227076 157360 227128 157412
rect 49148 157292 49200 157344
rect 156420 157292 156472 157344
rect 158720 157292 158772 157344
rect 219992 157292 220044 157344
rect 45744 157224 45796 157276
rect 153844 157224 153896 157276
rect 163780 157224 163832 157276
rect 166448 157224 166500 157276
rect 192116 157224 192168 157276
rect 265164 157224 265216 157276
rect 283840 157224 283892 157276
rect 335544 157224 335596 157276
rect 42432 157156 42484 157208
rect 151268 157156 151320 157208
rect 156512 157156 156564 157208
rect 159088 157156 159140 157208
rect 160100 157156 160152 157208
rect 166172 157156 166224 157208
rect 166264 157156 166316 157208
rect 171140 157156 171192 157208
rect 177028 157156 177080 157208
rect 254032 157156 254084 157208
rect 300676 157156 300728 157208
rect 348056 157156 348108 157208
rect 39028 157088 39080 157140
rect 148784 157088 148836 157140
rect 150072 157088 150124 157140
rect 233516 157088 233568 157140
rect 280436 157088 280488 157140
rect 333060 157088 333112 157140
rect 35716 157020 35768 157072
rect 146208 157020 146260 157072
rect 151728 157020 151780 157072
rect 234804 157020 234856 157072
rect 273720 157020 273772 157072
rect 327908 157020 327960 157072
rect 24768 156952 24820 157004
rect 137376 156952 137428 157004
rect 138296 156952 138348 157004
rect 224132 156952 224184 157004
rect 224960 156952 225012 157004
rect 272064 156952 272116 157004
rect 277124 156952 277176 157004
rect 330484 156952 330536 157004
rect 21364 156884 21416 156936
rect 135260 156884 135312 156936
rect 135812 156884 135864 156936
rect 222568 156884 222620 156936
rect 226616 156884 226668 156936
rect 291936 156884 291988 156936
rect 293868 156884 293920 156936
rect 342720 156884 342772 156936
rect 18052 156816 18104 156868
rect 132500 156816 132552 156868
rect 134892 156816 134944 156868
rect 221372 156816 221424 156868
rect 223212 156816 223264 156868
rect 289360 156816 289412 156868
rect 290556 156816 290608 156868
rect 340052 156816 340104 156868
rect 14648 156748 14700 156800
rect 130108 156748 130160 156800
rect 139124 156748 139176 156800
rect 225144 156748 225196 156800
rect 230020 156748 230072 156800
rect 294052 156748 294104 156800
rect 297272 156748 297324 156800
rect 345112 156748 345164 156800
rect 11244 156680 11296 156732
rect 127532 156680 127584 156732
rect 128176 156680 128228 156732
rect 212540 156680 212592 156732
rect 2044 156612 2096 156664
rect 120448 156612 120500 156664
rect 124864 156612 124916 156664
rect 211804 156612 211856 156664
rect 52460 156544 52512 156596
rect 158996 156544 159048 156596
rect 159088 156544 159140 156596
rect 215484 156680 215536 156732
rect 219900 156680 219952 156732
rect 286232 156680 286284 156732
rect 287152 156680 287204 156732
rect 338120 156680 338172 156732
rect 216496 156612 216548 156664
rect 283104 156612 283156 156664
rect 498292 156612 498344 156664
rect 499304 156612 499356 156664
rect 213828 156544 213880 156596
rect 281632 156544 281684 156596
rect 59268 156476 59320 156528
rect 164148 156476 164200 156528
rect 166172 156476 166224 156528
rect 69296 156408 69348 156460
rect 166264 156408 166316 156460
rect 166448 156476 166500 156528
rect 225052 156476 225104 156528
rect 228364 156408 228416 156460
rect 82820 156340 82872 156392
rect 182088 156340 182140 156392
rect 198832 156340 198884 156392
rect 200856 156340 200908 156392
rect 209780 156340 209832 156392
rect 279056 156340 279108 156392
rect 99564 156272 99616 156324
rect 194968 156272 195020 156324
rect 101312 156204 101364 156256
rect 196256 156204 196308 156256
rect 108028 156136 108080 156188
rect 200396 156136 200448 156188
rect 118148 156068 118200 156120
rect 209136 156272 209188 156324
rect 212540 156272 212592 156324
rect 216772 156272 216824 156324
rect 218060 156272 218112 156324
rect 266912 156272 266964 156324
rect 200672 156204 200724 156256
rect 201316 156204 201368 156256
rect 203064 156204 203116 156256
rect 121460 156000 121512 156052
rect 211620 156136 211672 156188
rect 211804 156136 211856 156188
rect 213920 156136 213972 156188
rect 230756 156204 230808 156256
rect 277124 156204 277176 156256
rect 273904 156136 273956 156188
rect 202328 156068 202380 156120
rect 273260 156068 273312 156120
rect 200856 156000 200908 156052
rect 270500 156000 270552 156052
rect 145012 155932 145064 155984
rect 229652 155932 229704 155984
rect 66812 155864 66864 155916
rect 82820 155864 82872 155916
rect 89536 155864 89588 155916
rect 186320 155864 186372 155916
rect 186412 155864 186464 155916
rect 192852 155864 192904 155916
rect 192944 155864 192996 155916
rect 266268 155864 266320 155916
rect 296444 155864 296496 155916
rect 345204 155864 345256 155916
rect 60096 155796 60148 155848
rect 79324 155796 79376 155848
rect 88708 155796 88760 155848
rect 186872 155796 186924 155848
rect 189632 155796 189684 155848
rect 263784 155796 263836 155848
rect 293040 155796 293092 155848
rect 342352 155796 342404 155848
rect 12164 155728 12216 155780
rect 109132 155728 109184 155780
rect 112260 155728 112312 155780
rect 204628 155728 204680 155780
rect 206468 155728 206520 155780
rect 276112 155728 276164 155780
rect 289728 155728 289780 155780
rect 339592 155728 339644 155780
rect 46572 155660 46624 155712
rect 75460 155660 75512 155712
rect 81900 155660 81952 155712
rect 180984 155660 181036 155712
rect 186228 155660 186280 155712
rect 260840 155660 260892 155712
rect 270316 155660 270368 155712
rect 325332 155660 325384 155712
rect 344376 155660 344428 155712
rect 381820 155660 381872 155712
rect 53380 155592 53432 155644
rect 67088 155592 67140 155644
rect 71872 155592 71924 155644
rect 172704 155592 172756 155644
rect 176292 155592 176344 155644
rect 253388 155592 253440 155644
rect 267004 155592 267056 155644
rect 321744 155592 321796 155644
rect 340972 155592 341024 155644
rect 378140 155592 378192 155644
rect 39856 155524 39908 155576
rect 68836 155524 68888 155576
rect 75184 155524 75236 155576
rect 176384 155524 176436 155576
rect 179512 155524 179564 155576
rect 255780 155524 255832 155576
rect 263600 155524 263652 155576
rect 320180 155524 320232 155576
rect 337660 155524 337712 155576
rect 375564 155524 375616 155576
rect 65156 155456 65208 155508
rect 168656 155456 168708 155508
rect 169392 155456 169444 155508
rect 248236 155456 248288 155508
rect 260288 155456 260340 155508
rect 317604 155456 317656 155508
rect 333428 155456 333480 155508
rect 373448 155456 373500 155508
rect 8760 155388 8812 155440
rect 125692 155388 125744 155440
rect 145840 155388 145892 155440
rect 229192 155388 229244 155440
rect 253572 155388 253624 155440
rect 312452 155388 312504 155440
rect 330116 155388 330168 155440
rect 370872 155388 370924 155440
rect 7932 155320 7984 155372
rect 124680 155320 124732 155372
rect 142528 155320 142580 155372
rect 227812 155320 227864 155372
rect 250168 155320 250220 155372
rect 309876 155320 309928 155372
rect 319996 155320 320048 155372
rect 363236 155320 363288 155372
rect 4528 155252 4580 155304
rect 122012 155252 122064 155304
rect 125784 155252 125836 155304
rect 214840 155252 214892 155304
rect 240048 155252 240100 155304
rect 302332 155252 302384 155304
rect 306564 155252 306616 155304
rect 352472 155252 352524 155304
rect 373816 155252 373868 155304
rect 404084 155252 404136 155304
rect 5356 155184 5408 155236
rect 123024 155184 123076 155236
rect 129004 155184 129056 155236
rect 217416 155184 217468 155236
rect 233332 155184 233384 155236
rect 297088 155184 297140 155236
rect 299756 155184 299808 155236
rect 347872 155184 347924 155236
rect 370412 155184 370464 155236
rect 401692 155184 401744 155236
rect 92020 155116 92072 155168
rect 189172 155116 189224 155168
rect 192852 155116 192904 155168
rect 194324 155116 194376 155168
rect 196348 155116 196400 155168
rect 268844 155116 268896 155168
rect 303160 155116 303212 155168
rect 350356 155116 350408 155168
rect 95424 155048 95476 155100
rect 98736 154980 98788 155032
rect 186320 154980 186372 155032
rect 186780 155048 186832 155100
rect 191748 154980 191800 155032
rect 199660 155048 199712 155100
rect 271420 155048 271472 155100
rect 200120 154980 200172 155032
rect 207020 154980 207072 155032
rect 269488 154980 269540 155032
rect 15476 154912 15528 154964
rect 109040 154912 109092 154964
rect 122288 154912 122340 154964
rect 211252 154912 211304 154964
rect 214564 154912 214616 154964
rect 261392 154912 261444 154964
rect 106372 154844 106424 154896
rect 186412 154844 186464 154896
rect 186688 154844 186740 154896
rect 245844 154844 245896 154896
rect 110512 154776 110564 154828
rect 139308 154776 139360 154828
rect 149244 154776 149296 154828
rect 232872 154776 232924 154828
rect 109224 154708 109276 154760
rect 133052 154708 133104 154760
rect 151912 154708 151964 154760
rect 153108 154708 153160 154760
rect 155960 154708 156012 154760
rect 238024 154708 238076 154760
rect 159364 154640 159416 154692
rect 240600 154640 240652 154692
rect 118608 154572 118660 154624
rect 119988 154572 120040 154624
rect 137100 154572 137152 154624
rect 138020 154572 138072 154624
rect 48320 154504 48372 154556
rect 152648 154572 152700 154624
rect 162676 154572 162728 154624
rect 243084 154572 243136 154624
rect 152464 154504 152516 154556
rect 202696 154504 202748 154556
rect 218336 154504 218388 154556
rect 44180 154436 44232 154488
rect 142896 154436 142948 154488
rect 142988 154436 143040 154488
rect 188252 154436 188304 154488
rect 114468 154368 114520 154420
rect 118608 154368 118660 154420
rect 118700 154368 118752 154420
rect 119896 154368 119948 154420
rect 119988 154368 120040 154420
rect 189816 154436 189868 154488
rect 191012 154436 191064 154488
rect 188436 154368 188488 154420
rect 197544 154368 197596 154420
rect 198464 154436 198516 154488
rect 210424 154436 210476 154488
rect 215300 154436 215352 154488
rect 283656 154504 283708 154556
rect 285588 154504 285640 154556
rect 285680 154504 285732 154556
rect 337476 154504 337528 154556
rect 353668 154504 353720 154556
rect 388904 154504 388956 154556
rect 283288 154436 283340 154488
rect 334900 154436 334952 154488
rect 349528 154436 349580 154488
rect 386236 154436 386288 154488
rect 390652 154436 390704 154488
rect 417148 154436 417200 154488
rect 202052 154368 202104 154420
rect 205088 154368 205140 154420
rect 275836 154368 275888 154420
rect 276204 154368 276256 154420
rect 329932 154368 329984 154420
rect 346400 154368 346452 154420
rect 383752 154368 383804 154420
rect 397368 154368 397420 154420
rect 422300 154368 422352 154420
rect 34520 154300 34572 154352
rect 142620 154300 142672 154352
rect 142712 154300 142764 154352
rect 205272 154300 205324 154352
rect 208400 154300 208452 154352
rect 278412 154300 278464 154352
rect 278872 154300 278924 154352
rect 332416 154300 332468 154352
rect 342812 154300 342864 154352
rect 381176 154300 381228 154352
rect 393320 154300 393372 154352
rect 419724 154300 419776 154352
rect 434720 154300 434772 154352
rect 444288 154300 444340 154352
rect 37924 154232 37976 154284
rect 27252 154164 27304 154216
rect 136916 154164 136968 154216
rect 143080 154232 143132 154284
rect 152464 154232 152516 154284
rect 152648 154232 152700 154284
rect 155776 154232 155828 154284
rect 161480 154232 161532 154284
rect 166080 154232 166132 154284
rect 176660 154232 176712 154284
rect 179696 154232 179748 154284
rect 182180 154232 182232 154284
rect 258540 154232 258592 154284
rect 262220 154232 262272 154284
rect 319536 154232 319588 154284
rect 339500 154232 339552 154284
rect 378600 154232 378652 154284
rect 386512 154232 386564 154284
rect 414572 154232 414624 154284
rect 23480 154096 23532 154148
rect 137008 154096 137060 154148
rect 13820 154028 13872 154080
rect 129280 154028 129332 154080
rect 9680 153960 9732 154012
rect 126888 153960 126940 154012
rect 127624 153960 127676 154012
rect 129372 153960 129424 154012
rect 7104 153892 7156 153944
rect 124312 153892 124364 153944
rect 125508 153892 125560 153944
rect 129648 153960 129700 154012
rect 142436 154096 142488 154148
rect 142896 154164 142948 154216
rect 137284 154028 137336 154080
rect 139768 154028 139820 154080
rect 139860 154028 139912 154080
rect 142528 154028 142580 154080
rect 148140 154096 148192 154148
rect 148324 154096 148376 154148
rect 152280 154164 152332 154216
rect 163504 154164 163556 154216
rect 172520 154164 172572 154216
rect 250812 154164 250864 154216
rect 255320 154164 255372 154216
rect 314384 154164 314436 154216
rect 336832 154164 336884 154216
rect 376024 154164 376076 154216
rect 383660 154164 383712 154216
rect 411996 154164 412048 154216
rect 142988 154028 143040 154080
rect 143540 154028 143592 154080
rect 150624 154028 150676 154080
rect 153200 154096 153252 154148
rect 153292 154096 153344 154148
rect 158444 154096 158496 154148
rect 160192 154096 160244 154148
rect 152188 154028 152240 154080
rect 152372 154028 152424 154080
rect 161572 154028 161624 154080
rect 165620 154096 165672 154148
rect 245660 154096 245712 154148
rect 245936 154096 245988 154148
rect 306656 154096 306708 154148
rect 326712 154096 326764 154148
rect 368296 154096 368348 154148
rect 376852 154096 376904 154148
rect 406844 154096 406896 154148
rect 241244 154028 241296 154080
rect 248604 154028 248656 154080
rect 309232 154028 309284 154080
rect 323308 154028 323360 154080
rect 365812 154028 365864 154080
rect 380164 154028 380216 154080
rect 409420 154028 409472 154080
rect 132408 153892 132460 153944
rect 219900 153960 219952 154012
rect 222384 153960 222436 154012
rect 288716 153960 288768 154012
rect 313280 153960 313332 154012
rect 357900 153960 357952 154012
rect 367100 153960 367152 154012
rect 399116 153960 399168 154012
rect 138020 153892 138072 153944
rect 143080 153892 143132 153944
rect 143264 153892 143316 153944
rect 145564 153892 145616 153944
rect 480 153824 532 153876
rect 119804 153824 119856 153876
rect 119896 153824 119948 153876
rect 142804 153824 142856 153876
rect 143356 153824 143408 153876
rect 223212 153892 223264 153944
rect 225236 153892 225288 153944
rect 291292 153892 291344 153944
rect 316040 153892 316092 153944
rect 360660 153892 360712 153944
rect 363052 153892 363104 153944
rect 396540 153892 396592 153944
rect 401600 153892 401652 153944
rect 425520 153892 425572 153944
rect 147404 153824 147456 153876
rect 152372 153824 152424 153876
rect 51080 153756 51132 153808
rect 158352 153824 158404 153876
rect 158444 153824 158496 153876
rect 235448 153824 235500 153876
rect 241888 153824 241940 153876
rect 304080 153824 304132 153876
rect 309140 153824 309192 153876
rect 355508 153824 355560 153876
rect 356244 153824 356296 153876
rect 391480 153824 391532 153876
rect 397460 153824 397512 153876
rect 422852 153824 422904 153876
rect 152648 153756 152700 153808
rect 212908 153756 212960 153808
rect 231860 153756 231912 153808
rect 296444 153756 296496 153808
rect 360384 153756 360436 153808
rect 394056 153756 394108 153808
rect 61108 153688 61160 153740
rect 57980 153620 58032 153672
rect 152280 153620 152332 153672
rect 161480 153688 161532 153740
rect 161572 153688 161624 153740
rect 198464 153688 198516 153740
rect 198556 153688 198608 153740
rect 209780 153688 209832 153740
rect 229100 153688 229152 153740
rect 293868 153688 293920 153740
rect 154488 153620 154540 153672
rect 218060 153620 218112 153672
rect 235080 153620 235132 153672
rect 299020 153620 299072 153672
rect 78680 153552 78732 153604
rect 179604 153552 179656 153604
rect 179696 153552 179748 153604
rect 230940 153552 230992 153604
rect 238852 153552 238904 153604
rect 301596 153552 301648 153604
rect 102140 153484 102192 153536
rect 196900 153484 196952 153536
rect 197268 153484 197320 153536
rect 198648 153484 198700 153536
rect 198924 153484 198976 153536
rect 248880 153484 248932 153536
rect 252652 153484 252704 153536
rect 311808 153484 311860 153536
rect 104900 153416 104952 153468
rect 199476 153416 199528 153468
rect 108304 153348 108356 153400
rect 191012 153348 191064 153400
rect 191656 153348 191708 153400
rect 200212 153348 200264 153400
rect 115940 153280 115992 153332
rect 207848 153416 207900 153468
rect 207940 153416 207992 153468
rect 259184 153416 259236 153468
rect 265440 153416 265492 153468
rect 322204 153416 322256 153468
rect 41604 153212 41656 153264
rect 138388 153212 138440 153264
rect 142804 153212 142856 153264
rect 198556 153212 198608 153264
rect 198648 153212 198700 153264
rect 243728 153348 243780 153400
rect 259460 153348 259512 153400
rect 316960 153348 317012 153400
rect 200580 153280 200632 153332
rect 238668 153280 238720 153332
rect 269212 153280 269264 153332
rect 324688 153280 324740 153332
rect 201408 153212 201460 153264
rect 207940 153212 207992 153264
rect 272892 153212 272944 153264
rect 327264 153212 327316 153264
rect 113180 153144 113232 153196
rect 205916 153144 205968 153196
rect 215392 153144 215444 153196
rect 279700 153144 279752 153196
rect 285496 153144 285548 153196
rect 336832 153144 336884 153196
rect 339684 153144 339736 153196
rect 377312 153144 377364 153196
rect 378232 153144 378284 153196
rect 379888 153144 379940 153196
rect 385040 153144 385092 153196
rect 399760 153144 399812 153196
rect 402428 153144 402480 153196
rect 423496 153144 423548 153196
rect 423588 153144 423640 153196
rect 80060 153076 80112 153128
rect 175096 153076 175148 153128
rect 180800 153076 180852 153128
rect 257252 153076 257304 153128
rect 264980 153076 265032 153128
rect 321468 153076 321520 153128
rect 324320 153076 324372 153128
rect 367008 153076 367060 153128
rect 367192 153076 367244 153128
rect 368940 153076 368992 153128
rect 380992 153076 381044 153128
rect 410064 153076 410116 153128
rect 410708 153076 410760 153128
rect 421012 153076 421064 153128
rect 422576 153076 422628 153128
rect 429476 153076 429528 153128
rect 430212 153144 430264 153196
rect 447324 153144 447376 153196
rect 456800 153144 456852 153196
rect 459468 153144 459520 153196
rect 461676 153144 461728 153196
rect 465908 153144 465960 153196
rect 466460 153144 466512 153196
rect 470416 153144 470468 153196
rect 471796 153144 471848 153196
rect 472992 153144 473044 153196
rect 473360 153144 473412 153196
rect 475568 153144 475620 153196
rect 476120 153144 476172 153196
rect 478144 153144 478196 153196
rect 484032 153144 484084 153196
rect 488448 153144 488500 153196
rect 489920 153144 489972 153196
rect 492864 153144 492916 153196
rect 494060 153144 494112 153196
rect 496084 153144 496136 153196
rect 496636 153144 496688 153196
rect 498016 153144 498068 153196
rect 510988 153144 511040 153196
rect 513472 153144 513524 153196
rect 514208 153144 514260 153196
rect 517428 153144 517480 153196
rect 431868 153076 431920 153128
rect 431960 153076 432012 153128
rect 441988 153076 442040 153128
rect 103520 153008 103572 153060
rect 198188 153008 198240 153060
rect 204168 153008 204220 153060
rect 267556 153008 267608 153060
rect 272156 153008 272208 153060
rect 326620 153008 326672 153060
rect 330944 153008 330996 153060
rect 371516 153008 371568 153060
rect 375472 153008 375524 153060
rect 398104 153008 398156 153060
rect 405832 153008 405884 153060
rect 408776 153008 408828 153060
rect 413376 153008 413428 153060
rect 416504 153008 416556 153060
rect 419264 153008 419316 153060
rect 434628 153008 434680 153060
rect 436100 153008 436152 153060
rect 437756 153008 437808 153060
rect 437848 153008 437900 153060
rect 442172 153076 442224 153128
rect 92480 152940 92532 152992
rect 187884 152940 187936 152992
rect 195428 152940 195480 152992
rect 218704 152940 218756 152992
rect 220360 152940 220412 152992
rect 284852 152940 284904 152992
rect 288164 152940 288216 152992
rect 290004 152940 290056 152992
rect 291384 152940 291436 152992
rect 341340 152940 341392 152992
rect 342260 152940 342312 152992
rect 343916 152940 343968 152992
rect 345296 152940 345348 152992
rect 382464 152940 382516 152992
rect 382556 152940 382608 152992
rect 386972 152940 387024 152992
rect 390376 152940 390428 152992
rect 415216 152940 415268 152992
rect 415400 152940 415452 152992
rect 436376 152940 436428 152992
rect 437480 152940 437532 152992
rect 441896 152940 441948 152992
rect 96620 152872 96672 152924
rect 193036 152872 193088 152924
rect 212448 152872 212500 152924
rect 277768 152872 277820 152924
rect 278780 152872 278832 152924
rect 331772 152872 331824 152924
rect 335360 152872 335412 152924
rect 375380 152872 375432 152924
rect 382188 152872 382240 152924
rect 410708 152872 410760 152924
rect 411260 152872 411312 152924
rect 433156 152872 433208 152924
rect 433524 152872 433576 152924
rect 449900 153076 449952 153128
rect 463608 153076 463660 153128
rect 466552 153076 466604 153128
rect 466644 153076 466696 153128
rect 469772 153076 469824 153128
rect 471428 153076 471480 153128
rect 473636 153076 473688 153128
rect 474832 153076 474884 153128
rect 476856 153076 476908 153128
rect 484952 153076 485004 153128
rect 489644 153076 489696 153128
rect 491668 153076 491720 153128
rect 494796 153076 494848 153128
rect 494980 153076 495032 153128
rect 496728 153076 496780 153128
rect 496820 153076 496872 153128
rect 498660 153076 498712 153128
rect 512920 153076 512972 153128
rect 515220 153076 515272 153128
rect 33140 152804 33192 152856
rect 138020 152804 138072 152856
rect 138112 152804 138164 152856
rect 141700 152804 141752 152856
rect 146484 152804 146536 152856
rect 167368 152804 167420 152856
rect 173900 152804 173952 152856
rect 252100 152804 252152 152856
rect 255412 152804 255464 152856
rect 313096 152804 313148 152856
rect 313188 152804 313240 152856
rect 356152 152804 356204 152856
rect 357440 152804 357492 152856
rect 359372 152804 359424 152856
rect 361580 152804 361632 152856
rect 395252 152804 395304 152856
rect 395528 152804 395580 152856
rect 397828 152804 397880 152856
rect 399208 152804 399260 152856
rect 424232 152804 424284 152856
rect 26424 152736 26476 152788
rect 139124 152736 139176 152788
rect 140780 152736 140832 152788
rect 144276 152736 144328 152788
rect 144368 152736 144420 152788
rect 162216 152736 162268 152788
rect 164424 152736 164476 152788
rect 244372 152736 244424 152788
rect 257712 152736 257764 152788
rect 315672 152736 315724 152788
rect 317052 152736 317104 152788
rect 318248 152736 318300 152788
rect 320272 152736 320324 152788
rect 323124 152736 323176 152788
rect 324228 152736 324280 152788
rect 366364 152736 366416 152788
rect 372620 152736 372672 152788
rect 403624 152736 403676 152788
rect 406660 152736 406712 152788
rect 422944 152736 422996 152788
rect 423496 152736 423548 152788
rect 426164 152804 426216 152856
rect 426440 152804 426492 152856
rect 440148 152804 440200 152856
rect 440240 152804 440292 152856
rect 455052 153008 455104 153060
rect 463148 153008 463200 153060
rect 467196 153008 467248 153060
rect 472164 153008 472216 153060
rect 474280 153008 474332 153060
rect 484400 153008 484452 153060
rect 489000 153008 489052 153060
rect 492680 153008 492732 153060
rect 495440 153008 495492 153060
rect 495532 153008 495584 153060
rect 497372 153008 497424 153060
rect 442540 152940 442592 152992
rect 453120 152940 453172 152992
rect 464528 152940 464580 152992
rect 468392 152940 468444 152992
rect 472348 152940 472400 152992
rect 474924 152940 474976 152992
rect 483112 152940 483164 152992
rect 487804 152940 487856 152992
rect 491300 152940 491352 152992
rect 494152 152940 494204 152992
rect 512276 152940 512328 152992
rect 514760 152940 514812 152992
rect 443000 152872 443052 152924
rect 451188 152872 451240 152924
rect 465080 152872 465132 152924
rect 469128 152872 469180 152924
rect 490012 152872 490064 152924
rect 493508 152872 493560 152924
rect 442448 152804 442500 152856
rect 444380 152804 444432 152856
rect 446312 152804 446364 152856
rect 460020 152804 460072 152856
rect 510344 152804 510396 152856
rect 512000 152804 512052 152856
rect 425244 152736 425296 152788
rect 434260 152736 434312 152788
rect 434352 152736 434404 152788
rect 450544 152736 450596 152788
rect 28172 152668 28224 152720
rect 141056 152668 141108 152720
rect 142804 152668 142856 152720
rect 149428 152668 149480 152720
rect 149520 152668 149572 152720
rect 231584 152668 231636 152720
rect 240324 152668 240376 152720
rect 241888 152668 241940 152720
rect 247040 152668 247092 152720
rect 307944 152668 307996 152720
rect 318340 152668 318392 152720
rect 361948 152668 362000 152720
rect 368480 152668 368532 152720
rect 400404 152668 400456 152720
rect 404360 152668 404412 152720
rect 428004 152668 428056 152720
rect 430580 152668 430632 152720
rect 447968 152668 448020 152720
rect 22192 152600 22244 152652
rect 135904 152600 135956 152652
rect 19340 152532 19392 152584
rect 133972 152532 134024 152584
rect 136824 152532 136876 152584
rect 151912 152600 151964 152652
rect 153568 152600 153620 152652
rect 236736 152600 236788 152652
rect 244464 152600 244516 152652
rect 306012 152600 306064 152652
rect 311532 152600 311584 152652
rect 356796 152600 356848 152652
rect 358820 152600 358872 152652
rect 393412 152600 393464 152652
rect 394884 152600 394936 152652
rect 420368 152600 420420 152652
rect 421380 152600 421432 152652
rect 138112 152532 138164 152584
rect 144276 152532 144328 152584
rect 144368 152532 144420 152584
rect 226432 152532 226484 152584
rect 234160 152532 234212 152584
rect 297732 152532 297784 152584
rect 304816 152532 304868 152584
rect 351644 152532 351696 152584
rect 352012 152532 352064 152584
rect 388260 152532 388312 152584
rect 388352 152532 388404 152584
rect 392216 152532 392268 152584
rect 393136 152532 393188 152584
rect 419080 152532 419132 152584
rect 419540 152532 419592 152584
rect 419816 152532 419868 152584
rect 421012 152532 421064 152584
rect 423312 152532 423364 152584
rect 423404 152532 423456 152584
rect 434260 152600 434312 152652
rect 436928 152600 436980 152652
rect 437020 152600 437072 152652
rect 438952 152600 439004 152652
rect 440332 152600 440384 152652
rect 455696 152600 455748 152652
rect 2872 152464 2924 152516
rect 121092 152464 121144 152516
rect 126980 152464 127032 152516
rect 216128 152464 216180 152516
rect 227720 152464 227772 152516
rect 293224 152464 293276 152516
rect 298652 152464 298704 152516
rect 347136 152464 347188 152516
rect 347964 152464 348016 152516
rect 385040 152464 385092 152516
rect 386420 152464 386472 152516
rect 413928 152464 413980 152516
rect 414388 152464 414440 152516
rect 67088 152396 67140 152448
rect 159640 152396 159692 152448
rect 173256 152396 173308 152448
rect 249524 152396 249576 152448
rect 251180 152396 251232 152448
rect 311164 152396 311216 152448
rect 317420 152396 317472 152448
rect 361304 152396 361356 152448
rect 365720 152396 365772 152448
rect 398472 152396 398524 152448
rect 398564 152396 398616 152448
rect 408132 152396 408184 152448
rect 412824 152396 412876 152448
rect 120080 152328 120132 152380
rect 211068 152328 211120 152380
rect 224592 152328 224644 152380
rect 288072 152328 288124 152380
rect 292212 152328 292264 152380
rect 341984 152328 342036 152380
rect 343640 152328 343692 152380
rect 349804 152328 349856 152380
rect 349896 152328 349948 152380
rect 385684 152328 385736 152380
rect 385776 152328 385828 152380
rect 387616 152328 387668 152380
rect 389180 152328 389232 152380
rect 412640 152328 412692 152380
rect 415860 152328 415912 152380
rect 426808 152328 426860 152380
rect 426900 152328 426952 152380
rect 432052 152328 432104 152380
rect 433800 152328 433852 152380
rect 440884 152532 440936 152584
rect 442080 152532 442132 152584
rect 456984 152532 457036 152584
rect 459560 152532 459612 152584
rect 464620 152532 464672 152584
rect 442172 152396 442224 152448
rect 434536 152328 434588 152380
rect 434628 152328 434680 152380
rect 437020 152328 437072 152380
rect 437756 152328 437808 152380
rect 91100 152260 91152 152312
rect 180248 152260 180300 152312
rect 187976 152260 188028 152312
rect 262404 152260 262456 152312
rect 266360 152260 266412 152312
rect 320824 152260 320876 152312
rect 325884 152260 325936 152312
rect 367652 152260 367704 152312
rect 371332 152260 371384 152312
rect 402336 152260 402388 152312
rect 404268 152260 404320 152312
rect 405096 152260 405148 152312
rect 409236 152260 409288 152312
rect 417884 152260 417936 152312
rect 419908 152260 419960 152312
rect 428648 152260 428700 152312
rect 429292 152260 429344 152312
rect 438400 152260 438452 152312
rect 109040 152192 109092 152244
rect 130752 152192 130804 152244
rect 134064 152192 134116 152244
rect 221280 152192 221332 152244
rect 221464 152192 221516 152244
rect 282920 152192 282972 152244
rect 285772 152192 285824 152244
rect 336188 152192 336240 152244
rect 342444 152192 342496 152244
rect 344560 152192 344612 152244
rect 349160 152192 349212 152244
rect 349896 152192 349948 152244
rect 354496 152192 354548 152244
rect 389548 152192 389600 152244
rect 394608 152192 394660 152244
rect 417792 152192 417844 152244
rect 419816 152192 419868 152244
rect 421748 152192 421800 152244
rect 422944 152192 422996 152244
rect 429384 152192 429436 152244
rect 429476 152192 429528 152244
rect 431960 152192 432012 152244
rect 432052 152192 432104 152244
rect 438308 152192 438360 152244
rect 438860 152328 438912 152380
rect 454408 152464 454460 152516
rect 444196 152328 444248 152380
rect 452476 152396 452528 152448
rect 444380 152328 444432 152380
rect 453764 152328 453816 152380
rect 511632 152328 511684 152380
rect 513564 152328 513616 152380
rect 438584 152260 438636 152312
rect 446680 152260 446732 152312
rect 441436 152192 441488 152244
rect 441620 152192 441672 152244
rect 456340 152192 456392 152244
rect 513564 152192 513616 152244
rect 516140 152192 516192 152244
rect 82820 152124 82872 152176
rect 169944 152124 169996 152176
rect 172152 152124 172204 152176
rect 190460 152124 190512 152176
rect 194140 152124 194192 152176
rect 213552 152124 213604 152176
rect 79324 152056 79376 152108
rect 164792 152056 164844 152108
rect 167000 152056 167052 152108
rect 182732 152056 182784 152108
rect 183468 152056 183520 152108
rect 200764 152056 200816 152108
rect 212724 152056 212776 152108
rect 274548 152124 274600 152176
rect 277400 152124 277452 152176
rect 331128 152124 331180 152176
rect 332600 152124 332652 152176
rect 372804 152124 372856 152176
rect 384948 152124 385000 152176
rect 392124 152124 392176 152176
rect 392216 152124 392268 152176
rect 407488 152124 407540 152176
rect 408500 152124 408552 152176
rect 423588 152124 423640 152176
rect 423680 152124 423732 152176
rect 427084 152124 427136 152176
rect 427820 152124 427872 152176
rect 225328 152056 225380 152108
rect 229008 152056 229060 152108
rect 243360 152056 243412 152108
rect 302884 152056 302936 152108
rect 303712 152056 303764 152108
rect 351000 152056 351052 152108
rect 354680 152056 354732 152108
rect 390192 152056 390244 152108
rect 398840 152056 398892 152108
rect 68836 151988 68888 152040
rect 142804 151988 142856 152040
rect 143448 151988 143500 152040
rect 146944 151988 146996 152040
rect 156328 151988 156380 152040
rect 172520 151988 172572 152040
rect 191472 151988 191524 152040
rect 208492 151988 208544 152040
rect 242440 151988 242492 152040
rect 300952 151988 301004 152040
rect 307392 151988 307444 152040
rect 352288 151988 352340 152040
rect 364524 151988 364576 152040
rect 397184 151988 397236 152040
rect 75460 151920 75512 151972
rect 154488 151920 154540 151972
rect 162492 151920 162544 151972
rect 177672 151920 177724 151972
rect 184388 151920 184440 151972
rect 195612 151920 195664 151972
rect 213736 151920 213788 151972
rect 272708 151920 272760 151972
rect 272800 151920 272852 151972
rect 325976 151920 326028 151972
rect 331220 151920 331272 151972
rect 372160 151920 372212 151972
rect 378784 151920 378836 151972
rect 384396 151920 384448 151972
rect 388444 151920 388496 151972
rect 404912 151920 404964 151972
rect 405648 152056 405700 152108
rect 421012 152056 421064 152108
rect 405096 151988 405148 152040
rect 418436 151988 418488 152040
rect 419632 151988 419684 152040
rect 434444 152056 434496 152108
rect 434720 152056 434772 152108
rect 435732 152056 435784 152108
rect 436836 152124 436888 152176
rect 443460 152124 443512 152176
rect 445208 152124 445260 152176
rect 445300 152124 445352 152176
rect 458824 152124 458876 152176
rect 444380 152056 444432 152108
rect 449256 152056 449308 152108
rect 425060 151988 425112 152040
rect 436836 151988 436888 152040
rect 436928 151988 436980 152040
rect 444104 151988 444156 152040
rect 444472 151988 444524 152040
rect 458180 151988 458232 152040
rect 467840 151988 467892 152040
rect 471704 151988 471756 152040
rect 485780 151988 485832 152040
rect 490288 151988 490340 152040
rect 516692 151988 516744 152040
rect 520280 151988 520332 152040
rect 413284 151920 413336 151972
rect 417240 151920 417292 151972
rect 431776 151920 431828 151972
rect 431868 151920 431920 151972
rect 439596 151920 439648 151972
rect 440148 151920 440200 151972
rect 26700 151852 26752 151904
rect 71688 151852 71740 151904
rect 109132 151852 109184 151904
rect 33600 151784 33652 151836
rect 82820 151784 82872 151836
rect 105820 151784 105872 151836
rect 110328 151784 110380 151836
rect 110512 151852 110564 151904
rect 138480 151852 138532 151904
rect 139308 151852 139360 151904
rect 203340 151852 203392 151904
rect 260932 151852 260984 151904
rect 316316 151852 316368 151904
rect 321560 151852 321612 151904
rect 362592 151852 362644 151904
rect 363144 151852 363196 151904
rect 364524 151852 364576 151904
rect 386328 151852 386380 151904
rect 394700 151852 394752 151904
rect 396172 151852 396224 151904
rect 402980 151852 403032 151904
rect 404176 151852 404228 151904
rect 128176 151784 128228 151836
rect 129740 151784 129792 151836
rect 146852 151784 146904 151836
rect 146944 151784 146996 151836
rect 157064 151784 157116 151836
rect 169760 151784 169812 151836
rect 185308 151784 185360 151836
rect 283196 151784 283248 151836
rect 287428 151784 287480 151836
rect 299572 151784 299624 151836
rect 346492 151784 346544 151836
rect 349804 151784 349856 151836
rect 380532 151784 380584 151836
rect 398104 151784 398156 151836
rect 405556 151784 405608 151836
rect 413192 151852 413244 151904
rect 415860 151784 415912 151836
rect 418528 151852 418580 151904
rect 426900 151852 426952 151904
rect 421656 151784 421708 151836
rect 421748 151784 421800 151836
rect 437020 151852 437072 151904
rect 437112 151852 437164 151904
rect 443828 151852 443880 151904
rect 444288 151920 444340 151972
rect 451096 151920 451148 151972
rect 451188 151920 451240 151972
rect 457628 151920 457680 151972
rect 469220 151920 469272 151972
rect 472348 151920 472400 151972
rect 487344 151920 487396 151972
rect 490932 151920 490984 151972
rect 509056 151920 509108 151972
rect 510896 151920 510948 151972
rect 515496 151920 515548 151972
rect 518900 151920 518952 151972
rect 444472 151852 444524 151904
rect 427084 151784 427136 151836
rect 431224 151784 431276 151836
rect 431960 151784 432012 151836
rect 441528 151784 441580 151836
rect 441988 151784 442040 151836
rect 444380 151784 444432 151836
rect 441436 151648 441488 151700
rect 451832 151852 451884 151904
rect 464344 151852 464396 151904
rect 467840 151852 467892 151904
rect 467932 151852 467984 151904
rect 471060 151852 471112 151904
rect 488540 151852 488592 151904
rect 492220 151852 492272 151904
rect 507768 151852 507820 151904
rect 509516 151852 509568 151904
rect 516048 151852 516100 151904
rect 519452 151852 519504 151904
rect 445208 151784 445260 151836
rect 446036 151784 446088 151836
rect 488172 151784 488224 151836
rect 491576 151784 491628 151836
rect 499120 151784 499172 151836
rect 499948 151784 500000 151836
rect 517428 151784 517480 151836
rect 521568 151784 521620 151836
rect 82820 151376 82872 151428
rect 117228 151376 117280 151428
rect 68008 151308 68060 151360
rect 112720 151308 112772 151360
rect 71688 151240 71740 151292
rect 117044 151240 117096 151292
rect 64512 151172 64564 151224
rect 112628 151172 112680 151224
rect 61108 151104 61160 151156
rect 112536 151104 112588 151156
rect 57704 151036 57756 151088
rect 111708 151036 111760 151088
rect 54208 150968 54260 151020
rect 112444 150968 112496 151020
rect 50804 150900 50856 150952
rect 111616 150900 111668 150952
rect 47308 150832 47360 150884
rect 111524 150832 111576 150884
rect 43904 150764 43956 150816
rect 111432 150764 111484 150816
rect 40500 150696 40552 150748
rect 111340 150696 111392 150748
rect 37004 150628 37056 150680
rect 111248 150628 111300 150680
rect 23296 150560 23348 150612
rect 116952 150560 117004 150612
rect 12992 150492 13044 150544
rect 116676 150492 116728 150544
rect 2688 150424 2740 150476
rect 111064 150424 111116 150476
rect 263692 150288 263744 150340
rect 122840 150152 122892 150204
rect 123714 150152 123766 150204
rect 146392 150152 146444 150204
rect 147542 150152 147594 150204
rect 164332 150152 164384 150204
rect 165482 150152 165534 150204
rect 168380 150152 168432 150204
rect 169346 150152 169398 150204
rect 171140 150152 171192 150204
rect 171922 150152 171974 150204
rect 172704 150152 172756 150204
rect 173854 150152 173906 150204
rect 182272 150152 182324 150204
rect 183422 150152 183474 150204
rect 211252 150152 211304 150204
rect 212310 150152 212362 150204
rect 225052 150152 225104 150204
rect 225834 150152 225886 150204
rect 229192 150152 229244 150204
rect 230342 150152 230394 150204
rect 233240 150152 233292 150204
rect 234206 150152 234258 150204
rect 238944 150152 238996 150204
rect 240002 150152 240054 150204
rect 253940 150152 253992 150204
rect 254722 150152 254774 150204
rect 256792 150152 256844 150204
rect 257942 150152 257994 150204
rect 264382 150152 264434 150204
rect 269120 150152 269172 150204
rect 270178 150152 270230 150204
rect 281540 150152 281592 150204
rect 282322 150152 282374 150204
rect 283104 150152 283156 150204
rect 284254 150152 284306 150204
rect 284392 150152 284444 150204
rect 285542 150152 285594 150204
rect 299480 150152 299532 150204
rect 300354 150152 300406 150204
rect 321744 150152 321796 150204
rect 322802 150152 322854 150204
rect 328460 150152 328512 150204
rect 329242 150152 329294 150204
rect 332692 150152 332744 150204
rect 333750 150152 333802 150204
rect 338396 150152 338448 150204
rect 339454 150152 339506 150204
rect 345112 150152 345164 150204
rect 345894 150152 345946 150204
rect 358912 150152 358964 150204
rect 360062 150152 360114 150204
rect 362960 150152 363012 150204
rect 363926 150152 363978 150204
rect 375564 150152 375616 150204
rect 376714 150152 376766 150204
rect 378140 150152 378192 150204
rect 379290 150152 379342 150204
rect 394976 150152 395028 150204
rect 396034 150152 396086 150204
rect 462320 150152 462372 150204
rect 463378 150152 463430 150204
rect 477684 150152 477736 150204
rect 478834 150152 478886 150204
rect 478972 150152 479024 150204
rect 480122 150152 480174 150204
rect 481640 150152 481692 150204
rect 482698 150152 482750 150204
rect 483204 150152 483256 150204
rect 483986 150152 484038 150204
rect 518026 150152 518078 150204
rect 518808 150152 518860 150204
rect 102600 150016 102652 150068
rect 116216 150016 116268 150068
rect 20168 149948 20220 150000
rect 116860 149948 116912 150000
rect 16488 149880 16540 149932
rect 116768 149880 116820 149932
rect 9588 149812 9640 149864
rect 116584 149812 116636 149864
rect 6368 149744 6420 149796
rect 111156 149744 111208 149796
rect 85488 149676 85540 149728
rect 112352 149676 112404 149728
rect 81992 149608 82044 149660
rect 113088 149608 113140 149660
rect 78588 149540 78640 149592
rect 112996 149540 113048 149592
rect 75184 149472 75236 149524
rect 112904 149472 112956 149524
rect 71688 149404 71740 149456
rect 112812 149404 112864 149456
rect 30288 149336 30340 149388
rect 117136 149336 117188 149388
rect 88984 149268 89036 149320
rect 92020 149200 92072 149252
rect 95792 149268 95844 149320
rect 99288 149268 99340 149320
rect 116032 149268 116084 149320
rect 116400 149200 116452 149252
rect 116492 149132 116544 149184
rect 112260 149064 112312 149116
rect 109592 148996 109644 149048
rect 116124 148996 116176 149048
rect 110328 147568 110380 147620
rect 116124 147568 116176 147620
rect 112260 140700 112312 140752
rect 116124 140700 116176 140752
rect 112352 136552 112404 136604
rect 116124 136552 116176 136604
rect 113088 133832 113140 133884
rect 116032 133832 116084 133884
rect 114192 132608 114244 132660
rect 115204 132608 115256 132660
rect 112996 132404 113048 132456
rect 116124 132404 116176 132456
rect 112904 131044 112956 131096
rect 116124 131044 116176 131096
rect 112812 128256 112864 128308
rect 116124 128256 116176 128308
rect 112720 126896 112772 126948
rect 116032 126896 116084 126948
rect 112628 124108 112680 124160
rect 116124 124108 116176 124160
rect 112536 122748 112588 122800
rect 115940 122748 115992 122800
rect 111708 121388 111760 121440
rect 116124 121388 116176 121440
rect 112444 118600 112496 118652
rect 116124 118600 116176 118652
rect 116492 117988 116544 118040
rect 117228 117988 117280 118040
rect 111616 117240 111668 117292
rect 116124 117240 116176 117292
rect 111524 114452 111576 114504
rect 116124 114452 116176 114504
rect 111432 113092 111484 113144
rect 115940 113092 115992 113144
rect 111340 111732 111392 111784
rect 116124 111732 116176 111784
rect 111248 108944 111300 108996
rect 116124 108944 116176 108996
rect 111156 92420 111208 92472
rect 116124 92420 116176 92472
rect 111064 89632 111116 89684
rect 116124 89632 116176 89684
rect 113824 88272 113876 88324
rect 116032 88272 116084 88324
rect 114468 87184 114520 87236
rect 116492 87184 116544 87236
rect 113916 83920 113968 83972
rect 116584 83920 116636 83972
rect 114008 82764 114060 82816
rect 116216 82764 116268 82816
rect 114100 79976 114152 80028
rect 115940 79976 115992 80028
rect 114192 71748 114244 71800
rect 116584 71748 116636 71800
rect 114100 69028 114152 69080
rect 116308 69028 116360 69080
rect 114008 67600 114060 67652
rect 116124 67600 116176 67652
rect 113916 66240 113968 66292
rect 116584 66240 116636 66292
rect 114468 64540 114520 64592
rect 116584 64540 116636 64592
rect 113824 63520 113876 63572
rect 116216 63520 116268 63572
rect 109684 41420 109736 41472
rect 116124 41420 116176 41472
rect 114100 38632 114152 38684
rect 116400 38632 116452 38684
rect 116216 38496 116268 38548
rect 116400 38496 116452 38548
rect 114192 37272 114244 37324
rect 116216 37272 116268 37324
rect 111064 34484 111116 34536
rect 116124 34484 116176 34536
rect 112444 33124 112496 33176
rect 116124 33124 116176 33176
rect 112536 31764 112588 31816
rect 116124 31764 116176 31816
rect 112628 28976 112680 29028
rect 116124 28976 116176 29028
rect 112720 27616 112772 27668
rect 116124 27616 116176 27668
rect 112812 24828 112864 24880
rect 116124 24828 116176 24880
rect 111156 23468 111208 23520
rect 116124 23468 116176 23520
rect 111248 22108 111300 22160
rect 116032 22108 116084 22160
rect 116032 16464 116084 16516
rect 116216 16464 116268 16516
rect 116216 11840 116268 11892
rect 116308 11636 116360 11688
rect 116952 11364 117004 11416
rect 117320 11364 117372 11416
rect 116952 5448 117004 5500
rect 117136 5448 117188 5500
rect 116308 5312 116360 5364
rect 116952 5312 117004 5364
rect 115940 5176 115992 5228
rect 116308 5176 116360 5228
rect 115940 5040 115992 5092
rect 116124 5040 116176 5092
rect 109776 4156 109828 4208
rect 116124 4156 116176 4208
rect 2504 2592 2556 2644
rect 39396 2592 39448 2644
rect 39764 2592 39816 2644
rect 42984 2592 43036 2644
rect 43536 2592 43588 2644
rect 46112 2592 46164 2644
rect 50620 2592 50672 2644
rect 53656 2592 53708 2644
rect 111064 3884 111116 3936
rect 112444 3816 112496 3868
rect 58716 2592 58768 2644
rect 58808 2592 58860 2644
rect 62856 2592 62908 2644
rect 32772 2456 32824 2508
rect 43536 2456 43588 2508
rect 58624 2524 58676 2576
rect 59728 2524 59780 2576
rect 112536 3748 112588 3800
rect 112628 3680 112680 3732
rect 112720 3612 112772 3664
rect 112812 3544 112864 3596
rect 111156 3476 111208 3528
rect 63316 2592 63368 2644
rect 63500 2592 63552 2644
rect 66996 2592 67048 2644
rect 68008 2592 68060 2644
rect 80152 2592 80204 2644
rect 80244 2592 80296 2644
rect 80336 2592 80388 2644
rect 80428 2592 80480 2644
rect 81532 2592 81584 2644
rect 81624 2592 81676 2644
rect 81808 2592 81860 2644
rect 81900 2592 81952 2644
rect 81992 2592 82044 2644
rect 82452 2592 82504 2644
rect 111248 3408 111300 3460
rect 114192 3340 114244 3392
rect 114100 3272 114152 3324
rect 112444 3204 112496 3256
rect 82728 2592 82780 2644
rect 73252 2524 73304 2576
rect 82360 2524 82412 2576
rect 73068 2456 73120 2508
rect 73344 2456 73396 2508
rect 82268 2456 82320 2508
rect 36360 2388 36412 2440
rect 39764 2388 39816 2440
rect 50620 2388 50672 2440
rect 56140 2388 56192 2440
rect 58624 2388 58676 2440
rect 68008 2388 68060 2440
rect 80152 2388 80204 2440
rect 81900 2388 81952 2440
rect 83004 2592 83056 2644
rect 83096 2592 83148 2644
rect 52920 2320 52972 2372
rect 66996 2320 67048 2372
rect 69664 2320 69716 2372
rect 82268 2320 82320 2372
rect 117964 3000 118016 3052
rect 112444 2932 112496 2984
rect 117688 2932 117740 2984
rect 98368 2592 98420 2644
rect 98460 2592 98512 2644
rect 100024 2592 100076 2644
rect 116124 2864 116176 2916
rect 98368 2456 98420 2508
rect 100024 2456 100076 2508
rect 109592 2456 109644 2508
rect 116584 2456 116636 2508
rect 294788 2456 294840 2508
rect 425796 2456 425848 2508
rect 443644 2456 443696 2508
rect 106188 2388 106240 2440
rect 116676 2388 116728 2440
rect 102968 2320 103020 2372
rect 116768 2320 116820 2372
rect 49608 2252 49660 2304
rect 58808 2252 58860 2304
rect 81992 2252 82044 2304
rect 99656 2252 99708 2304
rect 116860 2252 116912 2304
rect 56232 2184 56284 2236
rect 73068 2184 73120 2236
rect 80244 2184 80296 2236
rect 81532 2184 81584 2236
rect 82084 2184 82136 2236
rect 82452 2184 82504 2236
rect 96344 2184 96396 2236
rect 117044 2184 117096 2236
rect 63316 2116 63368 2168
rect 80336 2116 80388 2168
rect 81808 2116 81860 2168
rect 93032 2116 93084 2168
rect 117228 2116 117280 2168
rect 80428 2048 80480 2100
rect 81624 2048 81676 2100
rect 89628 2048 89680 2100
rect 117320 2048 117372 2100
rect 86408 1980 86460 2032
rect 117136 1980 117188 2032
rect 82636 1912 82688 1964
rect 116492 1912 116544 1964
rect 79324 1844 79376 1896
rect 116400 1844 116452 1896
rect 72700 1776 72752 1828
rect 109684 1776 109736 1828
rect 76012 1708 76064 1760
rect 116216 1708 116268 1760
rect 32680 1640 32732 1692
rect 116032 1640 116084 1692
rect 29276 1572 29328 1624
rect 115940 1572 115992 1624
rect 25964 1504 26016 1556
rect 116952 1504 117004 1556
rect 22652 1436 22704 1488
rect 116308 1436 116360 1488
rect 117688 1436 117740 1488
rect 143632 1436 143684 1488
rect 6000 1368 6052 1420
rect 109776 1368 109828 1420
rect 117964 1368 118016 1420
rect 193588 1368 193640 1420
rect 294788 1368 294840 1420
rect 343640 1368 343692 1420
rect 491300 1368 491352 1420
rect 493600 1368 493652 1420
<< metal2 >>
rect 386 163200 442 164400
rect 492 163254 1164 163282
rect 400 158030 428 163200
rect 388 158024 440 158030
rect 388 157966 440 157972
rect 492 153882 520 163254
rect 1136 163146 1164 163254
rect 1214 163200 1270 164400
rect 2042 163200 2098 164400
rect 2870 163200 2926 164400
rect 2976 163254 3648 163282
rect 1228 163146 1256 163200
rect 1136 163118 1256 163146
rect 2056 156670 2084 163200
rect 2044 156664 2096 156670
rect 2044 156606 2096 156612
rect 480 153876 532 153882
rect 480 153818 532 153824
rect 2884 152522 2912 163200
rect 2976 153785 3004 163254
rect 3620 163146 3648 163254
rect 3698 163200 3754 164400
rect 4526 163200 4582 164400
rect 5354 163200 5410 164400
rect 6274 163200 6330 164400
rect 7102 163200 7158 164400
rect 7930 163200 7986 164400
rect 8758 163200 8814 164400
rect 8864 163254 9536 163282
rect 3712 163146 3740 163200
rect 3620 163118 3740 163146
rect 4540 155310 4568 163200
rect 4528 155304 4580 155310
rect 4528 155246 4580 155252
rect 5368 155242 5396 163200
rect 6288 159390 6316 163200
rect 6276 159384 6328 159390
rect 6276 159326 6328 159332
rect 5356 155236 5408 155242
rect 5356 155178 5408 155184
rect 7116 153950 7144 163200
rect 7944 155378 7972 163200
rect 8772 155446 8800 163200
rect 8760 155440 8812 155446
rect 8760 155382 8812 155388
rect 7932 155372 7984 155378
rect 7932 155314 7984 155320
rect 7104 153944 7156 153950
rect 7104 153886 7156 153892
rect 2962 153776 3018 153785
rect 2962 153711 3018 153720
rect 2872 152516 2924 152522
rect 2872 152458 2924 152464
rect 8864 152425 8892 163254
rect 9508 163146 9536 163254
rect 9586 163200 9642 164400
rect 9692 163254 10364 163282
rect 9600 163146 9628 163200
rect 9508 163118 9628 163146
rect 9692 154018 9720 163254
rect 10336 163146 10364 163254
rect 10414 163200 10470 164400
rect 11242 163200 11298 164400
rect 12162 163200 12218 164400
rect 12452 163254 12940 163282
rect 10428 163146 10456 163200
rect 10336 163118 10456 163146
rect 11256 156738 11284 163200
rect 11244 156732 11296 156738
rect 11244 156674 11296 156680
rect 12176 155786 12204 163200
rect 12164 155780 12216 155786
rect 12164 155722 12216 155728
rect 9680 154012 9732 154018
rect 9680 153954 9732 153960
rect 12452 152561 12480 163254
rect 12912 163146 12940 163254
rect 12990 163200 13046 164400
rect 13818 163200 13874 164400
rect 14646 163200 14702 164400
rect 15474 163200 15530 164400
rect 16302 163200 16358 164400
rect 16592 163254 17080 163282
rect 13004 163146 13032 163200
rect 12912 163118 13032 163146
rect 13832 154086 13860 163200
rect 14660 156806 14688 163200
rect 14648 156800 14700 156806
rect 14648 156742 14700 156748
rect 15488 154970 15516 163200
rect 16316 159361 16344 163200
rect 16302 159352 16358 159361
rect 16302 159287 16358 159296
rect 15476 154964 15528 154970
rect 15476 154906 15528 154912
rect 13820 154080 13872 154086
rect 13820 154022 13872 154028
rect 16592 153921 16620 163254
rect 17052 163146 17080 163254
rect 17130 163200 17186 164400
rect 18050 163200 18106 164400
rect 18878 163200 18934 164400
rect 19352 163254 19656 163282
rect 17144 163146 17172 163200
rect 17052 163118 17172 163146
rect 18064 156874 18092 163200
rect 18892 159730 18920 163200
rect 18880 159724 18932 159730
rect 18880 159666 18932 159672
rect 18052 156868 18104 156874
rect 18052 156810 18104 156816
rect 16578 153912 16634 153921
rect 16578 153847 16634 153856
rect 19352 152590 19380 163254
rect 19628 163146 19656 163254
rect 19706 163200 19762 164400
rect 19904 163254 20484 163282
rect 19720 163146 19748 163200
rect 19628 163118 19748 163146
rect 19904 154057 19932 163254
rect 20456 163146 20484 163254
rect 20534 163200 20590 164400
rect 21362 163200 21418 164400
rect 22190 163200 22246 164400
rect 23018 163200 23074 164400
rect 23492 163254 23888 163282
rect 20548 163146 20576 163200
rect 20456 163118 20576 163146
rect 21376 156942 21404 163200
rect 21364 156936 21416 156942
rect 21364 156878 21416 156884
rect 19890 154048 19946 154057
rect 19890 153983 19946 153992
rect 22204 152658 22232 163200
rect 23032 159497 23060 163200
rect 23018 159488 23074 159497
rect 23018 159423 23074 159432
rect 23492 154154 23520 163254
rect 23860 163146 23888 163254
rect 23938 163200 23994 164400
rect 24766 163200 24822 164400
rect 25594 163200 25650 164400
rect 26422 163200 26478 164400
rect 27250 163200 27306 164400
rect 28078 163200 28134 164400
rect 28184 163254 28856 163282
rect 23952 163146 23980 163200
rect 23860 163118 23980 163146
rect 24780 157010 24808 163200
rect 25608 160002 25636 163200
rect 25596 159996 25648 160002
rect 25596 159938 25648 159944
rect 24768 157004 24820 157010
rect 24768 156946 24820 156952
rect 23480 154148 23532 154154
rect 23480 154090 23532 154096
rect 26436 152794 26464 163200
rect 27264 154222 27292 163200
rect 28092 156777 28120 163200
rect 28078 156768 28134 156777
rect 28078 156703 28134 156712
rect 27252 154216 27304 154222
rect 27252 154158 27304 154164
rect 26424 152788 26476 152794
rect 26424 152730 26476 152736
rect 28184 152726 28212 163254
rect 28828 163146 28856 163254
rect 28906 163200 28962 164400
rect 29826 163200 29882 164400
rect 30392 163254 30604 163282
rect 28920 163146 28948 163200
rect 28828 163118 28948 163146
rect 29840 159633 29868 163200
rect 29826 159624 29882 159633
rect 29826 159559 29882 159568
rect 30392 154193 30420 163254
rect 30576 163146 30604 163254
rect 30654 163200 30710 164400
rect 31482 163200 31538 164400
rect 32310 163200 32366 164400
rect 33138 163200 33194 164400
rect 33966 163200 34022 164400
rect 34532 163254 34744 163282
rect 30668 163146 30696 163200
rect 30576 163118 30696 163146
rect 31496 156641 31524 163200
rect 32324 159458 32352 163200
rect 32312 159452 32364 159458
rect 32312 159394 32364 159400
rect 31482 156632 31538 156641
rect 31482 156567 31538 156576
rect 30378 154184 30434 154193
rect 30378 154119 30434 154128
rect 33152 152862 33180 163200
rect 33980 158001 34008 163200
rect 33966 157992 34022 158001
rect 33966 157927 34022 157936
rect 34532 154358 34560 163254
rect 34716 163146 34744 163254
rect 34794 163200 34850 164400
rect 35714 163200 35770 164400
rect 36542 163200 36598 164400
rect 37370 163200 37426 164400
rect 37936 163254 38148 163282
rect 34808 163146 34836 163200
rect 34716 163118 34836 163146
rect 35728 157078 35756 163200
rect 36556 159526 36584 163200
rect 36544 159520 36596 159526
rect 36544 159462 36596 159468
rect 37384 158098 37412 163200
rect 37372 158092 37424 158098
rect 37372 158034 37424 158040
rect 35716 157072 35768 157078
rect 35716 157014 35768 157020
rect 34520 154352 34572 154358
rect 34520 154294 34572 154300
rect 37936 154290 37964 163254
rect 38120 163146 38148 163254
rect 38198 163200 38254 164400
rect 39026 163200 39082 164400
rect 39854 163200 39910 164400
rect 40682 163200 40738 164400
rect 41602 163200 41658 164400
rect 42430 163200 42486 164400
rect 43258 163200 43314 164400
rect 44086 163200 44142 164400
rect 44192 163254 44864 163282
rect 38212 163146 38240 163200
rect 38120 163118 38240 163146
rect 39040 157146 39068 163200
rect 39028 157140 39080 157146
rect 39028 157082 39080 157088
rect 39868 155582 39896 163200
rect 40696 158273 40724 163200
rect 40682 158264 40738 158273
rect 40682 158199 40738 158208
rect 39856 155576 39908 155582
rect 39856 155518 39908 155524
rect 37924 154284 37976 154290
rect 37924 154226 37976 154232
rect 41616 153270 41644 163200
rect 42444 157214 42472 163200
rect 43272 159594 43300 163200
rect 43260 159588 43312 159594
rect 43260 159530 43312 159536
rect 44100 158137 44128 163200
rect 44086 158128 44142 158137
rect 44086 158063 44142 158072
rect 42432 157208 42484 157214
rect 42432 157150 42484 157156
rect 44192 154494 44220 163254
rect 44836 163146 44864 163254
rect 44914 163200 44970 164400
rect 45742 163200 45798 164400
rect 46570 163200 46626 164400
rect 47490 163200 47546 164400
rect 48318 163200 48374 164400
rect 49146 163200 49202 164400
rect 49974 163200 50030 164400
rect 50802 163200 50858 164400
rect 51092 163254 51580 163282
rect 44928 163146 44956 163200
rect 44836 163118 44956 163146
rect 45756 157282 45784 163200
rect 45744 157276 45796 157282
rect 45744 157218 45796 157224
rect 46584 155718 46612 163200
rect 47504 158166 47532 163200
rect 47492 158160 47544 158166
rect 47492 158102 47544 158108
rect 46572 155712 46624 155718
rect 46572 155654 46624 155660
rect 48332 154562 48360 163200
rect 49160 157350 49188 163200
rect 49988 159662 50016 163200
rect 49976 159656 50028 159662
rect 49976 159598 50028 159604
rect 50816 158234 50844 163200
rect 50804 158228 50856 158234
rect 50804 158170 50856 158176
rect 49148 157344 49200 157350
rect 49148 157286 49200 157292
rect 48320 154556 48372 154562
rect 48320 154498 48372 154504
rect 44180 154488 44232 154494
rect 44180 154430 44232 154436
rect 51092 153814 51120 163254
rect 51552 163146 51580 163254
rect 51630 163200 51686 164400
rect 52458 163200 52514 164400
rect 53378 163200 53434 164400
rect 54206 163200 54262 164400
rect 54312 163254 54984 163282
rect 51644 163146 51672 163200
rect 51552 163118 51672 163146
rect 52472 156602 52500 163200
rect 52460 156596 52512 156602
rect 52460 156538 52512 156544
rect 53392 155650 53420 163200
rect 54220 158302 54248 163200
rect 54208 158296 54260 158302
rect 54208 158238 54260 158244
rect 53380 155644 53432 155650
rect 53380 155586 53432 155592
rect 54312 154329 54340 163254
rect 54956 163146 54984 163254
rect 55034 163200 55090 164400
rect 55862 163200 55918 164400
rect 56690 163200 56746 164400
rect 57518 163200 57574 164400
rect 57992 163254 58296 163282
rect 55048 163146 55076 163200
rect 54956 163118 55076 163146
rect 55876 156913 55904 163200
rect 56704 159798 56732 163200
rect 56692 159792 56744 159798
rect 56692 159734 56744 159740
rect 57532 158409 57560 163200
rect 57518 158400 57574 158409
rect 57518 158335 57574 158344
rect 55862 156904 55918 156913
rect 55862 156839 55918 156848
rect 54298 154320 54354 154329
rect 54298 154255 54354 154264
rect 51080 153808 51132 153814
rect 51080 153750 51132 153756
rect 57992 153678 58020 163254
rect 58268 163146 58296 163254
rect 58346 163200 58402 164400
rect 59266 163200 59322 164400
rect 60094 163200 60150 164400
rect 60922 163200 60978 164400
rect 61120 163254 61700 163282
rect 58360 163146 58388 163200
rect 58268 163118 58388 163146
rect 59280 156534 59308 163200
rect 59268 156528 59320 156534
rect 59268 156470 59320 156476
rect 60108 155854 60136 163200
rect 60936 158370 60964 163200
rect 60924 158364 60976 158370
rect 60924 158306 60976 158312
rect 60096 155848 60148 155854
rect 60096 155790 60148 155796
rect 61120 153746 61148 163254
rect 61672 163146 61700 163254
rect 61750 163200 61806 164400
rect 62578 163200 62634 164400
rect 63406 163200 63462 164400
rect 64234 163200 64290 164400
rect 65154 163200 65210 164400
rect 65982 163200 66038 164400
rect 66810 163200 66866 164400
rect 67638 163200 67694 164400
rect 68466 163200 68522 164400
rect 69294 163200 69350 164400
rect 70122 163200 70178 164400
rect 71042 163200 71098 164400
rect 71870 163200 71926 164400
rect 72698 163200 72754 164400
rect 73526 163200 73582 164400
rect 74354 163200 74410 164400
rect 75182 163200 75238 164400
rect 76010 163200 76066 164400
rect 76930 163200 76986 164400
rect 77758 163200 77814 164400
rect 78586 163200 78642 164400
rect 78692 163254 79364 163282
rect 61764 163146 61792 163200
rect 61672 163118 61792 163146
rect 62592 155553 62620 163200
rect 63420 160070 63448 163200
rect 63408 160064 63460 160070
rect 63408 160006 63460 160012
rect 64248 158438 64276 163200
rect 64236 158432 64288 158438
rect 64236 158374 64288 158380
rect 62578 155544 62634 155553
rect 65168 155514 65196 163200
rect 62578 155479 62634 155488
rect 65156 155508 65208 155514
rect 65156 155450 65208 155456
rect 65996 155417 66024 163200
rect 66824 155922 66852 163200
rect 67652 158642 67680 163200
rect 67640 158636 67692 158642
rect 67640 158578 67692 158584
rect 66812 155916 66864 155922
rect 66812 155858 66864 155864
rect 67088 155644 67140 155650
rect 67088 155586 67140 155592
rect 65982 155408 66038 155417
rect 65982 155343 66038 155352
rect 61108 153740 61160 153746
rect 61108 153682 61160 153688
rect 57980 153672 58032 153678
rect 57980 153614 58032 153620
rect 41604 153264 41656 153270
rect 41604 153206 41656 153212
rect 33140 152856 33192 152862
rect 33140 152798 33192 152804
rect 28172 152720 28224 152726
rect 28172 152662 28224 152668
rect 22192 152652 22244 152658
rect 22192 152594 22244 152600
rect 19340 152584 19392 152590
rect 12438 152552 12494 152561
rect 19340 152526 19392 152532
rect 12438 152487 12494 152496
rect 67100 152454 67128 155586
rect 68480 155281 68508 163200
rect 69308 156466 69336 163200
rect 70136 159866 70164 163200
rect 70124 159860 70176 159866
rect 70124 159802 70176 159808
rect 71056 158506 71084 163200
rect 71044 158500 71096 158506
rect 71044 158442 71096 158448
rect 69296 156460 69348 156466
rect 69296 156402 69348 156408
rect 71884 155650 71912 163200
rect 72712 157049 72740 163200
rect 73540 159322 73568 163200
rect 73528 159316 73580 159322
rect 73528 159258 73580 159264
rect 74368 158574 74396 163200
rect 74356 158568 74408 158574
rect 74356 158510 74408 158516
rect 72698 157040 72754 157049
rect 72698 156975 72754 156984
rect 71872 155644 71924 155650
rect 71872 155586 71924 155592
rect 75196 155582 75224 163200
rect 76024 155825 76052 163200
rect 76944 159934 76972 163200
rect 76932 159928 76984 159934
rect 76932 159870 76984 159876
rect 77772 157962 77800 163200
rect 77760 157956 77812 157962
rect 77760 157898 77812 157904
rect 76010 155816 76066 155825
rect 76010 155751 76066 155760
rect 75460 155712 75512 155718
rect 78600 155689 78628 163200
rect 75460 155654 75512 155660
rect 78586 155680 78642 155689
rect 68836 155576 68888 155582
rect 68836 155518 68888 155524
rect 75184 155576 75236 155582
rect 75184 155518 75236 155524
rect 68466 155272 68522 155281
rect 68466 155207 68522 155216
rect 67088 152448 67140 152454
rect 8850 152416 8906 152425
rect 67088 152390 67140 152396
rect 8850 152351 8906 152360
rect 68848 152046 68876 155518
rect 68836 152040 68888 152046
rect 68836 151982 68888 151988
rect 75472 151978 75500 155654
rect 78586 155615 78642 155624
rect 78692 153610 78720 163254
rect 79336 163146 79364 163254
rect 79414 163200 79470 164400
rect 80242 163200 80298 164400
rect 81070 163200 81126 164400
rect 81898 163200 81954 164400
rect 82818 163200 82874 164400
rect 83646 163200 83702 164400
rect 84474 163200 84530 164400
rect 85302 163200 85358 164400
rect 85592 163254 86080 163282
rect 79428 163146 79456 163200
rect 79336 163118 79456 163146
rect 80060 159316 80112 159322
rect 80060 159258 80112 159264
rect 79324 155848 79376 155854
rect 79324 155790 79376 155796
rect 78680 153604 78732 153610
rect 78680 153546 78732 153552
rect 79336 152114 79364 155790
rect 80072 153134 80100 159258
rect 80256 159254 80284 163200
rect 80244 159248 80296 159254
rect 80244 159190 80296 159196
rect 81084 158710 81112 163200
rect 81072 158704 81124 158710
rect 81072 158646 81124 158652
rect 81912 155718 81940 163200
rect 82832 156398 82860 163200
rect 83660 159322 83688 163200
rect 83648 159316 83700 159322
rect 83648 159258 83700 159264
rect 84488 157826 84516 163200
rect 84476 157820 84528 157826
rect 84476 157762 84528 157768
rect 82820 156392 82872 156398
rect 82820 156334 82872 156340
rect 85316 155961 85344 163200
rect 85302 155952 85358 155961
rect 82820 155916 82872 155922
rect 85302 155887 85358 155896
rect 82820 155858 82872 155864
rect 81900 155712 81952 155718
rect 81900 155654 81952 155660
rect 80060 153128 80112 153134
rect 80060 153070 80112 153076
rect 82832 152182 82860 155858
rect 85592 154465 85620 163254
rect 86052 163146 86080 163254
rect 86130 163200 86186 164400
rect 86958 163200 87014 164400
rect 87786 163200 87842 164400
rect 88706 163200 88762 164400
rect 89534 163200 89590 164400
rect 90362 163200 90418 164400
rect 91190 163200 91246 164400
rect 92018 163200 92074 164400
rect 92846 163200 92902 164400
rect 93674 163200 93730 164400
rect 94594 163200 94650 164400
rect 95422 163200 95478 164400
rect 96250 163200 96306 164400
rect 96632 163254 97028 163282
rect 86144 163146 86172 163200
rect 86052 163118 86172 163146
rect 86972 159186 87000 163200
rect 86960 159180 87012 159186
rect 86960 159122 87012 159128
rect 87800 157894 87828 163200
rect 87788 157888 87840 157894
rect 87788 157830 87840 157836
rect 88720 155854 88748 163200
rect 89548 155922 89576 163200
rect 90376 158778 90404 163200
rect 91100 159248 91152 159254
rect 91100 159190 91152 159196
rect 90364 158772 90416 158778
rect 90364 158714 90416 158720
rect 89536 155916 89588 155922
rect 89536 155858 89588 155864
rect 88708 155848 88760 155854
rect 88708 155790 88760 155796
rect 85578 154456 85634 154465
rect 85578 154391 85634 154400
rect 91112 152318 91140 159190
rect 91204 157758 91232 163200
rect 91192 157752 91244 157758
rect 91192 157694 91244 157700
rect 92032 155174 92060 163200
rect 92860 158778 92888 163200
rect 93688 159118 93716 163200
rect 93676 159112 93728 159118
rect 93676 159054 93728 159060
rect 92480 158772 92532 158778
rect 92480 158714 92532 158720
rect 92848 158772 92900 158778
rect 92848 158714 92900 158720
rect 92020 155168 92072 155174
rect 92020 155110 92072 155116
rect 92492 152998 92520 158714
rect 94608 157690 94636 163200
rect 94596 157684 94648 157690
rect 94596 157626 94648 157632
rect 95436 155106 95464 163200
rect 96264 158982 96292 163200
rect 96252 158976 96304 158982
rect 96252 158918 96304 158924
rect 95424 155100 95476 155106
rect 95424 155042 95476 155048
rect 92480 152992 92532 152998
rect 92480 152934 92532 152940
rect 96632 152930 96660 163254
rect 97000 163146 97028 163254
rect 97078 163200 97134 164400
rect 97906 163200 97962 164400
rect 98734 163200 98790 164400
rect 99562 163200 99618 164400
rect 100482 163200 100538 164400
rect 101310 163200 101366 164400
rect 102138 163200 102194 164400
rect 102966 163200 103022 164400
rect 103532 163254 103744 163282
rect 97092 163146 97120 163200
rect 97000 163118 97120 163146
rect 97920 157622 97948 163200
rect 97908 157616 97960 157622
rect 97908 157558 97960 157564
rect 98748 155038 98776 163200
rect 99576 156330 99604 163200
rect 100496 159254 100524 163200
rect 100484 159248 100536 159254
rect 100484 159190 100536 159196
rect 99564 156324 99616 156330
rect 99564 156266 99616 156272
rect 101324 156262 101352 163200
rect 101312 156256 101364 156262
rect 101312 156198 101364 156204
rect 98736 155032 98788 155038
rect 98736 154974 98788 154980
rect 102152 153542 102180 163200
rect 102980 158914 103008 163200
rect 102968 158908 103020 158914
rect 102968 158850 103020 158856
rect 102140 153536 102192 153542
rect 102140 153478 102192 153484
rect 103532 153066 103560 163254
rect 103716 163146 103744 163254
rect 103794 163200 103850 164400
rect 104622 163200 104678 164400
rect 104912 163254 105400 163282
rect 103808 163146 103836 163200
rect 103716 163118 103836 163146
rect 104636 158545 104664 163200
rect 104622 158536 104678 158545
rect 104622 158471 104678 158480
rect 104912 153474 104940 163254
rect 105372 163146 105400 163254
rect 105450 163200 105506 164400
rect 106370 163200 106426 164400
rect 107198 163200 107254 164400
rect 108026 163200 108082 164400
rect 108316 163254 108804 163282
rect 105464 163146 105492 163200
rect 105372 163118 105492 163146
rect 106384 154902 106412 163200
rect 107212 159050 107240 163200
rect 107200 159044 107252 159050
rect 107200 158986 107252 158992
rect 108040 156194 108068 163200
rect 108028 156188 108080 156194
rect 108028 156130 108080 156136
rect 106372 154896 106424 154902
rect 106372 154838 106424 154844
rect 104900 153468 104952 153474
rect 104900 153410 104952 153416
rect 108316 153406 108344 163254
rect 108776 163146 108804 163254
rect 108854 163200 108910 164400
rect 109682 163200 109738 164400
rect 110510 163200 110566 164400
rect 111338 163200 111394 164400
rect 112258 163200 112314 164400
rect 113086 163200 113142 164400
rect 113192 163254 113864 163282
rect 108868 163146 108896 163200
rect 108776 163118 108896 163146
rect 109224 159724 109276 159730
rect 109224 159666 109276 159672
rect 109132 155780 109184 155786
rect 109132 155722 109184 155728
rect 109040 154964 109092 154970
rect 109040 154906 109092 154912
rect 108304 153400 108356 153406
rect 108304 153342 108356 153348
rect 103520 153060 103572 153066
rect 103520 153002 103572 153008
rect 96620 152924 96672 152930
rect 96620 152866 96672 152872
rect 91100 152312 91152 152318
rect 91100 152254 91152 152260
rect 109052 152250 109080 154906
rect 109040 152244 109092 152250
rect 109040 152186 109092 152192
rect 82820 152176 82872 152182
rect 82820 152118 82872 152124
rect 79324 152108 79376 152114
rect 79324 152050 79376 152056
rect 75460 151972 75512 151978
rect 75460 151914 75512 151920
rect 109144 151910 109172 155722
rect 109236 154766 109264 159666
rect 109696 158846 109724 163200
rect 110328 159996 110380 160002
rect 110328 159938 110380 159944
rect 109684 158840 109736 158846
rect 109684 158782 109736 158788
rect 109224 154760 109276 154766
rect 109224 154702 109276 154708
rect 110340 151994 110368 159938
rect 110524 154834 110552 163200
rect 111352 157554 111380 163200
rect 111340 157548 111392 157554
rect 111340 157490 111392 157496
rect 112272 155786 112300 163200
rect 113100 159730 113128 163200
rect 113088 159724 113140 159730
rect 113088 159666 113140 159672
rect 112260 155780 112312 155786
rect 112260 155722 112312 155728
rect 110512 154828 110564 154834
rect 110512 154770 110564 154776
rect 113192 153202 113220 163254
rect 113836 163146 113864 163254
rect 113914 163200 113970 164400
rect 114742 163200 114798 164400
rect 115570 163200 115626 164400
rect 115952 163254 116348 163282
rect 113928 163146 113956 163200
rect 113836 163118 113956 163146
rect 114468 158772 114520 158778
rect 114468 158714 114520 158720
rect 114480 154426 114508 158714
rect 114756 157486 114784 163200
rect 114744 157480 114796 157486
rect 114744 157422 114796 157428
rect 115584 157185 115612 163200
rect 115570 157176 115626 157185
rect 115570 157111 115626 157120
rect 114468 154420 114520 154426
rect 114468 154362 114520 154368
rect 115952 153338 115980 163254
rect 116320 163146 116348 163254
rect 116398 163200 116454 164400
rect 117226 163200 117282 164400
rect 118146 163200 118202 164400
rect 118712 163254 118924 163282
rect 116412 163146 116440 163200
rect 116320 163118 116440 163146
rect 117240 160002 117268 163200
rect 117228 159996 117280 160002
rect 117228 159938 117280 159944
rect 118160 156126 118188 163200
rect 118148 156120 118200 156126
rect 118148 156062 118200 156068
rect 118608 154624 118660 154630
rect 118608 154566 118660 154572
rect 118620 154426 118648 154566
rect 118712 154426 118740 163254
rect 118896 163146 118924 163254
rect 118974 163200 119030 164400
rect 119802 163200 119858 164400
rect 120092 163254 120580 163282
rect 118988 163146 119016 163200
rect 118896 163118 119016 163146
rect 119816 158778 119844 163200
rect 119804 158772 119856 158778
rect 119804 158714 119856 158720
rect 118884 158024 118936 158030
rect 118884 157966 118936 157972
rect 118608 154420 118660 154426
rect 118608 154362 118660 154368
rect 118700 154420 118752 154426
rect 118700 154362 118752 154368
rect 115940 153332 115992 153338
rect 115940 153274 115992 153280
rect 113180 153196 113232 153202
rect 113180 153138 113232 153144
rect 110340 151966 110552 151994
rect 110524 151910 110552 151966
rect 26700 151904 26752 151910
rect 26700 151846 26752 151852
rect 71688 151904 71740 151910
rect 71688 151846 71740 151852
rect 109132 151904 109184 151910
rect 109132 151846 109184 151852
rect 110512 151904 110564 151910
rect 110512 151846 110564 151852
rect 23296 150612 23348 150618
rect 23296 150554 23348 150560
rect 12992 150544 13044 150550
rect 12992 150486 13044 150492
rect 2688 150476 2740 150482
rect 2688 150418 2740 150424
rect 2700 149940 2728 150418
rect 13004 149940 13032 150486
rect 20168 150000 20220 150006
rect 16422 149938 16528 149954
rect 19826 149948 20168 149954
rect 19826 149942 20220 149948
rect 16422 149932 16540 149938
rect 16422 149926 16488 149932
rect 19826 149926 20208 149942
rect 23308 149940 23336 150554
rect 26712 149940 26740 151846
rect 33600 151836 33652 151842
rect 33600 151778 33652 151784
rect 33612 149940 33640 151778
rect 68008 151360 68060 151366
rect 68008 151302 68060 151308
rect 64512 151224 64564 151230
rect 64512 151166 64564 151172
rect 61108 151156 61160 151162
rect 61108 151098 61160 151104
rect 57704 151088 57756 151094
rect 57704 151030 57756 151036
rect 54208 151020 54260 151026
rect 54208 150962 54260 150968
rect 50804 150952 50856 150958
rect 50804 150894 50856 150900
rect 47308 150884 47360 150890
rect 47308 150826 47360 150832
rect 43904 150816 43956 150822
rect 43904 150758 43956 150764
rect 40500 150748 40552 150754
rect 40500 150690 40552 150696
rect 37004 150680 37056 150686
rect 37004 150622 37056 150628
rect 37016 149940 37044 150622
rect 40512 149940 40540 150690
rect 43916 149940 43944 150758
rect 47320 149940 47348 150826
rect 50816 149940 50844 150894
rect 54220 149940 54248 150962
rect 57716 149940 57744 151030
rect 61120 149940 61148 151098
rect 64524 149940 64552 151166
rect 68020 149940 68048 151302
rect 71700 151298 71728 151846
rect 82820 151836 82872 151842
rect 105820 151836 105872 151842
rect 82820 151778 82872 151784
rect 105740 151786 105820 151814
rect 82832 151434 82860 151778
rect 82820 151428 82872 151434
rect 82820 151370 82872 151376
rect 71688 151292 71740 151298
rect 71688 151234 71740 151240
rect 102600 150068 102652 150074
rect 102600 150010 102652 150016
rect 102612 149954 102640 150010
rect 102350 149926 102640 149954
rect 105740 149954 105768 151786
rect 105820 151778 105872 151784
rect 110328 151836 110380 151842
rect 110328 151778 110380 151784
rect 105740 149926 105846 149954
rect 16488 149874 16540 149880
rect 9588 149864 9640 149870
rect 6118 149802 6408 149818
rect 9522 149812 9588 149818
rect 9522 149806 9640 149812
rect 6118 149796 6420 149802
rect 6118 149790 6368 149796
rect 9522 149790 9628 149806
rect 6368 149738 6420 149744
rect 85488 149728 85540 149734
rect 81742 149666 82032 149682
rect 85238 149676 85488 149682
rect 85238 149670 85540 149676
rect 81742 149660 82044 149666
rect 81742 149654 81992 149660
rect 85238 149654 85528 149670
rect 81992 149602 82044 149608
rect 78588 149592 78640 149598
rect 74842 149530 75224 149546
rect 78338 149540 78588 149546
rect 78338 149534 78640 149540
rect 74842 149524 75236 149530
rect 74842 149518 75184 149524
rect 78338 149518 78628 149534
rect 75184 149466 75236 149472
rect 71688 149456 71740 149462
rect 30222 149394 30328 149410
rect 71438 149404 71688 149410
rect 71438 149398 71740 149404
rect 30222 149388 30340 149394
rect 30222 149382 30288 149388
rect 71438 149382 71728 149398
rect 88642 149382 89024 149410
rect 95542 149382 95832 149410
rect 98946 149382 99328 149410
rect 109250 149382 109632 149410
rect 30288 149330 30340 149336
rect 88996 149326 89024 149382
rect 95804 149326 95832 149382
rect 99300 149326 99328 149382
rect 88984 149320 89036 149326
rect 88984 149262 89036 149268
rect 95792 149320 95844 149326
rect 95792 149262 95844 149268
rect 99288 149320 99340 149326
rect 99288 149262 99340 149268
rect 92032 149258 92060 149260
rect 92020 149252 92072 149258
rect 92020 149194 92072 149200
rect 109604 149054 109632 149382
rect 109592 149048 109644 149054
rect 109592 148990 109644 148996
rect 110340 147626 110368 151778
rect 117228 151428 117280 151434
rect 117228 151370 117280 151376
rect 112720 151360 112772 151366
rect 112720 151302 112772 151308
rect 112628 151224 112680 151230
rect 112628 151166 112680 151172
rect 112536 151156 112588 151162
rect 112536 151098 112588 151104
rect 111708 151088 111760 151094
rect 111708 151030 111760 151036
rect 111616 150952 111668 150958
rect 111616 150894 111668 150900
rect 111524 150884 111576 150890
rect 111524 150826 111576 150832
rect 111432 150816 111484 150822
rect 111432 150758 111484 150764
rect 111340 150748 111392 150754
rect 111340 150690 111392 150696
rect 111248 150680 111300 150686
rect 111248 150622 111300 150628
rect 111064 150476 111116 150482
rect 111064 150418 111116 150424
rect 110328 147620 110380 147626
rect 110328 147562 110380 147568
rect 111076 89690 111104 150418
rect 111156 149796 111208 149802
rect 111156 149738 111208 149744
rect 111168 92478 111196 149738
rect 111260 109002 111288 150622
rect 111352 111790 111380 150690
rect 111444 113150 111472 150758
rect 111536 114510 111564 150826
rect 111628 117298 111656 150894
rect 111720 121446 111748 151030
rect 112444 151020 112496 151026
rect 112444 150962 112496 150968
rect 112352 149728 112404 149734
rect 112352 149670 112404 149676
rect 112260 149116 112312 149122
rect 112260 149058 112312 149064
rect 112272 140758 112300 149058
rect 112260 140752 112312 140758
rect 112260 140694 112312 140700
rect 112364 136610 112392 149670
rect 112352 136604 112404 136610
rect 112352 136546 112404 136552
rect 111708 121440 111760 121446
rect 111708 121382 111760 121388
rect 112456 118658 112484 150962
rect 112548 122806 112576 151098
rect 112640 124166 112668 151166
rect 112732 126954 112760 151302
rect 117044 151292 117096 151298
rect 117044 151234 117096 151240
rect 116952 150612 117004 150618
rect 116952 150554 117004 150560
rect 116676 150544 116728 150550
rect 116676 150486 116728 150492
rect 116216 150068 116268 150074
rect 116216 150010 116268 150016
rect 113088 149660 113140 149666
rect 113088 149602 113140 149608
rect 112996 149592 113048 149598
rect 112996 149534 113048 149540
rect 112904 149524 112956 149530
rect 112904 149466 112956 149472
rect 112812 149456 112864 149462
rect 112812 149398 112864 149404
rect 112824 128314 112852 149398
rect 112916 131102 112944 149466
rect 113008 132462 113036 149534
rect 113100 133890 113128 149602
rect 116032 149320 116084 149326
rect 116032 149262 116084 149268
rect 113822 144256 113878 144265
rect 113822 144191 113878 144200
rect 113088 133884 113140 133890
rect 113088 133826 113140 133832
rect 112996 132456 113048 132462
rect 112996 132398 113048 132404
rect 112904 131096 112956 131102
rect 112904 131038 112956 131044
rect 112812 128308 112864 128314
rect 112812 128250 112864 128256
rect 112720 126948 112772 126954
rect 112720 126890 112772 126896
rect 112628 124160 112680 124166
rect 112628 124102 112680 124108
rect 112536 122800 112588 122806
rect 112536 122742 112588 122748
rect 112444 118652 112496 118658
rect 112444 118594 112496 118600
rect 111616 117292 111668 117298
rect 111616 117234 111668 117240
rect 111524 114504 111576 114510
rect 111524 114446 111576 114452
rect 111432 113144 111484 113150
rect 111432 113086 111484 113092
rect 111340 111784 111392 111790
rect 111340 111726 111392 111732
rect 111248 108996 111300 109002
rect 111248 108938 111300 108944
rect 111156 92472 111208 92478
rect 111156 92414 111208 92420
rect 111064 89684 111116 89690
rect 111064 89626 111116 89632
rect 113836 88330 113864 144191
rect 116044 143313 116072 149262
rect 116124 149048 116176 149054
rect 116122 149016 116124 149025
rect 116176 149016 116178 149025
rect 116122 148951 116178 148960
rect 116124 147620 116176 147626
rect 116124 147562 116176 147568
rect 116136 147121 116164 147562
rect 116122 147112 116178 147121
rect 116122 147047 116178 147056
rect 116228 145217 116256 150010
rect 116584 149864 116636 149870
rect 116584 149806 116636 149812
rect 116400 149252 116452 149258
rect 116400 149194 116452 149200
rect 116214 145208 116270 145217
rect 116214 145143 116270 145152
rect 116030 143304 116086 143313
rect 116030 143239 116086 143248
rect 116412 141409 116440 149194
rect 116492 149184 116544 149190
rect 116492 149126 116544 149132
rect 116398 141400 116454 141409
rect 116398 141335 116454 141344
rect 116124 140752 116176 140758
rect 116124 140694 116176 140700
rect 116136 139505 116164 140694
rect 116122 139496 116178 139505
rect 116122 139431 116178 139440
rect 116504 137601 116532 149126
rect 116490 137592 116546 137601
rect 116490 137527 116546 137536
rect 116124 136604 116176 136610
rect 116124 136546 116176 136552
rect 116136 135561 116164 136546
rect 116122 135552 116178 135561
rect 116122 135487 116178 135496
rect 116032 133884 116084 133890
rect 116032 133826 116084 133832
rect 116044 133657 116072 133826
rect 116030 133648 116086 133657
rect 116030 133583 116086 133592
rect 114190 132832 114246 132841
rect 114190 132767 114246 132776
rect 114204 132666 114232 132767
rect 114192 132660 114244 132666
rect 114192 132602 114244 132608
rect 115204 132660 115256 132666
rect 115204 132602 115256 132608
rect 113914 121408 113970 121417
rect 113914 121343 113970 121352
rect 113824 88324 113876 88330
rect 113824 88266 113876 88272
rect 113928 83978 113956 121343
rect 114006 110120 114062 110129
rect 114006 110055 114062 110064
rect 113916 83972 113968 83978
rect 113916 83914 113968 83920
rect 114020 82822 114048 110055
rect 114098 98696 114154 98705
rect 114098 98631 114154 98640
rect 114008 82816 114060 82822
rect 114008 82758 114060 82764
rect 114112 80034 114140 98631
rect 114466 87272 114522 87281
rect 114466 87207 114468 87216
rect 114520 87207 114522 87216
rect 114468 87178 114520 87184
rect 115216 85649 115244 132602
rect 116124 132456 116176 132462
rect 116124 132398 116176 132404
rect 116136 131753 116164 132398
rect 116122 131744 116178 131753
rect 116122 131679 116178 131688
rect 116124 131096 116176 131102
rect 116124 131038 116176 131044
rect 116136 129849 116164 131038
rect 116122 129840 116178 129849
rect 116122 129775 116178 129784
rect 116124 128308 116176 128314
rect 116124 128250 116176 128256
rect 116136 127945 116164 128250
rect 116122 127936 116178 127945
rect 116122 127871 116178 127880
rect 116032 126948 116084 126954
rect 116032 126890 116084 126896
rect 116044 126041 116072 126890
rect 116030 126032 116086 126041
rect 116030 125967 116086 125976
rect 116124 124160 116176 124166
rect 116122 124128 116124 124137
rect 116176 124128 116178 124137
rect 116122 124063 116178 124072
rect 115940 122800 115992 122806
rect 115940 122742 115992 122748
rect 115952 122233 115980 122742
rect 115938 122224 115994 122233
rect 115938 122159 115994 122168
rect 116124 121440 116176 121446
rect 116124 121382 116176 121388
rect 116136 120193 116164 121382
rect 116122 120184 116178 120193
rect 116122 120119 116178 120128
rect 116124 118652 116176 118658
rect 116124 118594 116176 118600
rect 116136 118289 116164 118594
rect 116122 118280 116178 118289
rect 116122 118215 116178 118224
rect 116492 118040 116544 118046
rect 116492 117982 116544 117988
rect 116124 117292 116176 117298
rect 116124 117234 116176 117240
rect 116136 116385 116164 117234
rect 116122 116376 116178 116385
rect 116122 116311 116178 116320
rect 116124 114504 116176 114510
rect 116122 114472 116124 114481
rect 116176 114472 116178 114481
rect 116122 114407 116178 114416
rect 115940 113144 115992 113150
rect 115940 113086 115992 113092
rect 115952 112577 115980 113086
rect 115938 112568 115994 112577
rect 115938 112503 115994 112512
rect 116124 111784 116176 111790
rect 116124 111726 116176 111732
rect 116136 110673 116164 111726
rect 116122 110664 116178 110673
rect 116122 110599 116178 110608
rect 116124 108996 116176 109002
rect 116124 108938 116176 108944
rect 116136 108769 116164 108938
rect 116122 108760 116178 108769
rect 116122 108695 116178 108704
rect 116504 106865 116532 117982
rect 116490 106856 116546 106865
rect 116490 106791 116546 106800
rect 116596 93401 116624 149806
rect 116688 95305 116716 150486
rect 116860 150000 116912 150006
rect 116860 149942 116912 149948
rect 116768 149932 116820 149938
rect 116768 149874 116820 149880
rect 116780 97209 116808 149874
rect 116872 99113 116900 149942
rect 116964 101017 116992 150554
rect 117056 102921 117084 151234
rect 117136 149388 117188 149394
rect 117136 149330 117188 149336
rect 117148 104825 117176 149330
rect 117240 118046 117268 151370
rect 118896 149954 118924 157966
rect 119988 154624 120040 154630
rect 119988 154566 120040 154572
rect 120000 154426 120028 154566
rect 119896 154420 119948 154426
rect 119896 154362 119948 154368
rect 119988 154420 120040 154426
rect 119988 154362 120040 154368
rect 119908 153882 119936 154362
rect 119804 153876 119856 153882
rect 119804 153818 119856 153824
rect 119896 153876 119948 153882
rect 119896 153818 119948 153824
rect 119816 150192 119844 153818
rect 120092 152386 120120 163254
rect 120552 163146 120580 163254
rect 120630 163200 120686 164400
rect 121458 163200 121514 164400
rect 122286 163200 122342 164400
rect 123114 163200 123170 164400
rect 124034 163200 124090 164400
rect 124862 163200 124918 164400
rect 125690 163200 125746 164400
rect 126518 163200 126574 164400
rect 126992 163254 127296 163282
rect 120644 163146 120672 163200
rect 120552 163118 120672 163146
rect 120448 156664 120500 156670
rect 120448 156606 120500 156612
rect 120080 152380 120132 152386
rect 120080 152322 120132 152328
rect 120460 150192 120488 156606
rect 121472 156058 121500 163200
rect 121920 158976 121972 158982
rect 121920 158918 121972 158924
rect 121460 156052 121512 156058
rect 121460 155994 121512 156000
rect 121932 153785 121960 158918
rect 122012 155304 122064 155310
rect 122012 155246 122064 155252
rect 121734 153776 121790 153785
rect 121734 153711 121790 153720
rect 121918 153776 121974 153785
rect 121918 153711 121974 153720
rect 121092 152516 121144 152522
rect 121092 152458 121144 152464
rect 121104 150192 121132 152458
rect 121748 150192 121776 153711
rect 122024 151814 122052 155246
rect 122300 154970 122328 163200
rect 123128 159390 123156 163200
rect 122840 159384 122892 159390
rect 122840 159326 122892 159332
rect 123116 159384 123168 159390
rect 123116 159326 123168 159332
rect 122288 154964 122340 154970
rect 122288 154906 122340 154912
rect 122024 151786 122420 151814
rect 122392 150226 122420 151786
rect 122392 150198 122466 150226
rect 122852 150210 122880 159326
rect 124048 158982 124076 163200
rect 124036 158976 124088 158982
rect 124036 158918 124088 158924
rect 124876 156670 124904 163200
rect 125704 161474 125732 163200
rect 125704 161446 125824 161474
rect 125508 158908 125560 158914
rect 125508 158850 125560 158856
rect 124864 156664 124916 156670
rect 124864 156606 124916 156612
rect 124680 155372 124732 155378
rect 124680 155314 124732 155320
rect 123024 155236 123076 155242
rect 123024 155178 123076 155184
rect 123036 150226 123064 155178
rect 124312 153944 124364 153950
rect 124312 153886 124364 153892
rect 124324 150226 124352 153886
rect 124692 151814 124720 155314
rect 125520 153950 125548 158850
rect 125692 155440 125744 155446
rect 125692 155382 125744 155388
rect 125508 153944 125560 153950
rect 125508 153886 125560 153892
rect 124692 151786 124996 151814
rect 124968 150226 124996 151786
rect 125704 150226 125732 155382
rect 125796 155310 125824 161446
rect 126532 159730 126560 163200
rect 126428 159724 126480 159730
rect 126428 159666 126480 159672
rect 126520 159724 126572 159730
rect 126520 159666 126572 159672
rect 126440 159526 126468 159666
rect 126336 159520 126388 159526
rect 126336 159462 126388 159468
rect 126428 159520 126480 159526
rect 126428 159462 126480 159468
rect 126348 158914 126376 159462
rect 126612 159452 126664 159458
rect 126612 159394 126664 159400
rect 126336 158908 126388 158914
rect 126336 158850 126388 158856
rect 125784 155304 125836 155310
rect 125784 155246 125836 155252
rect 126624 152425 126652 159394
rect 126888 154012 126940 154018
rect 126888 153954 126940 153960
rect 126242 152416 126298 152425
rect 126242 152351 126298 152360
rect 126610 152416 126666 152425
rect 126610 152351 126666 152360
rect 119816 150164 119890 150192
rect 120460 150164 120534 150192
rect 121104 150164 121178 150192
rect 121748 150164 121822 150192
rect 118896 149926 119324 149954
rect 119862 149940 119890 150164
rect 120506 149940 120534 150164
rect 121150 149940 121178 150164
rect 121794 149940 121822 150164
rect 122438 149940 122466 150198
rect 122840 150204 122892 150210
rect 123036 150198 123110 150226
rect 122840 150146 122892 150152
rect 123082 149940 123110 150198
rect 123714 150204 123766 150210
rect 124324 150198 124398 150226
rect 124968 150198 125042 150226
rect 123714 150146 123766 150152
rect 123726 149940 123754 150146
rect 124370 149940 124398 150198
rect 125014 149940 125042 150198
rect 125658 150198 125732 150226
rect 126256 150226 126284 152351
rect 126900 150226 126928 153954
rect 126992 152522 127020 163254
rect 127268 163146 127296 163254
rect 127346 163200 127402 164400
rect 128174 163200 128230 164400
rect 129002 163200 129058 164400
rect 129922 163200 129978 164400
rect 130750 163200 130806 164400
rect 131578 163200 131634 164400
rect 132406 163200 132462 164400
rect 133234 163200 133290 164400
rect 134062 163200 134118 164400
rect 134890 163200 134946 164400
rect 135810 163200 135866 164400
rect 136638 163200 136694 164400
rect 136744 163254 137416 163282
rect 127360 163146 127388 163200
rect 127268 163118 127388 163146
rect 127624 159520 127676 159526
rect 127624 159462 127676 159468
rect 127532 156732 127584 156738
rect 127532 156674 127584 156680
rect 126980 152516 127032 152522
rect 126980 152458 127032 152464
rect 127544 150226 127572 156674
rect 127636 154018 127664 159462
rect 128188 156738 128216 163200
rect 128176 156732 128228 156738
rect 128176 156674 128228 156680
rect 129016 155242 129044 163200
rect 129936 159526 129964 163200
rect 129924 159520 129976 159526
rect 129924 159462 129976 159468
rect 130764 159458 130792 163200
rect 130752 159452 130804 159458
rect 130752 159394 130804 159400
rect 131026 159352 131082 159361
rect 131026 159287 131082 159296
rect 129740 158908 129792 158914
rect 129740 158850 129792 158856
rect 129004 155236 129056 155242
rect 129004 155178 129056 155184
rect 129384 154142 129688 154170
rect 129280 154080 129332 154086
rect 129280 154022 129332 154028
rect 127624 154012 127676 154018
rect 127624 153954 127676 153960
rect 128818 152552 128874 152561
rect 128818 152487 128874 152496
rect 128176 151836 128228 151842
rect 128176 151778 128228 151784
rect 128188 150226 128216 151778
rect 128832 150226 128860 152487
rect 129292 151814 129320 154022
rect 129384 154018 129412 154142
rect 129660 154018 129688 154142
rect 129372 154012 129424 154018
rect 129372 153954 129424 153960
rect 129648 154012 129700 154018
rect 129648 153954 129700 153960
rect 129752 151842 129780 158850
rect 130108 156800 130160 156806
rect 130108 156742 130160 156748
rect 129740 151836 129792 151842
rect 129292 151786 129504 151814
rect 129476 150226 129504 151786
rect 129740 151778 129792 151784
rect 130120 150226 130148 156742
rect 130752 152244 130804 152250
rect 130752 152186 130804 152192
rect 130764 150226 130792 152186
rect 131040 151814 131068 159287
rect 131592 158030 131620 163200
rect 131580 158024 131632 158030
rect 131580 157966 131632 157972
rect 132420 153950 132448 163200
rect 133248 158846 133276 163200
rect 133602 159488 133658 159497
rect 133602 159423 133658 159432
rect 133236 158840 133288 158846
rect 133236 158782 133288 158788
rect 132500 156868 132552 156874
rect 132500 156810 132552 156816
rect 132408 153944 132460 153950
rect 132038 153912 132094 153921
rect 132408 153886 132460 153892
rect 132038 153847 132094 153856
rect 131040 151786 131436 151814
rect 131408 150226 131436 151786
rect 132052 150226 132080 153847
rect 132512 151814 132540 156810
rect 133052 154760 133104 154766
rect 133052 154702 133104 154708
rect 133064 151814 133092 154702
rect 133616 153105 133644 159423
rect 133602 153096 133658 153105
rect 133602 153031 133658 153040
rect 133972 152584 134024 152590
rect 133972 152526 134024 152532
rect 132512 151786 132724 151814
rect 133064 151786 133368 151814
rect 132696 150226 132724 151786
rect 133340 150226 133368 151786
rect 133984 150226 134012 152526
rect 134076 152250 134104 163200
rect 134904 156874 134932 163200
rect 135824 156942 135852 163200
rect 136652 163146 136680 163200
rect 136744 163146 136772 163254
rect 136652 163118 136772 163146
rect 137388 159798 137416 163254
rect 137466 163200 137522 164400
rect 138294 163200 138350 164400
rect 139122 163200 139178 164400
rect 139950 163200 140006 164400
rect 140778 163200 140834 164400
rect 141698 163200 141754 164400
rect 142526 163200 142582 164400
rect 143354 163200 143410 164400
rect 144182 163200 144238 164400
rect 145010 163200 145066 164400
rect 145838 163200 145894 164400
rect 146666 163200 146722 164400
rect 147586 163200 147642 164400
rect 148414 163200 148470 164400
rect 149242 163200 149298 164400
rect 150070 163200 150126 164400
rect 150898 163200 150954 164400
rect 151726 163200 151782 164400
rect 151924 163254 152504 163282
rect 137284 159792 137336 159798
rect 137284 159734 137336 159740
rect 137376 159792 137428 159798
rect 137376 159734 137428 159740
rect 137296 159594 137324 159734
rect 136824 159588 136876 159594
rect 136824 159530 136876 159536
rect 137284 159588 137336 159594
rect 137284 159530 137336 159536
rect 135260 156936 135312 156942
rect 135260 156878 135312 156884
rect 135812 156936 135864 156942
rect 135812 156878 135864 156884
rect 134892 156868 134944 156874
rect 134892 156810 134944 156816
rect 134614 154048 134670 154057
rect 134614 153983 134670 153992
rect 134064 152244 134116 152250
rect 134064 152186 134116 152192
rect 134628 150226 134656 153983
rect 135272 150226 135300 156878
rect 136546 153096 136602 153105
rect 136546 153031 136602 153040
rect 135904 152652 135956 152658
rect 135904 152594 135956 152600
rect 135916 150226 135944 152594
rect 136560 150226 136588 153031
rect 136836 152590 136864 159530
rect 137192 159452 137244 159458
rect 137192 159394 137244 159400
rect 137204 158914 137232 159394
rect 137480 159390 137508 163200
rect 138018 159624 138074 159633
rect 138018 159559 138074 159568
rect 137468 159384 137520 159390
rect 137468 159326 137520 159332
rect 137100 158908 137152 158914
rect 137100 158850 137152 158856
rect 137192 158908 137244 158914
rect 137192 158850 137244 158856
rect 137112 154630 137140 158850
rect 138032 157334 138060 159559
rect 138032 157306 138152 157334
rect 137376 157004 137428 157010
rect 137376 156946 137428 156952
rect 137100 154624 137152 154630
rect 137100 154566 137152 154572
rect 136928 154278 137140 154306
rect 136928 154222 136956 154278
rect 136916 154216 136968 154222
rect 136916 154158 136968 154164
rect 137112 154170 137140 154278
rect 137008 154148 137060 154154
rect 137112 154142 137324 154170
rect 137008 154090 137060 154096
rect 136824 152584 136876 152590
rect 136824 152526 136876 152532
rect 137020 151814 137048 154090
rect 137296 154086 137324 154142
rect 137284 154080 137336 154086
rect 137284 154022 137336 154028
rect 137388 151814 137416 156946
rect 138020 154624 138072 154630
rect 138020 154566 138072 154572
rect 138032 153950 138060 154566
rect 138020 153944 138072 153950
rect 138020 153886 138072 153892
rect 138124 152862 138152 157306
rect 138308 157010 138336 163200
rect 138296 157004 138348 157010
rect 138296 156946 138348 156952
rect 139136 156806 139164 163200
rect 139964 159798 139992 163200
rect 139400 159792 139452 159798
rect 139400 159734 139452 159740
rect 139952 159792 140004 159798
rect 139952 159734 140004 159740
rect 139412 157334 139440 159734
rect 139412 157306 139900 157334
rect 139124 156800 139176 156806
rect 139124 156742 139176 156748
rect 139308 154828 139360 154834
rect 139308 154770 139360 154776
rect 138386 153640 138442 153649
rect 138386 153575 138442 153584
rect 138400 153270 138428 153575
rect 138388 153264 138440 153270
rect 138388 153206 138440 153212
rect 138020 152856 138072 152862
rect 138020 152798 138072 152804
rect 138112 152856 138164 152862
rect 138112 152798 138164 152804
rect 138032 152674 138060 152798
rect 139124 152788 139176 152794
rect 139124 152730 139176 152736
rect 138032 152646 138152 152674
rect 138124 152590 138152 152646
rect 138112 152584 138164 152590
rect 138112 152526 138164 152532
rect 138480 151904 138532 151910
rect 138480 151846 138532 151852
rect 137020 151786 137232 151814
rect 137388 151786 137876 151814
rect 137204 150226 137232 151786
rect 137848 150226 137876 151786
rect 126256 150198 126330 150226
rect 126900 150198 126974 150226
rect 127544 150198 127618 150226
rect 128188 150198 128262 150226
rect 128832 150198 128906 150226
rect 129476 150198 129550 150226
rect 130120 150198 130194 150226
rect 130764 150198 130838 150226
rect 131408 150198 131482 150226
rect 132052 150198 132126 150226
rect 132696 150198 132770 150226
rect 133340 150198 133414 150226
rect 133984 150198 134058 150226
rect 134628 150198 134702 150226
rect 135272 150198 135346 150226
rect 135916 150198 135990 150226
rect 136560 150198 136634 150226
rect 137204 150198 137278 150226
rect 137848 150198 137922 150226
rect 125658 149940 125686 150198
rect 126302 149940 126330 150198
rect 126946 149940 126974 150198
rect 127590 149940 127618 150198
rect 128234 149940 128262 150198
rect 128878 149940 128906 150198
rect 129522 149940 129550 150198
rect 130166 149940 130194 150198
rect 130810 149940 130838 150198
rect 131454 149940 131482 150198
rect 132098 149940 132126 150198
rect 132742 149940 132770 150198
rect 133386 149940 133414 150198
rect 134030 149940 134058 150198
rect 134674 149940 134702 150198
rect 135318 149940 135346 150198
rect 135962 149940 135990 150198
rect 136606 149940 136634 150198
rect 137250 149940 137278 150198
rect 137894 149940 137922 150198
rect 138492 150090 138520 151846
rect 139136 150090 139164 152730
rect 139320 151910 139348 154770
rect 139872 154086 139900 157306
rect 140410 156768 140466 156777
rect 140410 156703 140466 156712
rect 139768 154080 139820 154086
rect 139768 154022 139820 154028
rect 139860 154080 139912 154086
rect 139860 154022 139912 154028
rect 139308 151904 139360 151910
rect 139308 151846 139360 151852
rect 139780 150090 139808 154022
rect 140424 150090 140452 156703
rect 140792 152794 140820 163200
rect 141712 157418 141740 163200
rect 141700 157412 141752 157418
rect 141700 157354 141752 157360
rect 142540 155378 142568 163200
rect 143368 159662 143396 163200
rect 143264 159656 143316 159662
rect 143264 159598 143316 159604
rect 143356 159656 143408 159662
rect 143356 159598 143408 159604
rect 143276 157334 143304 159598
rect 144000 159588 144052 159594
rect 144000 159530 144052 159536
rect 144092 159588 144144 159594
rect 144092 159530 144144 159536
rect 144012 159338 144040 159530
rect 144104 159458 144132 159530
rect 144196 159458 144224 163200
rect 144092 159452 144144 159458
rect 144092 159394 144144 159400
rect 144184 159452 144236 159458
rect 144184 159394 144236 159400
rect 144012 159310 144408 159338
rect 143276 157306 143488 157334
rect 143170 156632 143226 156641
rect 143170 156567 143226 156576
rect 142528 155372 142580 155378
rect 142528 155314 142580 155320
rect 142896 154488 142948 154494
rect 142448 154414 142752 154442
rect 142896 154430 142948 154436
rect 142988 154488 143040 154494
rect 142988 154430 143040 154436
rect 142342 154184 142398 154193
rect 142448 154154 142476 154414
rect 142724 154358 142752 154414
rect 142620 154352 142672 154358
rect 142620 154294 142672 154300
rect 142712 154352 142764 154358
rect 142712 154294 142764 154300
rect 142342 154119 142398 154128
rect 142436 154148 142488 154154
rect 141700 152856 141752 152862
rect 141700 152798 141752 152804
rect 140780 152788 140832 152794
rect 140780 152730 140832 152736
rect 141056 152720 141108 152726
rect 141056 152662 141108 152668
rect 141068 150090 141096 152662
rect 141712 150090 141740 152798
rect 142356 150090 142384 154119
rect 142436 154090 142488 154096
rect 142528 154080 142580 154086
rect 142632 154057 142660 154294
rect 142908 154222 142936 154430
rect 142896 154216 142948 154222
rect 142896 154158 142948 154164
rect 143000 154086 143028 154430
rect 143080 154284 143132 154290
rect 143080 154226 143132 154232
rect 142988 154080 143040 154086
rect 142528 154022 142580 154028
rect 142618 154048 142674 154057
rect 142540 153921 142568 154022
rect 142988 154022 143040 154028
rect 142618 153983 142674 153992
rect 143092 153950 143120 154226
rect 143080 153944 143132 153950
rect 142526 153912 142582 153921
rect 143080 153886 143132 153892
rect 142526 153847 142582 153856
rect 142804 153876 142856 153882
rect 142804 153818 142856 153824
rect 142816 153270 142844 153818
rect 142804 153264 142856 153270
rect 142804 153206 142856 153212
rect 142804 152720 142856 152726
rect 142804 152662 142856 152668
rect 142816 152046 142844 152662
rect 142804 152040 142856 152046
rect 142804 151982 142856 151988
rect 143184 150226 143212 156567
rect 143262 154048 143318 154057
rect 143262 153983 143318 153992
rect 143276 153950 143304 153983
rect 143264 153944 143316 153950
rect 143264 153886 143316 153892
rect 143354 153912 143410 153921
rect 143354 153847 143356 153856
rect 143408 153847 143410 153856
rect 143356 153818 143408 153824
rect 143460 152046 143488 157306
rect 143540 154080 143592 154086
rect 143540 154022 143592 154028
rect 143552 153649 143580 154022
rect 143538 153640 143594 153649
rect 143538 153575 143594 153584
rect 144380 152794 144408 159310
rect 145024 155990 145052 163200
rect 145102 157992 145158 158001
rect 145102 157927 145158 157936
rect 145012 155984 145064 155990
rect 145012 155926 145064 155932
rect 144276 152788 144328 152794
rect 144276 152730 144328 152736
rect 144368 152788 144420 152794
rect 144368 152730 144420 152736
rect 144288 152674 144316 152730
rect 144288 152646 144408 152674
rect 144380 152590 144408 152646
rect 144276 152584 144328 152590
rect 144276 152526 144328 152532
rect 144368 152584 144420 152590
rect 144368 152526 144420 152532
rect 143630 152416 143686 152425
rect 143630 152351 143686 152360
rect 143448 152040 143500 152046
rect 143448 151982 143500 151988
rect 143046 150198 143212 150226
rect 138492 150062 138566 150090
rect 139136 150062 139210 150090
rect 139780 150062 139854 150090
rect 140424 150062 140498 150090
rect 141068 150062 141142 150090
rect 141712 150062 141786 150090
rect 142356 150062 142430 150090
rect 138538 149940 138566 150062
rect 139182 149940 139210 150062
rect 139826 149940 139854 150062
rect 140470 149940 140498 150062
rect 141114 149940 141142 150062
rect 141758 149940 141786 150062
rect 142402 149940 142430 150062
rect 143046 149940 143074 150198
rect 143644 150090 143672 152351
rect 144288 150090 144316 152526
rect 145116 150226 145144 157927
rect 145852 155446 145880 163200
rect 146484 160064 146536 160070
rect 146484 160006 146536 160012
rect 146392 158092 146444 158098
rect 146392 158034 146444 158040
rect 146208 157072 146260 157078
rect 146208 157014 146260 157020
rect 145840 155440 145892 155446
rect 145840 155382 145892 155388
rect 145564 153944 145616 153950
rect 145564 153886 145616 153892
rect 144978 150198 145144 150226
rect 143644 150062 143718 150090
rect 144288 150062 144362 150090
rect 143690 149940 143718 150062
rect 144334 149940 144362 150062
rect 144978 149940 145006 150198
rect 145576 150090 145604 153886
rect 146220 150090 146248 157014
rect 146404 150210 146432 158034
rect 146496 152862 146524 160006
rect 146680 158778 146708 163200
rect 146944 160064 146996 160070
rect 146944 160006 146996 160012
rect 146852 159588 146904 159594
rect 146852 159530 146904 159536
rect 146864 159338 146892 159530
rect 146956 159526 146984 160006
rect 147048 159854 147260 159882
rect 147048 159798 147076 159854
rect 147036 159792 147088 159798
rect 147036 159734 147088 159740
rect 147128 159792 147180 159798
rect 147128 159734 147180 159740
rect 146944 159520 146996 159526
rect 147140 159474 147168 159734
rect 147232 159594 147260 159854
rect 147220 159588 147272 159594
rect 147220 159530 147272 159536
rect 146944 159462 146996 159468
rect 147048 159446 147168 159474
rect 147600 159458 147628 163200
rect 148324 159792 148376 159798
rect 148324 159734 148376 159740
rect 147588 159452 147640 159458
rect 147048 159338 147076 159446
rect 147588 159394 147640 159400
rect 146864 159310 147076 159338
rect 146576 158772 146628 158778
rect 146576 158714 146628 158720
rect 146668 158772 146720 158778
rect 146668 158714 146720 158720
rect 146588 158658 146616 158714
rect 146588 158630 147444 158658
rect 147416 153882 147444 158630
rect 148336 154154 148364 159734
rect 148428 158098 148456 163200
rect 148416 158092 148468 158098
rect 148416 158034 148468 158040
rect 148784 157140 148836 157146
rect 148784 157082 148836 157088
rect 148140 154148 148192 154154
rect 148140 154090 148192 154096
rect 148324 154148 148376 154154
rect 148324 154090 148376 154096
rect 147404 153876 147456 153882
rect 147404 153818 147456 153824
rect 146484 152856 146536 152862
rect 146484 152798 146536 152804
rect 146944 152040 146996 152046
rect 146944 151982 146996 151988
rect 146956 151842 146984 151982
rect 146852 151836 146904 151842
rect 146852 151778 146904 151784
rect 146944 151836 146996 151842
rect 146944 151778 146996 151784
rect 146392 150204 146444 150210
rect 146392 150146 146444 150152
rect 146864 150090 146892 151778
rect 147542 150204 147594 150210
rect 147542 150146 147594 150152
rect 145576 150062 145650 150090
rect 146220 150062 146294 150090
rect 146864 150062 146938 150090
rect 145622 149940 145650 150062
rect 146266 149940 146294 150062
rect 146910 149940 146938 150062
rect 147554 149940 147582 150146
rect 148152 150090 148180 154090
rect 148796 150090 148824 157082
rect 149256 154834 149284 163200
rect 149520 159452 149572 159458
rect 149520 159394 149572 159400
rect 149244 154828 149296 154834
rect 149244 154770 149296 154776
rect 149532 152726 149560 159394
rect 149610 158264 149666 158273
rect 149610 158199 149666 158208
rect 149624 157334 149652 158199
rect 149624 157306 150020 157334
rect 149428 152720 149480 152726
rect 149428 152662 149480 152668
rect 149520 152720 149572 152726
rect 149520 152662 149572 152668
rect 149440 150090 149468 152662
rect 149992 150226 150020 157306
rect 150084 157146 150112 163200
rect 150912 159458 150940 163200
rect 150900 159452 150952 159458
rect 150900 159394 150952 159400
rect 151268 157208 151320 157214
rect 151268 157150 151320 157156
rect 150072 157140 150124 157146
rect 150072 157082 150124 157088
rect 150624 154080 150676 154086
rect 150624 154022 150676 154028
rect 149992 150198 150066 150226
rect 148152 150062 148226 150090
rect 148796 150062 148870 150090
rect 149440 150062 149514 150090
rect 148198 149940 148226 150062
rect 148842 149940 148870 150062
rect 149486 149940 149514 150062
rect 150038 149940 150066 150198
rect 150636 150090 150664 154022
rect 151280 150226 151308 157150
rect 151740 157078 151768 163200
rect 151728 157072 151780 157078
rect 151728 157014 151780 157020
rect 151924 154766 151952 163254
rect 152476 163146 152504 163254
rect 152554 163200 152610 164400
rect 153474 163200 153530 164400
rect 153580 163254 154252 163282
rect 152568 163146 152596 163200
rect 152476 163118 152596 163146
rect 153488 159798 153516 163200
rect 153476 159792 153528 159798
rect 153476 159734 153528 159740
rect 152554 158128 152610 158137
rect 152554 158063 152610 158072
rect 151912 154760 151964 154766
rect 151912 154702 151964 154708
rect 152464 154556 152516 154562
rect 152464 154498 152516 154504
rect 152476 154290 152504 154498
rect 152464 154284 152516 154290
rect 152464 154226 152516 154232
rect 152280 154216 152332 154222
rect 152280 154158 152332 154164
rect 152188 154080 152240 154086
rect 152188 154022 152240 154028
rect 152200 153921 152228 154022
rect 152186 153912 152242 153921
rect 152186 153847 152242 153856
rect 152292 153678 152320 154158
rect 152372 154080 152424 154086
rect 152372 154022 152424 154028
rect 152384 153882 152412 154022
rect 152372 153876 152424 153882
rect 152372 153818 152424 153824
rect 152280 153672 152332 153678
rect 152280 153614 152332 153620
rect 151912 152652 151964 152658
rect 151912 152594 151964 152600
rect 151280 150198 151354 150226
rect 150636 150062 150710 150090
rect 150682 149940 150710 150062
rect 151326 149940 151354 150198
rect 151924 150090 151952 152594
rect 152568 150226 152596 158063
rect 153108 154760 153160 154766
rect 153108 154702 153160 154708
rect 152648 154624 152700 154630
rect 152648 154566 152700 154572
rect 152660 154290 152688 154566
rect 153120 154306 153148 154702
rect 152648 154284 152700 154290
rect 153120 154278 153332 154306
rect 152648 154226 152700 154232
rect 153304 154154 153332 154278
rect 153200 154148 153252 154154
rect 153200 154090 153252 154096
rect 153292 154148 153344 154154
rect 153292 154090 153344 154096
rect 152646 153912 152702 153921
rect 152646 153847 152702 153856
rect 152660 153814 152688 153847
rect 152648 153808 152700 153814
rect 152648 153750 152700 153756
rect 152568 150198 152642 150226
rect 151924 150062 151998 150090
rect 151970 149940 151998 150062
rect 152614 149940 152642 150198
rect 153212 150090 153240 154090
rect 153580 152658 153608 163254
rect 154224 163146 154252 163254
rect 154302 163200 154358 164400
rect 155130 163200 155186 164400
rect 155958 163200 156014 164400
rect 156786 163200 156842 164400
rect 157614 163200 157670 164400
rect 158442 163200 158498 164400
rect 159362 163200 159418 164400
rect 160190 163200 160246 164400
rect 161018 163200 161074 164400
rect 161846 163200 161902 164400
rect 162674 163200 162730 164400
rect 163502 163200 163558 164400
rect 164330 163200 164386 164400
rect 165250 163200 165306 164400
rect 165632 163254 166028 163282
rect 154316 163146 154344 163200
rect 154224 163118 154344 163146
rect 154488 160064 154540 160070
rect 154488 160006 154540 160012
rect 153844 157276 153896 157282
rect 153844 157218 153896 157224
rect 153568 152652 153620 152658
rect 153568 152594 153620 152600
rect 153856 150090 153884 157218
rect 154500 153678 154528 160006
rect 155144 158166 155172 163200
rect 155040 158160 155092 158166
rect 155040 158102 155092 158108
rect 155132 158160 155184 158166
rect 155132 158102 155184 158108
rect 155052 157334 155080 158102
rect 155052 157306 155172 157334
rect 154488 153672 154540 153678
rect 154488 153614 154540 153620
rect 154488 151972 154540 151978
rect 154488 151914 154540 151920
rect 154500 150090 154528 151914
rect 155144 150226 155172 157306
rect 155972 154766 156000 163200
rect 156800 160070 156828 163200
rect 156788 160064 156840 160070
rect 156788 160006 156840 160012
rect 156328 159860 156380 159866
rect 156328 159802 156380 159808
rect 155960 154760 156012 154766
rect 155960 154702 156012 154708
rect 155776 154284 155828 154290
rect 155776 154226 155828 154232
rect 155144 150198 155218 150226
rect 153212 150062 153286 150090
rect 153856 150062 153930 150090
rect 154500 150062 154574 150090
rect 153258 149940 153286 150062
rect 153902 149940 153930 150062
rect 154546 149940 154574 150062
rect 155190 149940 155218 150198
rect 155788 150090 155816 154226
rect 156340 152046 156368 159802
rect 156604 159792 156656 159798
rect 156788 159792 156840 159798
rect 156656 159740 156788 159746
rect 156604 159734 156840 159740
rect 156512 159724 156564 159730
rect 156616 159718 156828 159734
rect 156512 159666 156564 159672
rect 156420 157344 156472 157350
rect 156420 157286 156472 157292
rect 156328 152040 156380 152046
rect 156328 151982 156380 151988
rect 156432 150090 156460 157286
rect 156524 157214 156552 159666
rect 157628 159594 157656 163200
rect 157616 159588 157668 159594
rect 157616 159530 157668 159536
rect 158456 158234 158484 163200
rect 158720 158840 158772 158846
rect 158720 158782 158772 158788
rect 157708 158228 157760 158234
rect 157708 158170 157760 158176
rect 158444 158228 158496 158234
rect 158444 158170 158496 158176
rect 156512 157208 156564 157214
rect 156512 157150 156564 157156
rect 157064 151836 157116 151842
rect 157064 151778 157116 151784
rect 157076 150090 157104 151778
rect 157720 150226 157748 158170
rect 158732 157350 158760 158782
rect 158720 157344 158772 157350
rect 158720 157286 158772 157292
rect 159088 157208 159140 157214
rect 159088 157150 159140 157156
rect 159100 156602 159128 157150
rect 158996 156596 159048 156602
rect 158996 156538 159048 156544
rect 159088 156596 159140 156602
rect 159088 156538 159140 156544
rect 158444 154148 158496 154154
rect 158444 154090 158496 154096
rect 158456 153882 158484 154090
rect 158352 153876 158404 153882
rect 158352 153818 158404 153824
rect 158444 153876 158496 153882
rect 158444 153818 158496 153824
rect 158364 150226 158392 153818
rect 159008 150226 159036 156538
rect 159376 154698 159404 163200
rect 160100 159860 160152 159866
rect 160100 159802 160152 159808
rect 160112 157214 160140 159802
rect 160100 157208 160152 157214
rect 160100 157150 160152 157156
rect 159364 154692 159416 154698
rect 159364 154634 159416 154640
rect 160204 154154 160232 163200
rect 161032 159662 161060 163200
rect 161020 159656 161072 159662
rect 161020 159598 161072 159604
rect 161860 158302 161888 163200
rect 162492 159928 162544 159934
rect 162492 159870 162544 159876
rect 160284 158296 160336 158302
rect 160284 158238 160336 158244
rect 161848 158296 161900 158302
rect 161848 158238 161900 158244
rect 160192 154148 160244 154154
rect 160192 154090 160244 154096
rect 159640 152448 159692 152454
rect 159640 152390 159692 152396
rect 159652 150226 159680 152390
rect 160296 150226 160324 158238
rect 161662 156904 161718 156913
rect 161662 156839 161718 156848
rect 160926 154320 160982 154329
rect 160926 154255 160982 154264
rect 161480 154284 161532 154290
rect 160940 150226 160968 154255
rect 161480 154226 161532 154232
rect 161492 153746 161520 154226
rect 161572 154080 161624 154086
rect 161572 154022 161624 154028
rect 161584 153746 161612 154022
rect 161480 153740 161532 153746
rect 161480 153682 161532 153688
rect 161572 153740 161624 153746
rect 161572 153682 161624 153688
rect 161676 150226 161704 156839
rect 162216 152788 162268 152794
rect 162216 152730 162268 152736
rect 157720 150198 157794 150226
rect 158364 150198 158438 150226
rect 159008 150198 159082 150226
rect 159652 150198 159726 150226
rect 160296 150198 160370 150226
rect 160940 150198 161014 150226
rect 155788 150062 155862 150090
rect 156432 150062 156506 150090
rect 157076 150062 157150 150090
rect 155834 149940 155862 150062
rect 156478 149940 156506 150062
rect 157122 149940 157150 150062
rect 157766 149940 157794 150198
rect 158410 149940 158438 150198
rect 159054 149940 159082 150198
rect 159698 149940 159726 150198
rect 160342 149940 160370 150198
rect 160986 149940 161014 150198
rect 161630 150198 161704 150226
rect 162228 150226 162256 152730
rect 162504 151978 162532 159870
rect 162688 154630 162716 163200
rect 162872 159186 163084 159202
rect 162872 159180 163096 159186
rect 162872 159174 163044 159180
rect 162872 159118 162900 159174
rect 163044 159122 163096 159128
rect 162860 159112 162912 159118
rect 162860 159054 162912 159060
rect 163516 158846 163544 163200
rect 164344 161474 164372 163200
rect 164344 161446 164464 161474
rect 163780 159724 163832 159730
rect 163780 159666 163832 159672
rect 163504 158840 163556 158846
rect 163504 158782 163556 158788
rect 162858 158400 162914 158409
rect 162858 158335 162914 158344
rect 162676 154624 162728 154630
rect 162676 154566 162728 154572
rect 162492 151972 162544 151978
rect 162492 151914 162544 151920
rect 162872 150226 162900 158335
rect 163792 157282 163820 159666
rect 164332 158364 164384 158370
rect 164332 158306 164384 158312
rect 163780 157276 163832 157282
rect 163780 157218 163832 157224
rect 164148 156528 164200 156534
rect 164148 156470 164200 156476
rect 163504 154216 163556 154222
rect 163504 154158 163556 154164
rect 163516 150226 163544 154158
rect 164160 150226 164188 156470
rect 162228 150198 162302 150226
rect 162872 150198 162946 150226
rect 163516 150198 163590 150226
rect 164160 150198 164234 150226
rect 164344 150210 164372 158306
rect 164436 152794 164464 161446
rect 165264 158370 165292 163200
rect 165252 158364 165304 158370
rect 165252 158306 165304 158312
rect 164884 157888 164936 157894
rect 164882 157856 164884 157865
rect 164936 157856 164938 157865
rect 164882 157791 164938 157800
rect 165632 154154 165660 163254
rect 166000 163146 166028 163254
rect 166078 163200 166134 164400
rect 166906 163200 166962 164400
rect 167734 163200 167790 164400
rect 168562 163200 168618 164400
rect 169390 163200 169446 164400
rect 170218 163200 170274 164400
rect 171138 163200 171194 164400
rect 171966 163200 172022 164400
rect 172532 163254 172744 163282
rect 166092 163146 166120 163200
rect 166000 163118 166120 163146
rect 166920 159934 166948 163200
rect 166908 159928 166960 159934
rect 166908 159870 166960 159876
rect 167748 159730 167776 163200
rect 168576 160342 168604 163200
rect 168564 160336 168616 160342
rect 168564 160278 168616 160284
rect 167736 159724 167788 159730
rect 167736 159666 167788 159672
rect 167000 159316 167052 159322
rect 167000 159258 167052 159264
rect 166080 158636 166132 158642
rect 166080 158578 166132 158584
rect 166540 158636 166592 158642
rect 166540 158578 166592 158584
rect 166092 158522 166120 158578
rect 166092 158506 166488 158522
rect 165988 158500 166040 158506
rect 166092 158500 166500 158506
rect 166092 158494 166448 158500
rect 165988 158442 166040 158448
rect 166448 158442 166500 158448
rect 166000 158386 166028 158442
rect 166552 158386 166580 158578
rect 166000 158358 166580 158386
rect 166448 157276 166500 157282
rect 166448 157218 166500 157224
rect 166172 157208 166224 157214
rect 166172 157150 166224 157156
rect 166264 157208 166316 157214
rect 166264 157150 166316 157156
rect 166184 156534 166212 157150
rect 166172 156528 166224 156534
rect 166172 156470 166224 156476
rect 166276 156466 166304 157150
rect 166460 156534 166488 157218
rect 166448 156528 166500 156534
rect 166448 156470 166500 156476
rect 166264 156460 166316 156466
rect 166264 156402 166316 156408
rect 166722 155544 166778 155553
rect 166722 155479 166778 155488
rect 166080 154284 166132 154290
rect 166080 154226 166132 154232
rect 165620 154148 165672 154154
rect 165620 154090 165672 154096
rect 164424 152788 164476 152794
rect 164424 152730 164476 152736
rect 164792 152108 164844 152114
rect 164792 152050 164844 152056
rect 164804 150226 164832 152050
rect 166092 150226 166120 154226
rect 166736 150226 166764 155479
rect 167012 152114 167040 159258
rect 167552 158432 167604 158438
rect 167552 158374 167604 158380
rect 167368 152856 167420 152862
rect 167368 152798 167420 152804
rect 167000 152108 167052 152114
rect 167000 152050 167052 152056
rect 167380 150226 167408 152798
rect 167564 151814 167592 158374
rect 169404 155514 169432 163200
rect 170232 159322 170260 163200
rect 171152 159798 171180 163200
rect 171140 159792 171192 159798
rect 171140 159734 171192 159740
rect 170220 159316 170272 159322
rect 170220 159258 170272 159264
rect 169760 159112 169812 159118
rect 169760 159054 169812 159060
rect 171784 159112 171836 159118
rect 171784 159054 171836 159060
rect 168656 155508 168708 155514
rect 168656 155450 168708 155456
rect 169392 155508 169444 155514
rect 169392 155450 169444 155456
rect 168378 155408 168434 155417
rect 168378 155343 168434 155352
rect 167564 151786 168052 151814
rect 168024 150226 168052 151786
rect 161630 149940 161658 150198
rect 162274 149940 162302 150198
rect 162918 149940 162946 150198
rect 163562 149940 163590 150198
rect 164206 149940 164234 150198
rect 164332 150204 164384 150210
rect 164804 150198 164878 150226
rect 164332 150146 164384 150152
rect 164850 149940 164878 150198
rect 165482 150204 165534 150210
rect 166092 150198 166166 150226
rect 166736 150198 166810 150226
rect 167380 150198 167454 150226
rect 168024 150198 168098 150226
rect 168392 150210 168420 155343
rect 168668 150226 168696 155450
rect 169772 151842 169800 159054
rect 171796 158778 171824 159054
rect 171784 158772 171836 158778
rect 171784 158714 171836 158720
rect 170404 158500 170456 158506
rect 170404 158442 170456 158448
rect 170220 157956 170272 157962
rect 170220 157898 170272 157904
rect 170036 157820 170088 157826
rect 170232 157808 170260 157898
rect 170088 157780 170260 157808
rect 170036 157762 170088 157768
rect 170416 157334 170444 158442
rect 171980 158438 172008 163200
rect 172152 159180 172204 159186
rect 172152 159122 172204 159128
rect 171968 158432 172020 158438
rect 171968 158374 172020 158380
rect 170496 157888 170548 157894
rect 170494 157856 170496 157865
rect 170548 157856 170550 157865
rect 170494 157791 170550 157800
rect 170324 157306 170444 157334
rect 169944 152176 169996 152182
rect 169944 152118 169996 152124
rect 169760 151836 169812 151842
rect 169760 151778 169812 151784
rect 169956 150226 169984 152118
rect 170324 151814 170352 157306
rect 171140 157208 171192 157214
rect 171140 157150 171192 157156
rect 170324 151786 170628 151814
rect 170600 150226 170628 151786
rect 165482 150146 165534 150152
rect 165494 149940 165522 150146
rect 166138 149940 166166 150198
rect 166782 149940 166810 150198
rect 167426 149940 167454 150198
rect 168070 149940 168098 150198
rect 168380 150204 168432 150210
rect 168668 150198 168742 150226
rect 168380 150146 168432 150152
rect 168714 149940 168742 150198
rect 169346 150204 169398 150210
rect 169956 150198 170030 150226
rect 170600 150198 170674 150226
rect 171152 150210 171180 157150
rect 171230 155272 171286 155281
rect 171230 155207 171286 155216
rect 171244 150226 171272 155207
rect 172164 152182 172192 159122
rect 172532 154222 172560 163254
rect 172716 163146 172744 163254
rect 172794 163200 172850 164400
rect 173622 163200 173678 164400
rect 173912 163254 174400 163282
rect 172808 163146 172836 163200
rect 172716 163118 172836 163146
rect 173348 160336 173400 160342
rect 173348 160278 173400 160284
rect 173256 159792 173308 159798
rect 173256 159734 173308 159740
rect 172900 158732 173204 158760
rect 172900 158574 172928 158732
rect 172980 158636 173032 158642
rect 173032 158596 173112 158624
rect 172980 158578 173032 158584
rect 172888 158568 172940 158574
rect 172888 158510 172940 158516
rect 172704 155644 172756 155650
rect 172704 155586 172756 155592
rect 172520 154216 172572 154222
rect 172520 154158 172572 154164
rect 172152 152176 172204 152182
rect 172152 152118 172204 152124
rect 172520 152040 172572 152046
rect 172520 151982 172572 151988
rect 172532 150226 172560 151982
rect 169346 150146 169398 150152
rect 169358 149940 169386 150146
rect 170002 149940 170030 150198
rect 170646 149940 170674 150198
rect 171140 150204 171192 150210
rect 171244 150198 171318 150226
rect 171140 150146 171192 150152
rect 171290 149940 171318 150198
rect 171922 150204 171974 150210
rect 172532 150198 172606 150226
rect 172716 150210 172744 155586
rect 173084 151814 173112 158596
rect 173176 158506 173204 158732
rect 173164 158500 173216 158506
rect 173164 158442 173216 158448
rect 173268 152454 173296 159734
rect 173360 158642 173388 160278
rect 173636 158778 173664 163200
rect 173624 158772 173676 158778
rect 173624 158714 173676 158720
rect 173348 158636 173400 158642
rect 173348 158578 173400 158584
rect 173912 152862 173940 163254
rect 174372 163146 174400 163254
rect 174450 163200 174506 164400
rect 175278 163200 175334 164400
rect 176106 163200 176162 164400
rect 177026 163200 177082 164400
rect 177854 163200 177910 164400
rect 178682 163200 178738 164400
rect 179510 163200 179566 164400
rect 180338 163200 180394 164400
rect 180812 163254 181116 163282
rect 174464 163146 174492 163200
rect 174372 163118 174492 163146
rect 175292 158506 175320 163200
rect 175188 158500 175240 158506
rect 175188 158442 175240 158448
rect 175280 158500 175332 158506
rect 175280 158442 175332 158448
rect 175200 158386 175228 158442
rect 175200 158358 175320 158386
rect 174450 157040 174506 157049
rect 174450 156975 174506 156984
rect 173900 152856 173952 152862
rect 173900 152798 173952 152804
rect 173256 152448 173308 152454
rect 173256 152390 173308 152396
rect 173084 151786 173204 151814
rect 173176 150226 173204 151786
rect 174464 150226 174492 156975
rect 175096 153128 175148 153134
rect 175096 153070 175148 153076
rect 175108 150226 175136 153070
rect 175292 151814 175320 158358
rect 176120 157334 176148 163200
rect 176660 159112 176712 159118
rect 176660 159054 176712 159060
rect 176120 157306 176332 157334
rect 176304 155650 176332 157306
rect 176292 155644 176344 155650
rect 176292 155586 176344 155592
rect 176384 155576 176436 155582
rect 176384 155518 176436 155524
rect 175292 151786 175780 151814
rect 175752 150226 175780 151786
rect 176396 150226 176424 155518
rect 176672 154290 176700 159054
rect 177040 157214 177068 163200
rect 177868 159798 177896 163200
rect 177856 159792 177908 159798
rect 177856 159734 177908 159740
rect 178696 158574 178724 163200
rect 179420 159860 179472 159866
rect 179420 159802 179472 159808
rect 178684 158568 178736 158574
rect 178684 158510 178736 158516
rect 179432 157826 179460 159802
rect 178040 157820 178092 157826
rect 178040 157762 178092 157768
rect 179420 157820 179472 157826
rect 179420 157762 179472 157768
rect 177028 157208 177080 157214
rect 177028 157150 177080 157156
rect 177026 155816 177082 155825
rect 177026 155751 177082 155760
rect 176660 154284 176712 154290
rect 176660 154226 176712 154232
rect 177040 150226 177068 155751
rect 177672 151972 177724 151978
rect 177672 151914 177724 151920
rect 177684 150226 177712 151914
rect 178052 151814 178080 157762
rect 178958 155680 179014 155689
rect 178958 155615 179014 155624
rect 178052 151786 178356 151814
rect 178328 150226 178356 151786
rect 178972 150226 179000 155615
rect 179524 155582 179552 163200
rect 180352 159118 180380 163200
rect 180340 159112 180392 159118
rect 180340 159054 180392 159060
rect 179512 155576 179564 155582
rect 179512 155518 179564 155524
rect 179696 154284 179748 154290
rect 179696 154226 179748 154232
rect 179708 153610 179736 154226
rect 179604 153604 179656 153610
rect 179604 153546 179656 153552
rect 179696 153604 179748 153610
rect 179696 153546 179748 153552
rect 179616 150226 179644 153546
rect 180812 153134 180840 163254
rect 181088 163146 181116 163254
rect 181166 163200 181222 164400
rect 181994 163200 182050 164400
rect 182192 163254 182864 163282
rect 181180 163146 181208 163200
rect 181088 163118 181208 163146
rect 182008 158710 182036 163200
rect 180892 158704 180944 158710
rect 180892 158646 180944 158652
rect 181996 158704 182048 158710
rect 181996 158646 182048 158652
rect 180800 153128 180852 153134
rect 180800 153070 180852 153076
rect 180248 152312 180300 152318
rect 180248 152254 180300 152260
rect 180260 150226 180288 152254
rect 180904 150226 180932 158646
rect 182088 156392 182140 156398
rect 182088 156334 182140 156340
rect 180984 155712 181036 155718
rect 180984 155654 181036 155660
rect 180996 151814 181024 155654
rect 180996 151786 181484 151814
rect 171922 150146 171974 150152
rect 171934 149940 171962 150146
rect 172578 149940 172606 150198
rect 172704 150204 172756 150210
rect 173176 150198 173250 150226
rect 172704 150146 172756 150152
rect 173222 149940 173250 150198
rect 173854 150204 173906 150210
rect 174464 150198 174538 150226
rect 175108 150198 175182 150226
rect 175752 150198 175826 150226
rect 176396 150198 176470 150226
rect 177040 150198 177114 150226
rect 177684 150198 177758 150226
rect 178328 150198 178402 150226
rect 178972 150198 179046 150226
rect 179616 150198 179690 150226
rect 180260 150198 180334 150226
rect 173854 150146 173906 150152
rect 173866 149940 173894 150146
rect 174510 149940 174538 150198
rect 175154 149940 175182 150198
rect 175798 149940 175826 150198
rect 176442 149940 176470 150198
rect 177086 149940 177114 150198
rect 177730 149940 177758 150198
rect 178374 149940 178402 150198
rect 179018 149940 179046 150198
rect 179662 149940 179690 150198
rect 180306 149940 180334 150198
rect 180858 150198 180932 150226
rect 181456 150226 181484 151786
rect 182100 150226 182128 156334
rect 182192 154290 182220 163254
rect 182836 163146 182864 163254
rect 182914 163200 182970 164400
rect 183742 163200 183798 164400
rect 184570 163200 184626 164400
rect 185398 163200 185454 164400
rect 186226 163200 186282 164400
rect 187054 163200 187110 164400
rect 187882 163200 187938 164400
rect 188802 163200 188858 164400
rect 189630 163200 189686 164400
rect 190458 163200 190514 164400
rect 191286 163200 191342 164400
rect 192114 163200 192170 164400
rect 192942 163200 192998 164400
rect 193770 163200 193826 164400
rect 194690 163200 194746 164400
rect 195518 163200 195574 164400
rect 196346 163200 196402 164400
rect 197174 163200 197230 164400
rect 198002 163200 198058 164400
rect 198830 163200 198886 164400
rect 199658 163200 199714 164400
rect 200578 163200 200634 164400
rect 201406 163200 201462 164400
rect 202234 163200 202290 164400
rect 203062 163200 203118 164400
rect 203890 163200 203946 164400
rect 204718 163200 204774 164400
rect 205100 163254 205496 163282
rect 182928 163146 182956 163200
rect 182836 163118 182956 163146
rect 183756 159050 183784 163200
rect 184584 159866 184612 163200
rect 184572 159860 184624 159866
rect 184572 159802 184624 159808
rect 184388 159248 184440 159254
rect 184388 159190 184440 159196
rect 183468 159044 183520 159050
rect 183468 158986 183520 158992
rect 183744 159044 183796 159050
rect 183744 158986 183796 158992
rect 182272 157956 182324 157962
rect 182272 157898 182324 157904
rect 182180 154284 182232 154290
rect 182180 154226 182232 154232
rect 181456 150198 181530 150226
rect 182100 150198 182174 150226
rect 182284 150210 182312 157898
rect 183480 152114 183508 158986
rect 184018 155952 184074 155961
rect 184018 155887 184074 155896
rect 182732 152108 182784 152114
rect 182732 152050 182784 152056
rect 183468 152108 183520 152114
rect 183468 152050 183520 152056
rect 182744 150226 182772 152050
rect 184032 150226 184060 155887
rect 184400 151978 184428 159190
rect 185412 157962 185440 163200
rect 185308 157956 185360 157962
rect 185308 157898 185360 157904
rect 185400 157956 185452 157962
rect 185400 157898 185452 157904
rect 185124 157888 185176 157894
rect 185124 157830 185176 157836
rect 185320 157842 185348 157898
rect 185136 157434 185164 157830
rect 185320 157814 185624 157842
rect 185308 157752 185360 157758
rect 185308 157694 185360 157700
rect 185320 157570 185348 157694
rect 185596 157690 185624 157814
rect 185676 157752 185728 157758
rect 185676 157694 185728 157700
rect 185584 157684 185636 157690
rect 185584 157626 185636 157632
rect 185688 157570 185716 157694
rect 185320 157542 185716 157570
rect 185136 157406 185440 157434
rect 184662 154456 184718 154465
rect 184662 154391 184718 154400
rect 184388 151972 184440 151978
rect 184388 151914 184440 151920
rect 184676 150226 184704 154391
rect 185308 151836 185360 151842
rect 185412 151814 185440 157406
rect 186240 155718 186268 163200
rect 186412 159928 186464 159934
rect 186412 159870 186464 159876
rect 186424 157334 186452 159870
rect 187068 159254 187096 163200
rect 187896 161474 187924 163200
rect 187896 161446 188016 161474
rect 187056 159248 187108 159254
rect 187056 159190 187108 159196
rect 186424 157306 186728 157334
rect 186320 155916 186372 155922
rect 186320 155858 186372 155864
rect 186412 155916 186464 155922
rect 186412 155858 186464 155864
rect 186228 155712 186280 155718
rect 186228 155654 186280 155660
rect 186332 155145 186360 155858
rect 186318 155136 186374 155145
rect 186318 155071 186374 155080
rect 186320 155032 186372 155038
rect 186424 155020 186452 155858
rect 186372 154992 186452 155020
rect 186320 154974 186372 154980
rect 186700 154902 186728 157306
rect 186872 155848 186924 155854
rect 186872 155790 186924 155796
rect 186780 155100 186832 155106
rect 186780 155042 186832 155048
rect 186412 154896 186464 154902
rect 186412 154838 186464 154844
rect 186688 154896 186740 154902
rect 186688 154838 186740 154844
rect 186424 154714 186452 154838
rect 186792 154714 186820 155042
rect 186424 154686 186820 154714
rect 185412 151786 185992 151814
rect 185308 151778 185360 151784
rect 185320 150226 185348 151778
rect 185964 150226 185992 151786
rect 186884 150226 186912 155790
rect 187238 155136 187294 155145
rect 187238 155071 187294 155080
rect 180858 149940 180886 150198
rect 181502 149940 181530 150198
rect 182146 149940 182174 150198
rect 182272 150204 182324 150210
rect 182744 150198 182818 150226
rect 182272 150146 182324 150152
rect 182790 149940 182818 150198
rect 183422 150204 183474 150210
rect 184032 150198 184106 150226
rect 184676 150198 184750 150226
rect 185320 150198 185394 150226
rect 185964 150198 186038 150226
rect 183422 150146 183474 150152
rect 183434 149940 183462 150146
rect 184078 149940 184106 150198
rect 184722 149940 184750 150198
rect 185366 149940 185394 150198
rect 186010 149940 186038 150198
rect 186654 150198 186912 150226
rect 186654 149940 186682 150198
rect 187252 150090 187280 155071
rect 187884 152992 187936 152998
rect 187884 152934 187936 152940
rect 187896 150090 187924 152934
rect 187988 152318 188016 161446
rect 188816 157894 188844 163200
rect 188804 157888 188856 157894
rect 188804 157830 188856 157836
rect 188528 157752 188580 157758
rect 188528 157694 188580 157700
rect 188252 154488 188304 154494
rect 188304 154436 188476 154442
rect 188252 154430 188476 154436
rect 188264 154426 188476 154430
rect 188264 154420 188488 154426
rect 188264 154414 188436 154420
rect 188436 154362 188488 154368
rect 187976 152312 188028 152318
rect 187976 152254 188028 152260
rect 188540 150226 188568 157694
rect 189644 155854 189672 163200
rect 190472 157758 190500 163200
rect 191300 159934 191328 163200
rect 191656 160064 191708 160070
rect 191656 160006 191708 160012
rect 191472 159996 191524 160002
rect 191472 159938 191524 159944
rect 191288 159928 191340 159934
rect 191288 159870 191340 159876
rect 190644 157820 190696 157826
rect 190644 157762 190696 157768
rect 190460 157752 190512 157758
rect 190460 157694 190512 157700
rect 190656 157334 190684 157762
rect 190656 157306 191144 157334
rect 189632 155848 189684 155854
rect 189632 155790 189684 155796
rect 189172 155168 189224 155174
rect 189172 155110 189224 155116
rect 188540 150198 188614 150226
rect 187252 150062 187326 150090
rect 187896 150062 187970 150090
rect 187298 149940 187326 150062
rect 187942 149940 187970 150062
rect 188586 149940 188614 150198
rect 189184 150090 189212 155110
rect 189816 154488 189868 154494
rect 189816 154430 189868 154436
rect 191012 154488 191064 154494
rect 191012 154430 191064 154436
rect 189828 150090 189856 154430
rect 191024 153406 191052 154430
rect 191012 153400 191064 153406
rect 191012 153342 191064 153348
rect 190460 152176 190512 152182
rect 190460 152118 190512 152124
rect 190472 150090 190500 152118
rect 191116 150226 191144 157306
rect 191484 152046 191512 159938
rect 191668 153406 191696 160006
rect 192128 157282 192156 163200
rect 192116 157276 192168 157282
rect 192116 157218 192168 157224
rect 192956 155922 192984 163200
rect 193784 159186 193812 163200
rect 193772 159180 193824 159186
rect 193772 159122 193824 159128
rect 194704 158982 194732 163200
rect 194140 158976 194192 158982
rect 194140 158918 194192 158924
rect 194692 158976 194744 158982
rect 194692 158918 194744 158924
rect 193220 157616 193272 157622
rect 193220 157558 193272 157564
rect 193232 157334 193260 157558
rect 193232 157306 193720 157334
rect 192852 155916 192904 155922
rect 192852 155858 192904 155864
rect 192944 155916 192996 155922
rect 192944 155858 192996 155864
rect 192864 155174 192892 155858
rect 192852 155168 192904 155174
rect 192852 155110 192904 155116
rect 191748 155032 191800 155038
rect 191748 154974 191800 154980
rect 191656 153400 191708 153406
rect 191656 153342 191708 153348
rect 191472 152040 191524 152046
rect 191472 151982 191524 151988
rect 191116 150198 191190 150226
rect 189184 150062 189258 150090
rect 189828 150062 189902 150090
rect 190472 150062 190546 150090
rect 189230 149940 189258 150062
rect 189874 149940 189902 150062
rect 190518 149940 190546 150062
rect 191162 149940 191190 150198
rect 191760 150090 191788 154974
rect 192390 153776 192446 153785
rect 192390 153711 192446 153720
rect 192404 150090 192432 153711
rect 193036 152924 193088 152930
rect 193036 152866 193088 152872
rect 193048 150090 193076 152866
rect 193692 150226 193720 157306
rect 194152 152182 194180 158918
rect 195428 158908 195480 158914
rect 195428 158850 195480 158856
rect 194968 156324 195020 156330
rect 194968 156266 195020 156272
rect 194324 155168 194376 155174
rect 194324 155110 194376 155116
rect 194140 152176 194192 152182
rect 194140 152118 194192 152124
rect 193692 150198 193766 150226
rect 191760 150062 191834 150090
rect 192404 150062 192478 150090
rect 193048 150062 193122 150090
rect 191806 149940 191834 150062
rect 192450 149940 192478 150062
rect 193094 149940 193122 150062
rect 193738 149940 193766 150198
rect 194336 150090 194364 155110
rect 194980 150090 195008 156266
rect 195440 152998 195468 158850
rect 195532 157826 195560 163200
rect 195520 157820 195572 157826
rect 195520 157762 195572 157768
rect 196256 156256 196308 156262
rect 196256 156198 196308 156204
rect 195428 152992 195480 152998
rect 195428 152934 195480 152940
rect 195612 151972 195664 151978
rect 195612 151914 195664 151920
rect 195624 150090 195652 151914
rect 196268 150090 196296 156198
rect 196360 155174 196388 163200
rect 197188 160070 197216 163200
rect 197176 160064 197228 160070
rect 197176 160006 197228 160012
rect 198016 160002 198044 163200
rect 198004 159996 198056 160002
rect 198004 159938 198056 159944
rect 197268 158840 197320 158846
rect 197268 158782 197320 158788
rect 196348 155168 196400 155174
rect 196348 155110 196400 155116
rect 197280 153542 197308 158782
rect 197360 158772 197412 158778
rect 197360 158714 197412 158720
rect 197372 157622 197400 158714
rect 198738 158536 198794 158545
rect 198738 158471 198794 158480
rect 197360 157616 197412 157622
rect 197360 157558 197412 157564
rect 198464 154488 198516 154494
rect 198464 154430 198516 154436
rect 197544 154420 197596 154426
rect 197544 154362 197596 154368
rect 196900 153536 196952 153542
rect 196900 153478 196952 153484
rect 197268 153536 197320 153542
rect 197268 153478 197320 153484
rect 196912 150090 196940 153478
rect 197556 150090 197584 154362
rect 198476 153746 198504 154430
rect 198464 153740 198516 153746
rect 198464 153682 198516 153688
rect 198556 153740 198608 153746
rect 198556 153682 198608 153688
rect 198568 153270 198596 153682
rect 198648 153536 198700 153542
rect 198648 153478 198700 153484
rect 198660 153270 198688 153478
rect 198556 153264 198608 153270
rect 198556 153206 198608 153212
rect 198648 153264 198700 153270
rect 198648 153206 198700 153212
rect 198188 153060 198240 153066
rect 198188 153002 198240 153008
rect 198200 150090 198228 153002
rect 198752 150226 198780 158471
rect 198844 156398 198872 163200
rect 198924 159316 198976 159322
rect 198924 159258 198976 159264
rect 198832 156392 198884 156398
rect 198832 156334 198884 156340
rect 198936 153542 198964 159258
rect 199672 155106 199700 163200
rect 200592 158778 200620 163200
rect 201420 159322 201448 163200
rect 202248 161474 202276 163200
rect 202248 161446 202368 161474
rect 201408 159316 201460 159322
rect 201408 159258 201460 159264
rect 201408 159044 201460 159050
rect 201408 158986 201460 158992
rect 200580 158772 200632 158778
rect 200580 158714 200632 158720
rect 200856 156392 200908 156398
rect 200856 156334 200908 156340
rect 200672 156256 200724 156262
rect 200408 156204 200672 156210
rect 200408 156198 200724 156204
rect 200408 156194 200712 156198
rect 200396 156188 200712 156194
rect 200448 156182 200712 156188
rect 200396 156130 200448 156136
rect 200868 156058 200896 156334
rect 201316 156256 201368 156262
rect 201316 156198 201368 156204
rect 200856 156052 200908 156058
rect 200856 155994 200908 156000
rect 199660 155100 199712 155106
rect 199660 155042 199712 155048
rect 200120 155032 200172 155038
rect 200120 154974 200172 154980
rect 198924 153536 198976 153542
rect 198924 153478 198976 153484
rect 199476 153468 199528 153474
rect 199476 153410 199528 153416
rect 198752 150198 198918 150226
rect 194336 150062 194410 150090
rect 194980 150062 195054 150090
rect 195624 150062 195698 150090
rect 196268 150062 196342 150090
rect 196912 150062 196986 150090
rect 197556 150062 197630 150090
rect 198200 150062 198274 150090
rect 194382 149940 194410 150062
rect 195026 149940 195054 150062
rect 195670 149940 195698 150062
rect 196314 149940 196342 150062
rect 196958 149940 196986 150062
rect 197602 149940 197630 150062
rect 198246 149940 198274 150062
rect 198890 149940 198918 150198
rect 199488 150090 199516 153410
rect 200132 150090 200160 154974
rect 200212 153400 200264 153406
rect 200264 153348 200620 153354
rect 200212 153342 200620 153348
rect 200224 153338 200620 153342
rect 200224 153332 200632 153338
rect 200224 153326 200580 153332
rect 200580 153274 200632 153280
rect 200764 152108 200816 152114
rect 200764 152050 200816 152056
rect 200776 150090 200804 152050
rect 201328 150226 201356 156198
rect 201420 153270 201448 158986
rect 202340 156126 202368 161446
rect 203076 156262 203104 163200
rect 203904 159050 203932 163200
rect 204732 159361 204760 163200
rect 204718 159352 204774 159361
rect 204718 159287 204774 159296
rect 204904 159112 204956 159118
rect 204904 159054 204956 159060
rect 203892 159044 203944 159050
rect 203892 158986 203944 158992
rect 204168 158976 204220 158982
rect 204168 158918 204220 158924
rect 203984 157548 204036 157554
rect 203984 157490 204036 157496
rect 203064 156256 203116 156262
rect 203064 156198 203116 156204
rect 202328 156120 202380 156126
rect 202328 156062 202380 156068
rect 202696 154556 202748 154562
rect 202696 154498 202748 154504
rect 202052 154420 202104 154426
rect 202052 154362 202104 154368
rect 201408 153264 201460 153270
rect 201408 153206 201460 153212
rect 201328 150198 201494 150226
rect 199488 150062 199562 150090
rect 200132 150062 200206 150090
rect 200776 150062 200850 150090
rect 199534 149940 199562 150062
rect 200178 149940 200206 150062
rect 200822 149940 200850 150062
rect 201466 149940 201494 150198
rect 202064 150090 202092 154362
rect 202708 150090 202736 154498
rect 203340 151904 203392 151910
rect 203340 151846 203392 151852
rect 203352 150090 203380 151846
rect 203996 150226 204024 157490
rect 204180 153066 204208 158918
rect 204916 157554 204944 159054
rect 204904 157548 204956 157554
rect 204904 157490 204956 157496
rect 204628 155780 204680 155786
rect 204628 155722 204680 155728
rect 204168 153060 204220 153066
rect 204168 153002 204220 153008
rect 203996 150198 204070 150226
rect 202064 150062 202138 150090
rect 202708 150062 202782 150090
rect 203352 150062 203426 150090
rect 202110 149940 202138 150062
rect 202754 149940 202782 150062
rect 203398 149940 203426 150062
rect 204042 149940 204070 150198
rect 204640 150090 204668 155722
rect 205100 154426 205128 163254
rect 205468 163146 205496 163254
rect 205546 163200 205602 164400
rect 206466 163200 206522 164400
rect 207294 163200 207350 164400
rect 208122 163200 208178 164400
rect 208412 163254 208900 163282
rect 205560 163146 205588 163200
rect 205468 163118 205588 163146
rect 206480 155786 206508 163200
rect 207020 160064 207072 160070
rect 207020 160006 207072 160012
rect 206560 157480 206612 157486
rect 206560 157422 206612 157428
rect 206468 155780 206520 155786
rect 206468 155722 206520 155728
rect 205088 154420 205140 154426
rect 205088 154362 205140 154368
rect 205272 154352 205324 154358
rect 205272 154294 205324 154300
rect 205284 150090 205312 154294
rect 205916 153196 205968 153202
rect 205916 153138 205968 153144
rect 205928 150226 205956 153138
rect 206572 150226 206600 157422
rect 207032 155038 207060 160006
rect 207308 158982 207336 163200
rect 207296 158976 207348 158982
rect 207296 158918 207348 158924
rect 208136 158846 208164 163200
rect 208124 158840 208176 158846
rect 208124 158782 208176 158788
rect 207202 157176 207258 157185
rect 207202 157111 207258 157120
rect 207020 155032 207072 155038
rect 207020 154974 207072 154980
rect 207216 150226 207244 157111
rect 208412 154358 208440 163254
rect 208872 163146 208900 163254
rect 208950 163200 209006 164400
rect 209778 163200 209834 164400
rect 210606 163200 210662 164400
rect 211434 163200 211490 164400
rect 211540 163254 212304 163282
rect 208964 163146 208992 163200
rect 208872 163118 208992 163146
rect 209792 156398 209820 163200
rect 210620 158914 210648 163200
rect 211448 160070 211476 163200
rect 211436 160064 211488 160070
rect 211436 160006 211488 160012
rect 210608 158908 210660 158914
rect 210608 158850 210660 158856
rect 209780 156392 209832 156398
rect 209780 156334 209832 156340
rect 209136 156324 209188 156330
rect 209136 156266 209188 156272
rect 208400 154352 208452 154358
rect 208400 154294 208452 154300
rect 207848 153468 207900 153474
rect 207848 153410 207900 153416
rect 207940 153468 207992 153474
rect 207940 153410 207992 153416
rect 207860 150226 207888 153410
rect 207952 153270 207980 153410
rect 207940 153264 207992 153270
rect 207940 153206 207992 153212
rect 208492 152040 208544 152046
rect 208492 151982 208544 151988
rect 208504 150226 208532 151982
rect 209148 150226 209176 156266
rect 211252 154964 211304 154970
rect 211252 154906 211304 154912
rect 210424 154488 210476 154494
rect 210424 154430 210476 154436
rect 209780 153740 209832 153746
rect 209780 153682 209832 153688
rect 209792 150226 209820 153682
rect 210436 150226 210464 154430
rect 211068 152380 211120 152386
rect 211068 152322 211120 152328
rect 211080 150226 211108 152322
rect 205928 150198 206002 150226
rect 206572 150198 206646 150226
rect 207216 150198 207290 150226
rect 207860 150198 207934 150226
rect 208504 150198 208578 150226
rect 209148 150198 209222 150226
rect 209792 150198 209866 150226
rect 210436 150198 210510 150226
rect 211080 150198 211154 150226
rect 211264 150210 211292 154906
rect 211540 153785 211568 163254
rect 212276 163146 212304 163254
rect 212354 163200 212410 164400
rect 213182 163200 213238 164400
rect 213288 163254 213868 163282
rect 212368 163146 212396 163200
rect 212276 163118 212396 163146
rect 213196 163146 213224 163200
rect 213288 163146 213316 163254
rect 213196 163118 213316 163146
rect 213736 159316 213788 159322
rect 213736 159258 213788 159264
rect 212724 159044 212776 159050
rect 212724 158986 212776 158992
rect 212448 158840 212500 158846
rect 212448 158782 212500 158788
rect 211804 156664 211856 156670
rect 211804 156606 211856 156612
rect 211816 156194 211844 156606
rect 211620 156188 211672 156194
rect 211620 156130 211672 156136
rect 211804 156188 211856 156194
rect 211804 156130 211856 156136
rect 211526 153776 211582 153785
rect 211526 153711 211582 153720
rect 211632 150226 211660 156130
rect 212460 152930 212488 158782
rect 212540 156732 212592 156738
rect 212540 156674 212592 156680
rect 212552 156330 212580 156674
rect 212540 156324 212592 156330
rect 212540 156266 212592 156272
rect 212448 152924 212500 152930
rect 212448 152866 212500 152872
rect 212736 152114 212764 158986
rect 212908 153808 212960 153814
rect 212908 153750 212960 153756
rect 212724 152108 212776 152114
rect 212724 152050 212776 152056
rect 212920 150226 212948 153750
rect 213552 152176 213604 152182
rect 213552 152118 213604 152124
rect 213564 150226 213592 152118
rect 213748 151978 213776 159258
rect 213840 156602 213868 163254
rect 214010 163200 214066 164400
rect 214838 163200 214894 164400
rect 215312 163254 215616 163282
rect 214024 159322 214052 163200
rect 214012 159316 214064 159322
rect 214012 159258 214064 159264
rect 214564 159248 214616 159254
rect 214564 159190 214616 159196
rect 213828 156596 213880 156602
rect 213828 156538 213880 156544
rect 213920 156188 213972 156194
rect 213920 156130 213972 156136
rect 213736 151972 213788 151978
rect 213736 151914 213788 151920
rect 213932 151814 213960 156130
rect 214576 154970 214604 159190
rect 214852 158846 214880 163200
rect 214840 158840 214892 158846
rect 214840 158782 214892 158788
rect 214840 155304 214892 155310
rect 214840 155246 214892 155252
rect 214564 154964 214616 154970
rect 214564 154906 214616 154912
rect 213932 151786 214236 151814
rect 214208 150226 214236 151786
rect 214852 150226 214880 155246
rect 215312 154494 215340 163254
rect 215588 163146 215616 163254
rect 215666 163200 215722 164400
rect 216494 163200 216550 164400
rect 217322 163200 217378 164400
rect 218242 163200 218298 164400
rect 218348 163254 219020 163282
rect 215680 163146 215708 163200
rect 215588 163118 215708 163146
rect 215392 158908 215444 158914
rect 215392 158850 215444 158856
rect 215300 154488 215352 154494
rect 215300 154430 215352 154436
rect 215404 153202 215432 158850
rect 215484 156732 215536 156738
rect 215484 156674 215536 156680
rect 215392 153196 215444 153202
rect 215392 153138 215444 153144
rect 215496 150226 215524 156674
rect 216508 156670 216536 163200
rect 217336 158914 217364 163200
rect 218256 159254 218284 163200
rect 218244 159248 218296 159254
rect 218244 159190 218296 159196
rect 218060 159180 218112 159186
rect 218060 159122 218112 159128
rect 217324 158908 217376 158914
rect 217324 158850 217376 158856
rect 216496 156664 216548 156670
rect 216496 156606 216548 156612
rect 218072 156330 218100 159122
rect 216772 156324 216824 156330
rect 216772 156266 216824 156272
rect 218060 156324 218112 156330
rect 218060 156266 218112 156272
rect 216128 152516 216180 152522
rect 216128 152458 216180 152464
rect 216140 150226 216168 152458
rect 216784 150226 216812 156266
rect 217416 155236 217468 155242
rect 217416 155178 217468 155184
rect 217428 150226 217456 155178
rect 218348 154562 218376 163254
rect 218992 163146 219020 163254
rect 219070 163200 219126 164400
rect 219898 163200 219954 164400
rect 220726 163200 220782 164400
rect 221554 163200 221610 164400
rect 222382 163200 222438 164400
rect 223210 163200 223266 164400
rect 224130 163200 224186 164400
rect 224958 163200 225014 164400
rect 225248 163254 225736 163282
rect 219084 163146 219112 163200
rect 218992 163118 219112 163146
rect 219348 158024 219400 158030
rect 219348 157966 219400 157972
rect 218336 154556 218388 154562
rect 218336 154498 218388 154504
rect 218060 153672 218112 153678
rect 218060 153614 218112 153620
rect 218072 150226 218100 153614
rect 218704 152992 218756 152998
rect 218704 152934 218756 152940
rect 218716 150226 218744 152934
rect 219360 150226 219388 157966
rect 219912 156738 219940 163200
rect 220740 159186 220768 163200
rect 220728 159180 220780 159186
rect 220728 159122 220780 159128
rect 220360 158908 220412 158914
rect 220360 158850 220412 158856
rect 219992 157344 220044 157350
rect 219992 157286 220044 157292
rect 219900 156732 219952 156738
rect 219900 156674 219952 156680
rect 219900 154012 219952 154018
rect 219900 153954 219952 153960
rect 204640 150062 204714 150090
rect 205284 150062 205358 150090
rect 204686 149940 204714 150062
rect 205330 149940 205358 150062
rect 205974 149940 206002 150198
rect 206618 149940 206646 150198
rect 207262 149940 207290 150198
rect 207906 149940 207934 150198
rect 208550 149940 208578 150198
rect 209194 149940 209222 150198
rect 209838 149940 209866 150198
rect 210482 149940 210510 150198
rect 211126 149940 211154 150198
rect 211252 150204 211304 150210
rect 211632 150198 211706 150226
rect 211252 150146 211304 150152
rect 211678 149940 211706 150198
rect 212310 150204 212362 150210
rect 212920 150198 212994 150226
rect 213564 150198 213638 150226
rect 214208 150198 214282 150226
rect 214852 150198 214926 150226
rect 215496 150198 215570 150226
rect 216140 150198 216214 150226
rect 216784 150198 216858 150226
rect 217428 150198 217502 150226
rect 218072 150198 218146 150226
rect 218716 150198 218790 150226
rect 219360 150198 219434 150226
rect 212310 150146 212362 150152
rect 212322 149940 212350 150146
rect 212966 149940 212994 150198
rect 213610 149940 213638 150198
rect 214254 149940 214282 150198
rect 214898 149940 214926 150198
rect 215542 149940 215570 150198
rect 216186 149940 216214 150198
rect 216830 149940 216858 150198
rect 217474 149940 217502 150198
rect 218118 149940 218146 150198
rect 218762 149940 218790 150198
rect 219406 149940 219434 150198
rect 219912 150192 219940 153954
rect 220004 151814 220032 157286
rect 220372 152998 220400 158850
rect 221568 158846 221596 163200
rect 221464 158840 221516 158846
rect 221464 158782 221516 158788
rect 221556 158840 221608 158846
rect 221556 158782 221608 158788
rect 221372 156868 221424 156874
rect 221372 156810 221424 156816
rect 220360 152992 220412 152998
rect 220360 152934 220412 152940
rect 221280 152244 221332 152250
rect 221280 152186 221332 152192
rect 220004 151786 220676 151814
rect 220648 150226 220676 151786
rect 221292 150226 221320 152186
rect 221384 151814 221412 156810
rect 221476 152250 221504 158782
rect 222396 154018 222424 163200
rect 222568 156936 222620 156942
rect 222568 156878 222620 156884
rect 222384 154012 222436 154018
rect 222384 153954 222436 153960
rect 221464 152244 221516 152250
rect 221464 152186 221516 152192
rect 221384 151786 221964 151814
rect 221936 150226 221964 151786
rect 222580 150226 222608 156878
rect 223224 156874 223252 163200
rect 223580 159384 223632 159390
rect 223580 159326 223632 159332
rect 223212 156868 223264 156874
rect 223212 156810 223264 156816
rect 223212 153944 223264 153950
rect 223212 153886 223264 153892
rect 223224 150226 223252 153886
rect 223592 151814 223620 159326
rect 224144 159118 224172 163200
rect 224972 159390 225000 163200
rect 224960 159384 225012 159390
rect 224960 159326 225012 159332
rect 224132 159112 224184 159118
rect 224132 159054 224184 159060
rect 224592 158840 224644 158846
rect 224592 158782 224644 158788
rect 224132 157004 224184 157010
rect 224132 156946 224184 156952
rect 224144 151814 224172 156946
rect 224604 152386 224632 158782
rect 224960 158772 225012 158778
rect 224960 158714 225012 158720
rect 224972 157010 225000 158714
rect 224960 157004 225012 157010
rect 224960 156946 225012 156952
rect 225144 156800 225196 156806
rect 225144 156742 225196 156748
rect 225052 156528 225104 156534
rect 225052 156470 225104 156476
rect 224592 152380 224644 152386
rect 224592 152322 224644 152328
rect 223592 151786 223896 151814
rect 224144 151786 224540 151814
rect 223868 150226 223896 151786
rect 224512 150226 224540 151786
rect 220648 150198 220722 150226
rect 221292 150198 221366 150226
rect 221936 150198 222010 150226
rect 222580 150198 222654 150226
rect 223224 150198 223298 150226
rect 223868 150198 223942 150226
rect 224512 150198 224586 150226
rect 225064 150210 225092 156470
rect 225156 150226 225184 156742
rect 225248 153950 225276 163254
rect 225708 163146 225736 163254
rect 225786 163200 225842 164400
rect 226614 163200 226670 164400
rect 227442 163200 227498 164400
rect 227732 163254 228220 163282
rect 225800 163146 225828 163200
rect 225708 163118 225828 163146
rect 225328 159520 225380 159526
rect 225328 159462 225380 159468
rect 225236 153944 225288 153950
rect 225236 153886 225288 153892
rect 225340 152114 225368 159462
rect 226628 156942 226656 163200
rect 227076 157412 227128 157418
rect 227076 157354 227128 157360
rect 226616 156936 226668 156942
rect 226616 156878 226668 156884
rect 226432 152584 226484 152590
rect 226432 152526 226484 152532
rect 225328 152108 225380 152114
rect 225328 152050 225380 152056
rect 226444 150226 226472 152526
rect 227088 150226 227116 157354
rect 227456 152425 227484 163200
rect 227732 152522 227760 163254
rect 228192 163146 228220 163254
rect 228270 163200 228326 164400
rect 229098 163200 229154 164400
rect 230018 163200 230074 164400
rect 230846 163200 230902 164400
rect 231674 163200 231730 164400
rect 231872 163254 232452 163282
rect 228284 163146 228312 163200
rect 228192 163118 228312 163146
rect 228364 156460 228416 156466
rect 228364 156402 228416 156408
rect 227812 155372 227864 155378
rect 227812 155314 227864 155320
rect 227720 152516 227772 152522
rect 227720 152458 227772 152464
rect 227442 152416 227498 152425
rect 227442 152351 227498 152360
rect 227824 150226 227852 155314
rect 219912 150164 220078 150192
rect 220050 149940 220078 150164
rect 220694 149940 220722 150198
rect 221338 149940 221366 150198
rect 221982 149940 222010 150198
rect 222626 149940 222654 150198
rect 223270 149940 223298 150198
rect 223914 149940 223942 150198
rect 224558 149940 224586 150198
rect 225052 150204 225104 150210
rect 225156 150198 225230 150226
rect 225052 150146 225104 150152
rect 225202 149940 225230 150198
rect 225834 150204 225886 150210
rect 226444 150198 226518 150226
rect 227088 150198 227162 150226
rect 225834 150146 225886 150152
rect 225846 149940 225874 150146
rect 226490 149940 226518 150198
rect 227134 149940 227162 150198
rect 227778 150198 227852 150226
rect 228376 150226 228404 156402
rect 229112 153746 229140 163200
rect 230032 156806 230060 163200
rect 230860 159050 230888 163200
rect 231688 159526 231716 163200
rect 231676 159520 231728 159526
rect 231676 159462 231728 159468
rect 230848 159044 230900 159050
rect 230848 158986 230900 158992
rect 230756 158976 230808 158982
rect 230756 158918 230808 158924
rect 230020 156800 230072 156806
rect 230020 156742 230072 156748
rect 230768 156262 230796 158918
rect 230756 156256 230808 156262
rect 230756 156198 230808 156204
rect 229652 155984 229704 155990
rect 229652 155926 229704 155932
rect 229192 155440 229244 155446
rect 229192 155382 229244 155388
rect 229100 153740 229152 153746
rect 229100 153682 229152 153688
rect 229008 152108 229060 152114
rect 229008 152050 229060 152056
rect 229020 150226 229048 152050
rect 228376 150198 228450 150226
rect 229020 150198 229094 150226
rect 229204 150210 229232 155382
rect 229664 150226 229692 155926
rect 231872 153814 231900 163254
rect 232424 163146 232452 163254
rect 232502 163200 232558 164400
rect 233330 163200 233386 164400
rect 234158 163200 234214 164400
rect 234986 163200 235042 164400
rect 235092 163254 235856 163282
rect 232516 163146 232544 163200
rect 232424 163118 232544 163146
rect 233240 159452 233292 159458
rect 233240 159394 233292 159400
rect 231952 158092 232004 158098
rect 231952 158034 232004 158040
rect 231860 153808 231912 153814
rect 231860 153750 231912 153756
rect 230940 153604 230992 153610
rect 230940 153546 230992 153552
rect 230952 150226 230980 153546
rect 231584 152720 231636 152726
rect 231584 152662 231636 152668
rect 231596 150226 231624 152662
rect 231964 151814 231992 158034
rect 232872 154828 232924 154834
rect 232872 154770 232924 154776
rect 231964 151786 232268 151814
rect 232240 150226 232268 151786
rect 232884 150226 232912 154770
rect 227778 149940 227806 150198
rect 228422 149940 228450 150198
rect 229066 149940 229094 150198
rect 229192 150204 229244 150210
rect 229664 150198 229738 150226
rect 229192 150146 229244 150152
rect 229710 149940 229738 150198
rect 230342 150204 230394 150210
rect 230952 150198 231026 150226
rect 231596 150198 231670 150226
rect 232240 150198 232314 150226
rect 232884 150198 232958 150226
rect 233252 150210 233280 159394
rect 233344 155242 233372 163200
rect 233516 157140 233568 157146
rect 233516 157082 233568 157088
rect 233332 155236 233384 155242
rect 233332 155178 233384 155184
rect 233528 150226 233556 157082
rect 234172 152590 234200 163200
rect 235000 159458 235028 163200
rect 234988 159452 235040 159458
rect 234988 159394 235040 159400
rect 234804 157072 234856 157078
rect 234804 157014 234856 157020
rect 234160 152584 234212 152590
rect 234160 152526 234212 152532
rect 234816 150226 234844 157014
rect 235092 153678 235120 163254
rect 235828 163146 235856 163254
rect 235906 163200 235962 164400
rect 236734 163200 236790 164400
rect 237562 163200 237618 164400
rect 238390 163200 238446 164400
rect 238864 163254 239168 163282
rect 235920 163146 235948 163200
rect 235828 163118 235948 163146
rect 236748 158030 236776 163200
rect 237576 158982 237604 163200
rect 237564 158976 237616 158982
rect 237564 158918 237616 158924
rect 238404 158914 238432 163200
rect 238392 158908 238444 158914
rect 238392 158850 238444 158856
rect 237380 158160 237432 158166
rect 237380 158102 237432 158108
rect 236736 158024 236788 158030
rect 236736 157966 236788 157972
rect 236092 157684 236144 157690
rect 236092 157626 236144 157632
rect 235448 153876 235500 153882
rect 235448 153818 235500 153824
rect 235080 153672 235132 153678
rect 235080 153614 235132 153620
rect 235460 150226 235488 153818
rect 236104 150226 236132 157626
rect 236736 152652 236788 152658
rect 236736 152594 236788 152600
rect 236748 150226 236776 152594
rect 237392 150226 237420 158102
rect 238024 154760 238076 154766
rect 238024 154702 238076 154708
rect 238036 150226 238064 154702
rect 238864 153610 238892 163254
rect 239140 163146 239168 163254
rect 239218 163200 239274 164400
rect 240046 163200 240102 164400
rect 240874 163200 240930 164400
rect 241794 163200 241850 164400
rect 241900 163254 242572 163282
rect 239232 163146 239260 163200
rect 239140 163118 239260 163146
rect 239312 159588 239364 159594
rect 239312 159530 239364 159536
rect 238944 158228 238996 158234
rect 238944 158170 238996 158176
rect 238852 153604 238904 153610
rect 238852 153546 238904 153552
rect 238668 153332 238720 153338
rect 238668 153274 238720 153280
rect 238680 150226 238708 153274
rect 230342 150146 230394 150152
rect 230354 149940 230382 150146
rect 230998 149940 231026 150198
rect 231642 149940 231670 150198
rect 232286 149940 232314 150198
rect 232930 149940 232958 150198
rect 233240 150204 233292 150210
rect 233528 150198 233602 150226
rect 233240 150146 233292 150152
rect 233574 149940 233602 150198
rect 234206 150204 234258 150210
rect 234816 150198 234890 150226
rect 235460 150198 235534 150226
rect 236104 150198 236178 150226
rect 236748 150198 236822 150226
rect 237392 150198 237466 150226
rect 238036 150198 238110 150226
rect 238680 150198 238754 150226
rect 238956 150210 238984 158170
rect 239324 150226 239352 159530
rect 240060 155310 240088 163200
rect 240324 159656 240376 159662
rect 240324 159598 240376 159604
rect 240048 155304 240100 155310
rect 240048 155246 240100 155252
rect 240336 152726 240364 159598
rect 240888 158778 240916 163200
rect 241808 159662 241836 163200
rect 241796 159656 241848 159662
rect 241796 159598 241848 159604
rect 240876 158772 240928 158778
rect 240876 158714 240928 158720
rect 240600 154692 240652 154698
rect 240600 154634 240652 154640
rect 240324 152720 240376 152726
rect 240324 152662 240376 152668
rect 240612 150226 240640 154634
rect 241244 154080 241296 154086
rect 241244 154022 241296 154028
rect 241256 150226 241284 154022
rect 241900 153882 241928 163254
rect 242544 163146 242572 163254
rect 242622 163200 242678 164400
rect 243450 163200 243506 164400
rect 244278 163200 244334 164400
rect 244476 163254 245056 163282
rect 242636 163146 242664 163200
rect 242544 163118 242664 163146
rect 242440 158908 242492 158914
rect 242440 158850 242492 158856
rect 242072 158296 242124 158302
rect 242072 158238 242124 158244
rect 241888 153876 241940 153882
rect 241888 153818 241940 153824
rect 241888 152720 241940 152726
rect 241888 152662 241940 152668
rect 241900 150226 241928 152662
rect 242084 151814 242112 158238
rect 242452 152046 242480 158850
rect 243360 158772 243412 158778
rect 243360 158714 243412 158720
rect 243084 154624 243136 154630
rect 243084 154566 243136 154572
rect 242440 152040 242492 152046
rect 242440 151982 242492 151988
rect 242084 151786 242480 151814
rect 242452 150226 242480 151786
rect 243096 150226 243124 154566
rect 243372 152114 243400 158714
rect 243464 158098 243492 163200
rect 244292 158914 244320 163200
rect 244280 158908 244332 158914
rect 244280 158850 244332 158856
rect 243452 158092 243504 158098
rect 243452 158034 243504 158040
rect 243728 153400 243780 153406
rect 243728 153342 243780 153348
rect 243360 152108 243412 152114
rect 243360 152050 243412 152056
rect 243740 150226 243768 153342
rect 244372 152788 244424 152794
rect 244372 152730 244424 152736
rect 244384 150226 244412 152730
rect 244476 152658 244504 163254
rect 245028 163146 245056 163254
rect 245106 163200 245162 164400
rect 245934 163200 245990 164400
rect 246762 163200 246818 164400
rect 247052 163254 247632 163282
rect 245120 163146 245148 163200
rect 245028 163118 245148 163146
rect 245016 158364 245068 158370
rect 245016 158306 245068 158312
rect 244464 152652 244516 152658
rect 244464 152594 244516 152600
rect 245028 150226 245056 158306
rect 245844 154896 245896 154902
rect 245844 154838 245896 154844
rect 245660 154148 245712 154154
rect 245660 154090 245712 154096
rect 245672 150226 245700 154090
rect 245856 151814 245884 154838
rect 245948 154154 245976 163200
rect 246776 158166 246804 163200
rect 246948 159724 247000 159730
rect 246948 159666 247000 159672
rect 246764 158160 246816 158166
rect 246764 158102 246816 158108
rect 245936 154148 245988 154154
rect 245936 154090 245988 154096
rect 245856 151786 246344 151814
rect 246316 150226 246344 151786
rect 246960 150226 246988 159666
rect 247052 152726 247080 163254
rect 247604 163146 247632 163254
rect 247682 163200 247738 164400
rect 248510 163200 248566 164400
rect 248616 163254 249288 163282
rect 247696 163146 247724 163200
rect 247604 163118 247724 163146
rect 248524 158846 248552 163200
rect 248512 158840 248564 158846
rect 248512 158782 248564 158788
rect 247132 158636 247184 158642
rect 247132 158578 247184 158584
rect 247040 152720 247092 152726
rect 247040 152662 247092 152668
rect 247144 151814 247172 158578
rect 248236 155508 248288 155514
rect 248236 155450 248288 155456
rect 247144 151786 247632 151814
rect 247604 150226 247632 151786
rect 248248 150226 248276 155450
rect 248616 154086 248644 163254
rect 249260 163146 249288 163254
rect 249338 163200 249394 164400
rect 250166 163200 250222 164400
rect 250994 163200 251050 164400
rect 251192 163254 251772 163282
rect 249352 163146 249380 163200
rect 249260 163118 249380 163146
rect 250076 158432 250128 158438
rect 250076 158374 250128 158380
rect 248604 154080 248656 154086
rect 248604 154022 248656 154028
rect 248880 153536 248932 153542
rect 248880 153478 248932 153484
rect 248892 150226 248920 153478
rect 249524 152448 249576 152454
rect 249524 152390 249576 152396
rect 249536 150226 249564 152390
rect 250088 151814 250116 158374
rect 250180 155378 250208 163200
rect 251008 159594 251036 163200
rect 250996 159588 251048 159594
rect 250996 159530 251048 159536
rect 250168 155372 250220 155378
rect 250168 155314 250220 155320
rect 250812 154216 250864 154222
rect 250812 154158 250864 154164
rect 250088 151786 250208 151814
rect 250180 150226 250208 151786
rect 250824 150226 250852 154158
rect 251192 152454 251220 163254
rect 251744 163146 251772 163254
rect 251822 163200 251878 164400
rect 252650 163200 252706 164400
rect 253570 163200 253626 164400
rect 254398 163200 254454 164400
rect 255226 163200 255282 164400
rect 255332 163254 256004 163282
rect 251836 163146 251864 163200
rect 251744 163118 251864 163146
rect 251456 157616 251508 157622
rect 251456 157558 251508 157564
rect 251180 152448 251232 152454
rect 251180 152390 251232 152396
rect 251468 150226 251496 157558
rect 252664 153542 252692 163200
rect 252744 158500 252796 158506
rect 252744 158442 252796 158448
rect 252652 153536 252704 153542
rect 252652 153478 252704 153484
rect 252100 152856 252152 152862
rect 252100 152798 252152 152804
rect 252112 150226 252140 152798
rect 252756 150226 252784 158442
rect 253388 155644 253440 155650
rect 253388 155586 253440 155592
rect 253400 150226 253428 155586
rect 253584 155446 253612 163200
rect 253940 159792 253992 159798
rect 253940 159734 253992 159740
rect 253572 155440 253624 155446
rect 253572 155382 253624 155388
rect 234206 150146 234258 150152
rect 234218 149940 234246 150146
rect 234862 149940 234890 150198
rect 235506 149940 235534 150198
rect 236150 149940 236178 150198
rect 236794 149940 236822 150198
rect 237438 149940 237466 150198
rect 238082 149940 238110 150198
rect 238726 149940 238754 150198
rect 238944 150204 238996 150210
rect 239324 150198 239398 150226
rect 238944 150146 238996 150152
rect 239370 149940 239398 150198
rect 240002 150204 240054 150210
rect 240612 150198 240686 150226
rect 241256 150198 241330 150226
rect 241900 150198 241974 150226
rect 242452 150198 242526 150226
rect 243096 150198 243170 150226
rect 243740 150198 243814 150226
rect 244384 150198 244458 150226
rect 245028 150198 245102 150226
rect 245672 150198 245746 150226
rect 246316 150198 246390 150226
rect 246960 150198 247034 150226
rect 247604 150198 247678 150226
rect 248248 150198 248322 150226
rect 248892 150198 248966 150226
rect 249536 150198 249610 150226
rect 250180 150198 250254 150226
rect 250824 150198 250898 150226
rect 251468 150198 251542 150226
rect 252112 150198 252186 150226
rect 252756 150198 252830 150226
rect 253400 150198 253474 150226
rect 253952 150210 253980 159734
rect 254412 158778 254440 163200
rect 255240 159730 255268 163200
rect 255228 159724 255280 159730
rect 255228 159666 255280 159672
rect 254400 158772 254452 158778
rect 254400 158714 254452 158720
rect 254032 157208 254084 157214
rect 254032 157150 254084 157156
rect 254044 150226 254072 157150
rect 255332 154222 255360 163254
rect 255976 163146 256004 163254
rect 256054 163200 256110 164400
rect 256882 163200 256938 164400
rect 257710 163200 257766 164400
rect 258538 163200 258594 164400
rect 259458 163200 259514 164400
rect 260286 163200 260342 164400
rect 261114 163200 261170 164400
rect 261942 163200 261998 164400
rect 262232 163254 262720 163282
rect 256068 163146 256096 163200
rect 255976 163118 256096 163146
rect 255412 158772 255464 158778
rect 255412 158714 255464 158720
rect 255320 154216 255372 154222
rect 255320 154158 255372 154164
rect 255424 152862 255452 158714
rect 256792 158704 256844 158710
rect 256792 158646 256844 158652
rect 255596 158568 255648 158574
rect 255596 158510 255648 158516
rect 255412 152856 255464 152862
rect 255412 152798 255464 152804
rect 255608 151814 255636 158510
rect 255872 157548 255924 157554
rect 255872 157490 255924 157496
rect 255780 155576 255832 155582
rect 255780 155518 255832 155524
rect 255424 151786 255636 151814
rect 255424 150226 255452 151786
rect 255792 150498 255820 155518
rect 255884 151814 255912 157490
rect 255884 151786 256648 151814
rect 255792 150470 256004 150498
rect 240002 150146 240054 150152
rect 240014 149940 240042 150146
rect 240658 149940 240686 150198
rect 241302 149940 241330 150198
rect 241946 149940 241974 150198
rect 242498 149940 242526 150198
rect 243142 149940 243170 150198
rect 243786 149940 243814 150198
rect 244430 149940 244458 150198
rect 245074 149940 245102 150198
rect 245718 149940 245746 150198
rect 246362 149940 246390 150198
rect 247006 149940 247034 150198
rect 247650 149940 247678 150198
rect 248294 149940 248322 150198
rect 248938 149940 248966 150198
rect 249582 149940 249610 150198
rect 250226 149940 250254 150198
rect 250870 149940 250898 150198
rect 251514 149940 251542 150198
rect 252158 149940 252186 150198
rect 252802 149940 252830 150198
rect 253446 149940 253474 150198
rect 253940 150204 253992 150210
rect 254044 150198 254118 150226
rect 253940 150146 253992 150152
rect 254090 149940 254118 150198
rect 254722 150204 254774 150210
rect 254722 150146 254774 150152
rect 255378 150198 255452 150226
rect 255976 150226 256004 150470
rect 256620 150226 256648 151786
rect 255976 150198 256050 150226
rect 256620 150198 256694 150226
rect 256804 150210 256832 158646
rect 256896 158234 256924 163200
rect 256884 158228 256936 158234
rect 256884 158170 256936 158176
rect 257252 153128 257304 153134
rect 257252 153070 257304 153076
rect 257264 150226 257292 153070
rect 257724 152794 257752 163200
rect 258552 158778 258580 163200
rect 258540 158772 258592 158778
rect 258540 158714 258592 158720
rect 258540 154284 258592 154290
rect 258540 154226 258592 154232
rect 257712 152788 257764 152794
rect 257712 152730 257764 152736
rect 258552 150226 258580 154226
rect 259184 153468 259236 153474
rect 259184 153410 259236 153416
rect 259196 150226 259224 153410
rect 259472 153406 259500 163200
rect 259552 159860 259604 159866
rect 259552 159802 259604 159808
rect 259460 153400 259512 153406
rect 259460 153342 259512 153348
rect 259564 151814 259592 159802
rect 260300 155514 260328 163200
rect 261128 159866 261156 163200
rect 261116 159860 261168 159866
rect 261116 159802 261168 159808
rect 261956 159798 261984 163200
rect 261944 159792 261996 159798
rect 261944 159734 261996 159740
rect 260932 158772 260984 158778
rect 260932 158714 260984 158720
rect 260472 157956 260524 157962
rect 260472 157898 260524 157904
rect 260288 155508 260340 155514
rect 260288 155450 260340 155456
rect 259564 151786 259868 151814
rect 259840 150226 259868 151786
rect 260484 150226 260512 157898
rect 260840 155712 260892 155718
rect 260840 155654 260892 155660
rect 260852 151814 260880 155654
rect 260944 151910 260972 158714
rect 261392 154964 261444 154970
rect 261392 154906 261444 154912
rect 260932 151904 260984 151910
rect 260932 151846 260984 151852
rect 261404 151814 261432 154906
rect 262232 154290 262260 163254
rect 262692 163146 262720 163254
rect 262770 163200 262826 164400
rect 263598 163200 263654 164400
rect 264426 163200 264482 164400
rect 264992 163254 265296 163282
rect 262784 163146 262812 163200
rect 262692 163118 262812 163146
rect 263048 157888 263100 157894
rect 263048 157830 263100 157836
rect 262220 154284 262272 154290
rect 262220 154226 262272 154232
rect 262404 152312 262456 152318
rect 262404 152254 262456 152260
rect 260852 151786 261156 151814
rect 261404 151786 261800 151814
rect 261128 150226 261156 151786
rect 261772 150226 261800 151786
rect 262416 150226 262444 152254
rect 263060 150226 263088 157830
rect 263612 155582 263640 163200
rect 264440 158778 264468 163200
rect 264888 159928 264940 159934
rect 264888 159870 264940 159876
rect 264428 158772 264480 158778
rect 264428 158714 264480 158720
rect 263692 157752 263744 157758
rect 263692 157694 263744 157700
rect 263600 155576 263652 155582
rect 263600 155518 263652 155524
rect 263704 150346 263732 157694
rect 263784 155848 263836 155854
rect 263784 155790 263836 155796
rect 263692 150340 263744 150346
rect 263692 150282 263744 150288
rect 263796 150226 263824 155790
rect 264900 151814 264928 159870
rect 264992 153134 265020 163254
rect 265268 163146 265296 163254
rect 265346 163200 265402 164400
rect 265452 163254 266124 163282
rect 265360 163146 265388 163200
rect 265268 163118 265388 163146
rect 265164 157276 265216 157282
rect 265164 157218 265216 157224
rect 264980 153128 265032 153134
rect 264980 153070 265032 153076
rect 265176 151814 265204 157218
rect 265452 153474 265480 163254
rect 266096 163146 266124 163254
rect 266174 163200 266230 164400
rect 267002 163200 267058 164400
rect 267830 163200 267886 164400
rect 268658 163200 268714 164400
rect 269224 163254 269436 163282
rect 266188 163146 266216 163200
rect 266096 163118 266216 163146
rect 266360 158772 266412 158778
rect 266360 158714 266412 158720
rect 266268 155916 266320 155922
rect 266268 155858 266320 155864
rect 265440 153468 265492 153474
rect 265440 153410 265492 153416
rect 264900 151786 265020 151814
rect 265176 151786 265664 151814
rect 254734 149940 254762 150146
rect 255378 149940 255406 150198
rect 256022 149940 256050 150198
rect 256666 149940 256694 150198
rect 256792 150204 256844 150210
rect 257264 150198 257338 150226
rect 256792 150146 256844 150152
rect 257310 149940 257338 150198
rect 257942 150204 257994 150210
rect 258552 150198 258626 150226
rect 259196 150198 259270 150226
rect 259840 150198 259914 150226
rect 260484 150198 260558 150226
rect 261128 150198 261202 150226
rect 261772 150198 261846 150226
rect 262416 150198 262490 150226
rect 263060 150198 263134 150226
rect 257942 150146 257994 150152
rect 257954 149940 257982 150146
rect 258598 149940 258626 150198
rect 259242 149940 259270 150198
rect 259886 149940 259914 150198
rect 260530 149940 260558 150198
rect 261174 149940 261202 150198
rect 261818 149940 261846 150198
rect 262462 149940 262490 150198
rect 263106 149940 263134 150198
rect 263750 150198 263824 150226
rect 264992 150226 265020 151786
rect 265636 150226 265664 151786
rect 266280 150226 266308 155858
rect 266372 152318 266400 158714
rect 266912 156324 266964 156330
rect 266912 156266 266964 156272
rect 266360 152312 266412 152318
rect 266360 152254 266412 152260
rect 266924 150226 266952 156266
rect 267016 155650 267044 163200
rect 267844 158778 267872 163200
rect 268672 159934 268700 163200
rect 269120 159996 269172 160002
rect 269120 159938 269172 159944
rect 268660 159928 268712 159934
rect 268660 159870 268712 159876
rect 267832 158772 267884 158778
rect 267832 158714 267884 158720
rect 267740 157820 267792 157826
rect 267740 157762 267792 157768
rect 267004 155644 267056 155650
rect 267004 155586 267056 155592
rect 267556 153060 267608 153066
rect 267556 153002 267608 153008
rect 267568 150226 267596 153002
rect 267752 151814 267780 157762
rect 268844 155168 268896 155174
rect 268844 155110 268896 155116
rect 267752 151786 268240 151814
rect 268212 150226 268240 151786
rect 268856 150226 268884 155110
rect 264382 150204 264434 150210
rect 263750 149940 263778 150198
rect 264992 150198 265066 150226
rect 265636 150198 265710 150226
rect 266280 150198 266354 150226
rect 266924 150198 266998 150226
rect 267568 150198 267642 150226
rect 268212 150198 268286 150226
rect 268856 150198 268930 150226
rect 269132 150210 269160 159938
rect 269224 153338 269252 163254
rect 269408 163146 269436 163254
rect 269486 163200 269542 164400
rect 270314 163200 270370 164400
rect 271234 163200 271290 164400
rect 272062 163200 272118 164400
rect 272890 163200 272946 164400
rect 273718 163200 273774 164400
rect 274546 163200 274602 164400
rect 275374 163200 275430 164400
rect 276202 163200 276258 164400
rect 277122 163200 277178 164400
rect 277412 163254 277900 163282
rect 269500 163146 269528 163200
rect 269408 163118 269528 163146
rect 270328 155718 270356 163200
rect 271248 160002 271276 163200
rect 272076 161474 272104 163200
rect 272076 161446 272196 161474
rect 271236 159996 271288 160002
rect 271236 159938 271288 159944
rect 272064 157004 272116 157010
rect 272064 156946 272116 156952
rect 270500 156052 270552 156058
rect 270500 155994 270552 156000
rect 270316 155712 270368 155718
rect 270316 155654 270368 155660
rect 269488 155032 269540 155038
rect 269488 154974 269540 154980
rect 269212 153332 269264 153338
rect 269212 153274 269264 153280
rect 269500 150226 269528 154974
rect 270512 151814 270540 155994
rect 271420 155100 271472 155106
rect 271420 155042 271472 155048
rect 270512 151786 270816 151814
rect 270788 150226 270816 151786
rect 271432 150226 271460 155042
rect 272076 150226 272104 156946
rect 272168 153066 272196 161446
rect 272800 159996 272852 160002
rect 272800 159938 272852 159944
rect 272156 153060 272208 153066
rect 272156 153002 272208 153008
rect 272812 151978 272840 159938
rect 272904 153270 272932 163200
rect 273732 157078 273760 163200
rect 274560 159497 274588 163200
rect 275388 160002 275416 163200
rect 275376 159996 275428 160002
rect 275376 159938 275428 159944
rect 274546 159488 274602 159497
rect 274546 159423 274602 159432
rect 275190 159352 275246 159361
rect 275190 159287 275246 159296
rect 273720 157072 273772 157078
rect 273720 157014 273772 157020
rect 273904 156188 273956 156194
rect 273904 156130 273956 156136
rect 273260 156120 273312 156126
rect 273260 156062 273312 156068
rect 272892 153264 272944 153270
rect 272892 153206 272944 153212
rect 272708 151972 272760 151978
rect 272708 151914 272760 151920
rect 272800 151972 272852 151978
rect 272800 151914 272852 151920
rect 272720 150226 272748 151914
rect 273272 150226 273300 156062
rect 273916 150226 273944 156130
rect 274548 152176 274600 152182
rect 274548 152118 274600 152124
rect 274560 150226 274588 152118
rect 275204 150226 275232 159287
rect 276112 155780 276164 155786
rect 276112 155722 276164 155728
rect 275836 154420 275888 154426
rect 275836 154362 275888 154368
rect 275848 150226 275876 154362
rect 276124 151814 276152 155722
rect 276216 154426 276244 163200
rect 277136 157010 277164 163200
rect 277124 157004 277176 157010
rect 277124 156946 277176 156952
rect 277124 156256 277176 156262
rect 277124 156198 277176 156204
rect 276204 154420 276256 154426
rect 276204 154362 276256 154368
rect 276124 151786 276520 151814
rect 276492 150226 276520 151786
rect 277136 150226 277164 156198
rect 277412 152182 277440 163254
rect 277872 163146 277900 163254
rect 277950 163200 278006 164400
rect 278778 163200 278834 164400
rect 278884 163254 279556 163282
rect 277964 163146 277992 163200
rect 277872 163118 277992 163146
rect 278412 154352 278464 154358
rect 278412 154294 278464 154300
rect 277768 152924 277820 152930
rect 277768 152866 277820 152872
rect 277400 152176 277452 152182
rect 277400 152118 277452 152124
rect 277780 150226 277808 152866
rect 278424 150226 278452 154294
rect 278792 152930 278820 163200
rect 278884 154358 278912 163254
rect 279528 163146 279556 163254
rect 279606 163200 279662 164400
rect 280434 163200 280490 164400
rect 281262 163200 281318 164400
rect 282090 163200 282146 164400
rect 283010 163200 283066 164400
rect 283116 163254 283328 163282
rect 279620 163146 279648 163200
rect 279528 163118 279648 163146
rect 280344 160064 280396 160070
rect 280344 160006 280396 160012
rect 279056 156392 279108 156398
rect 279056 156334 279108 156340
rect 278872 154352 278924 154358
rect 278872 154294 278924 154300
rect 278780 152924 278832 152930
rect 278780 152866 278832 152872
rect 279068 150226 279096 156334
rect 279700 153196 279752 153202
rect 279700 153138 279752 153144
rect 279712 150226 279740 153138
rect 280356 150226 280384 160006
rect 280448 157146 280476 163200
rect 281276 160070 281304 163200
rect 281264 160064 281316 160070
rect 281264 160006 281316 160012
rect 282104 159322 282132 163200
rect 283024 163146 283052 163200
rect 283116 163146 283144 163254
rect 283024 163118 283144 163146
rect 281540 159316 281592 159322
rect 281540 159258 281592 159264
rect 282092 159316 282144 159322
rect 282092 159258 282144 159264
rect 280436 157140 280488 157146
rect 280436 157082 280488 157088
rect 280986 153776 281042 153785
rect 280986 153711 281042 153720
rect 281000 150226 281028 153711
rect 264382 150146 264434 150152
rect 264394 149940 264422 150146
rect 265038 149940 265066 150198
rect 265682 149940 265710 150198
rect 266326 149940 266354 150198
rect 266970 149940 266998 150198
rect 267614 149940 267642 150198
rect 268258 149940 268286 150198
rect 268902 149940 268930 150198
rect 269120 150204 269172 150210
rect 269500 150198 269574 150226
rect 269120 150146 269172 150152
rect 269546 149940 269574 150198
rect 270178 150204 270230 150210
rect 270788 150198 270862 150226
rect 271432 150198 271506 150226
rect 272076 150198 272150 150226
rect 272720 150198 272794 150226
rect 273272 150198 273346 150226
rect 273916 150198 273990 150226
rect 274560 150198 274634 150226
rect 275204 150198 275278 150226
rect 275848 150198 275922 150226
rect 276492 150198 276566 150226
rect 277136 150198 277210 150226
rect 277780 150198 277854 150226
rect 278424 150198 278498 150226
rect 279068 150198 279142 150226
rect 279712 150198 279786 150226
rect 280356 150198 280430 150226
rect 281000 150198 281074 150226
rect 281552 150210 281580 159258
rect 283196 159180 283248 159186
rect 283196 159122 283248 159128
rect 283104 156664 283156 156670
rect 283104 156606 283156 156612
rect 281632 156596 281684 156602
rect 281632 156538 281684 156544
rect 281644 150226 281672 156538
rect 282920 152244 282972 152250
rect 282920 152186 282972 152192
rect 282932 150226 282960 152186
rect 270178 150146 270230 150152
rect 270190 149940 270218 150146
rect 270834 149940 270862 150198
rect 271478 149940 271506 150198
rect 272122 149940 272150 150198
rect 272766 149940 272794 150198
rect 273318 149940 273346 150198
rect 273962 149940 273990 150198
rect 274606 149940 274634 150198
rect 275250 149940 275278 150198
rect 275894 149940 275922 150198
rect 276538 149940 276566 150198
rect 277182 149940 277210 150198
rect 277826 149940 277854 150198
rect 278470 149940 278498 150198
rect 279114 149940 279142 150198
rect 279758 149940 279786 150198
rect 280402 149940 280430 150198
rect 281046 149940 281074 150198
rect 281540 150204 281592 150210
rect 281644 150198 281718 150226
rect 281540 150146 281592 150152
rect 281690 149940 281718 150198
rect 282322 150204 282374 150210
rect 282932 150198 283006 150226
rect 283116 150210 283144 156606
rect 283208 151842 283236 159122
rect 283300 154494 283328 163254
rect 283838 163200 283894 164400
rect 284666 163200 284722 164400
rect 285494 163200 285550 164400
rect 285692 163254 286272 163282
rect 283852 157282 283880 163200
rect 284392 159248 284444 159254
rect 284392 159190 284444 159196
rect 283840 157276 283892 157282
rect 283840 157218 283892 157224
rect 283656 154556 283708 154562
rect 283656 154498 283708 154504
rect 283288 154488 283340 154494
rect 283288 154430 283340 154436
rect 283196 151836 283248 151842
rect 283196 151778 283248 151784
rect 283668 150226 283696 154498
rect 282322 150146 282374 150152
rect 282334 149940 282362 150146
rect 282978 149940 283006 150198
rect 283104 150204 283156 150210
rect 283104 150146 283156 150152
rect 283622 150198 283696 150226
rect 284404 150210 284432 159190
rect 284680 159186 284708 163200
rect 284668 159180 284720 159186
rect 284668 159122 284720 159128
rect 285508 153202 285536 163200
rect 285692 154562 285720 163254
rect 286244 163146 286272 163254
rect 286322 163200 286378 164400
rect 287150 163200 287206 164400
rect 287978 163200 288034 164400
rect 288898 163200 288954 164400
rect 289726 163200 289782 164400
rect 290554 163200 290610 164400
rect 291382 163200 291438 164400
rect 292210 163200 292266 164400
rect 293038 163200 293094 164400
rect 293866 163200 293922 164400
rect 294786 163200 294842 164400
rect 295614 163200 295670 164400
rect 296442 163200 296498 164400
rect 297270 163200 297326 164400
rect 298098 163200 298154 164400
rect 298664 163254 298876 163282
rect 286336 163146 286364 163200
rect 286244 163118 286364 163146
rect 285772 159180 285824 159186
rect 285772 159122 285824 159128
rect 285588 154556 285640 154562
rect 285588 154498 285640 154504
rect 285680 154556 285732 154562
rect 285680 154498 285732 154504
rect 285600 154442 285628 154498
rect 285600 154414 285720 154442
rect 285496 153196 285548 153202
rect 285496 153138 285548 153144
rect 284852 152992 284904 152998
rect 284852 152934 284904 152940
rect 284864 150226 284892 152934
rect 285692 151814 285720 154414
rect 285784 152250 285812 159122
rect 287164 156738 287192 163200
rect 287992 159254 288020 163200
rect 287980 159248 288032 159254
rect 287980 159190 288032 159196
rect 288912 159186 288940 163200
rect 288164 159180 288216 159186
rect 288164 159122 288216 159128
rect 288900 159180 288952 159186
rect 288900 159122 288952 159128
rect 286232 156732 286284 156738
rect 286232 156674 286284 156680
rect 287152 156732 287204 156738
rect 287152 156674 287204 156680
rect 285772 152244 285824 152250
rect 285772 152186 285824 152192
rect 286244 151814 286272 156674
rect 288176 152998 288204 159122
rect 289360 156868 289412 156874
rect 289360 156810 289412 156816
rect 288716 154012 288768 154018
rect 288716 153954 288768 153960
rect 288164 152992 288216 152998
rect 288164 152934 288216 152940
rect 288072 152380 288124 152386
rect 288072 152322 288124 152328
rect 287428 151836 287480 151842
rect 285692 151786 286180 151814
rect 286244 151786 286824 151814
rect 286152 150226 286180 151786
rect 286796 150226 286824 151786
rect 287428 151778 287480 151784
rect 287440 150226 287468 151778
rect 288084 150226 288112 152322
rect 288728 150226 288756 153954
rect 289372 150226 289400 156810
rect 289740 155786 289768 163200
rect 290568 156874 290596 163200
rect 290648 159384 290700 159390
rect 290648 159326 290700 159332
rect 290556 156868 290608 156874
rect 290556 156810 290608 156816
rect 289728 155780 289780 155786
rect 289728 155722 289780 155728
rect 290004 152992 290056 152998
rect 290004 152934 290056 152940
rect 290016 150226 290044 152934
rect 290660 150226 290688 159326
rect 291292 153944 291344 153950
rect 291292 153886 291344 153892
rect 291304 150226 291332 153886
rect 291396 152998 291424 163200
rect 291936 156936 291988 156942
rect 291936 156878 291988 156884
rect 291384 152992 291436 152998
rect 291384 152934 291436 152940
rect 291948 150226 291976 156878
rect 292224 152386 292252 163200
rect 293052 155854 293080 163200
rect 293880 156942 293908 163200
rect 294800 159390 294828 163200
rect 295628 159526 295656 163200
rect 295524 159520 295576 159526
rect 295524 159462 295576 159468
rect 295616 159520 295668 159526
rect 295616 159462 295668 159468
rect 294788 159384 294840 159390
rect 294788 159326 294840 159332
rect 295156 159044 295208 159050
rect 295156 158986 295208 158992
rect 293868 156936 293920 156942
rect 293868 156878 293920 156884
rect 294052 156800 294104 156806
rect 294052 156742 294104 156748
rect 293040 155848 293092 155854
rect 293040 155790 293092 155796
rect 293868 153740 293920 153746
rect 293868 153682 293920 153688
rect 293224 152516 293276 152522
rect 293224 152458 293276 152464
rect 292578 152416 292634 152425
rect 292212 152380 292264 152386
rect 292578 152351 292634 152360
rect 292212 152322 292264 152328
rect 292592 150226 292620 152351
rect 293236 150226 293264 152458
rect 293880 150226 293908 153682
rect 294064 151814 294092 156742
rect 294064 151786 294552 151814
rect 294524 150226 294552 151786
rect 295168 150226 295196 158986
rect 295536 151814 295564 159462
rect 296456 155922 296484 163200
rect 297284 156806 297312 163200
rect 298008 159452 298060 159458
rect 298008 159394 298060 159400
rect 297272 156800 297324 156806
rect 297272 156742 297324 156748
rect 296444 155916 296496 155922
rect 296444 155858 296496 155864
rect 297088 155236 297140 155242
rect 297088 155178 297140 155184
rect 296444 153808 296496 153814
rect 296444 153750 296496 153756
rect 295536 151786 295840 151814
rect 295812 150226 295840 151786
rect 296456 150226 296484 153750
rect 297100 150226 297128 155178
rect 297732 152584 297784 152590
rect 297732 152526 297784 152532
rect 297744 150226 297772 152526
rect 298020 151814 298048 159394
rect 298112 159050 298140 163200
rect 298100 159044 298152 159050
rect 298100 158986 298152 158992
rect 298664 152522 298692 163254
rect 298848 163146 298876 163254
rect 298926 163200 298982 164400
rect 299754 163200 299810 164400
rect 300674 163200 300730 164400
rect 301502 163200 301558 164400
rect 302330 163200 302386 164400
rect 303158 163200 303214 164400
rect 303724 163254 303936 163282
rect 298940 163146 298968 163200
rect 298848 163118 298968 163146
rect 299572 159044 299624 159050
rect 299572 158986 299624 158992
rect 299480 158976 299532 158982
rect 299480 158918 299532 158924
rect 299020 153672 299072 153678
rect 299020 153614 299072 153620
rect 298652 152516 298704 152522
rect 298652 152458 298704 152464
rect 298020 151786 298416 151814
rect 298388 150226 298416 151786
rect 299032 150226 299060 153614
rect 284254 150204 284306 150210
rect 283622 149940 283650 150198
rect 284254 150146 284306 150152
rect 284392 150204 284444 150210
rect 284864 150198 284938 150226
rect 284392 150146 284444 150152
rect 284266 149940 284294 150146
rect 284910 149940 284938 150198
rect 285542 150204 285594 150210
rect 286152 150198 286226 150226
rect 286796 150198 286870 150226
rect 287440 150198 287514 150226
rect 288084 150198 288158 150226
rect 288728 150198 288802 150226
rect 289372 150198 289446 150226
rect 290016 150198 290090 150226
rect 290660 150198 290734 150226
rect 291304 150198 291378 150226
rect 291948 150198 292022 150226
rect 292592 150198 292666 150226
rect 293236 150198 293310 150226
rect 293880 150198 293954 150226
rect 294524 150198 294598 150226
rect 295168 150198 295242 150226
rect 295812 150198 295886 150226
rect 296456 150198 296530 150226
rect 297100 150198 297174 150226
rect 297744 150198 297818 150226
rect 298388 150198 298462 150226
rect 299032 150198 299106 150226
rect 299492 150210 299520 158918
rect 299584 151842 299612 158986
rect 299664 158024 299716 158030
rect 299664 157966 299716 157972
rect 299572 151836 299624 151842
rect 299572 151778 299624 151784
rect 299676 150226 299704 157966
rect 299768 155242 299796 163200
rect 300688 157214 300716 163200
rect 301516 159458 301544 163200
rect 302344 159662 302372 163200
rect 302240 159656 302292 159662
rect 302240 159598 302292 159604
rect 302332 159656 302384 159662
rect 302332 159598 302384 159604
rect 301504 159452 301556 159458
rect 301504 159394 301556 159400
rect 302252 159118 302280 159598
rect 302240 159112 302292 159118
rect 302240 159054 302292 159060
rect 300676 157208 300728 157214
rect 300676 157150 300728 157156
rect 302332 155304 302384 155310
rect 302332 155246 302384 155252
rect 299756 155236 299808 155242
rect 299756 155178 299808 155184
rect 301596 153604 301648 153610
rect 301596 153546 301648 153552
rect 300952 152040 301004 152046
rect 300952 151982 301004 151988
rect 300964 150226 300992 151982
rect 301608 150226 301636 153546
rect 302344 150226 302372 155246
rect 303172 155174 303200 163200
rect 303528 159112 303580 159118
rect 303528 159054 303580 159060
rect 303160 155168 303212 155174
rect 303160 155110 303212 155116
rect 302884 152108 302936 152114
rect 302884 152050 302936 152056
rect 285542 150146 285594 150152
rect 285554 149940 285582 150146
rect 286198 149940 286226 150198
rect 286842 149940 286870 150198
rect 287486 149940 287514 150198
rect 288130 149940 288158 150198
rect 288774 149940 288802 150198
rect 289418 149940 289446 150198
rect 290062 149940 290090 150198
rect 290706 149940 290734 150198
rect 291350 149940 291378 150198
rect 291994 149940 292022 150198
rect 292638 149940 292666 150198
rect 293282 149940 293310 150198
rect 293926 149940 293954 150198
rect 294570 149940 294598 150198
rect 295214 149940 295242 150198
rect 295858 149940 295886 150198
rect 296502 149940 296530 150198
rect 297146 149940 297174 150198
rect 297790 149940 297818 150198
rect 298434 149940 298462 150198
rect 299078 149940 299106 150198
rect 299480 150204 299532 150210
rect 299676 150198 299750 150226
rect 299480 150146 299532 150152
rect 299722 149940 299750 150198
rect 300354 150204 300406 150210
rect 300964 150198 301038 150226
rect 301608 150198 301682 150226
rect 300354 150146 300406 150152
rect 300366 149940 300394 150146
rect 301010 149940 301038 150198
rect 301654 149940 301682 150198
rect 302298 150198 302372 150226
rect 302896 150226 302924 152050
rect 303540 150226 303568 159054
rect 303724 152114 303752 163254
rect 303908 163146 303936 163254
rect 303986 163200 304042 164400
rect 304814 163200 304870 164400
rect 305642 163200 305698 164400
rect 306562 163200 306618 164400
rect 307390 163200 307446 164400
rect 308218 163200 308274 164400
rect 309046 163200 309102 164400
rect 309152 163254 309824 163282
rect 304000 163146 304028 163200
rect 303908 163118 304028 163146
rect 304724 158092 304776 158098
rect 304724 158034 304776 158040
rect 304080 153876 304132 153882
rect 304080 153818 304132 153824
rect 303712 152108 303764 152114
rect 303712 152050 303764 152056
rect 304092 150226 304120 153818
rect 304736 150226 304764 158034
rect 304828 152590 304856 163200
rect 305368 159044 305420 159050
rect 305368 158986 305420 158992
rect 304816 152584 304868 152590
rect 304816 152526 304868 152532
rect 305380 150226 305408 158986
rect 305656 158914 305684 163200
rect 305644 158908 305696 158914
rect 305644 158850 305696 158856
rect 306576 155310 306604 163200
rect 307404 159050 307432 163200
rect 307392 159044 307444 159050
rect 307392 158986 307444 158992
rect 308232 158982 308260 163200
rect 309060 159118 309088 163200
rect 309048 159112 309100 159118
rect 309048 159054 309100 159060
rect 308220 158976 308272 158982
rect 308220 158918 308272 158924
rect 307392 158908 307444 158914
rect 307392 158850 307444 158856
rect 308588 158908 308640 158914
rect 308588 158850 308640 158856
rect 306932 158160 306984 158166
rect 306932 158102 306984 158108
rect 306564 155304 306616 155310
rect 306564 155246 306616 155252
rect 306656 154148 306708 154154
rect 306656 154090 306708 154096
rect 306012 152652 306064 152658
rect 306012 152594 306064 152600
rect 306024 150226 306052 152594
rect 306668 150226 306696 154090
rect 306944 151814 306972 158102
rect 307404 152046 307432 158850
rect 307944 152720 307996 152726
rect 307944 152662 307996 152668
rect 307392 152040 307444 152046
rect 307392 151982 307444 151988
rect 306944 151786 307340 151814
rect 307312 150226 307340 151786
rect 307956 150226 307984 152662
rect 308600 150226 308628 158850
rect 309152 153882 309180 163254
rect 309796 163146 309824 163254
rect 309874 163200 309930 164400
rect 310702 163200 310758 164400
rect 311530 163200 311586 164400
rect 312450 163200 312506 164400
rect 313278 163200 313334 164400
rect 314106 163200 314162 164400
rect 314934 163200 314990 164400
rect 315762 163200 315818 164400
rect 316052 163254 316540 163282
rect 309888 163146 309916 163200
rect 309796 163118 309916 163146
rect 310612 159588 310664 159594
rect 310612 159530 310664 159536
rect 309876 155372 309928 155378
rect 309876 155314 309928 155320
rect 309232 154080 309284 154086
rect 309232 154022 309284 154028
rect 309140 153876 309192 153882
rect 309140 153818 309192 153824
rect 309244 150226 309272 154022
rect 309888 150226 309916 155314
rect 310624 150226 310652 159530
rect 310716 158846 310744 163200
rect 310704 158840 310756 158846
rect 310704 158782 310756 158788
rect 311544 152658 311572 163200
rect 312464 158914 312492 163200
rect 312452 158908 312504 158914
rect 312452 158850 312504 158856
rect 313188 158840 313240 158846
rect 313188 158782 313240 158788
rect 312452 155440 312504 155446
rect 312452 155382 312504 155388
rect 311808 153536 311860 153542
rect 311808 153478 311860 153484
rect 311532 152652 311584 152658
rect 311532 152594 311584 152600
rect 311164 152448 311216 152454
rect 311164 152390 311216 152396
rect 302896 150198 302970 150226
rect 303540 150198 303614 150226
rect 304092 150198 304166 150226
rect 304736 150198 304810 150226
rect 305380 150198 305454 150226
rect 306024 150198 306098 150226
rect 306668 150198 306742 150226
rect 307312 150198 307386 150226
rect 307956 150198 308030 150226
rect 308600 150198 308674 150226
rect 309244 150198 309318 150226
rect 309888 150198 309962 150226
rect 302298 149940 302326 150198
rect 302942 149940 302970 150198
rect 303586 149940 303614 150198
rect 304138 149940 304166 150198
rect 304782 149940 304810 150198
rect 305426 149940 305454 150198
rect 306070 149940 306098 150198
rect 306714 149940 306742 150198
rect 307358 149940 307386 150198
rect 308002 149940 308030 150198
rect 308646 149940 308674 150198
rect 309290 149940 309318 150198
rect 309934 149940 309962 150198
rect 310578 150198 310652 150226
rect 311176 150226 311204 152390
rect 311820 150226 311848 153478
rect 312464 150226 312492 155382
rect 313200 152862 313228 158782
rect 313292 154018 313320 163200
rect 314120 159730 314148 163200
rect 313372 159724 313424 159730
rect 313372 159666 313424 159672
rect 314108 159724 314160 159730
rect 314108 159666 314160 159672
rect 313280 154012 313332 154018
rect 313280 153954 313332 153960
rect 313096 152856 313148 152862
rect 313096 152798 313148 152804
rect 313188 152856 313240 152862
rect 313188 152798 313240 152804
rect 313108 150226 313136 152798
rect 313384 151814 313412 159666
rect 314948 158914 314976 163200
rect 315776 159594 315804 163200
rect 315764 159588 315816 159594
rect 315764 159530 315816 159536
rect 313648 158908 313700 158914
rect 313648 158850 313700 158856
rect 314936 158908 314988 158914
rect 314936 158850 314988 158856
rect 313660 152425 313688 158850
rect 315028 158228 315080 158234
rect 315028 158170 315080 158176
rect 314384 154216 314436 154222
rect 314384 154158 314436 154164
rect 313646 152416 313702 152425
rect 313646 152351 313702 152360
rect 313384 151786 313780 151814
rect 313752 150226 313780 151786
rect 314396 150226 314424 154158
rect 315040 150226 315068 158170
rect 316052 153950 316080 163254
rect 316512 163146 316540 163254
rect 316590 163200 316646 164400
rect 317418 163200 317474 164400
rect 318338 163200 318394 164400
rect 319166 163200 319222 164400
rect 319994 163200 320050 164400
rect 320822 163200 320878 164400
rect 321650 163200 321706 164400
rect 322478 163200 322534 164400
rect 323306 163200 323362 164400
rect 324226 163200 324282 164400
rect 324332 163254 325004 163282
rect 316604 163146 316632 163200
rect 316512 163118 316632 163146
rect 317052 159860 317104 159866
rect 317052 159802 317104 159808
rect 316040 153944 316092 153950
rect 316040 153886 316092 153892
rect 316960 153400 317012 153406
rect 316960 153342 317012 153348
rect 315672 152788 315724 152794
rect 315672 152730 315724 152736
rect 315684 150226 315712 152730
rect 316316 151904 316368 151910
rect 316316 151846 316368 151852
rect 316328 150226 316356 151846
rect 316972 150226 317000 153342
rect 317064 152794 317092 159802
rect 317052 152788 317104 152794
rect 317052 152730 317104 152736
rect 317432 152454 317460 163200
rect 317604 155508 317656 155514
rect 317604 155450 317656 155456
rect 317420 152448 317472 152454
rect 317420 152390 317472 152396
rect 317616 150226 317644 155450
rect 318248 152788 318300 152794
rect 318248 152730 318300 152736
rect 318260 150226 318288 152730
rect 318352 152726 318380 163200
rect 318892 159792 318944 159798
rect 318892 159734 318944 159740
rect 318340 152720 318392 152726
rect 318340 152662 318392 152668
rect 318904 150226 318932 159734
rect 319180 158846 319208 163200
rect 319168 158840 319220 158846
rect 319168 158782 319220 158788
rect 320008 155378 320036 163200
rect 320836 159866 320864 163200
rect 320824 159860 320876 159866
rect 320824 159802 320876 159808
rect 321664 158846 321692 163200
rect 322492 159798 322520 163200
rect 322480 159792 322532 159798
rect 322480 159734 322532 159740
rect 321560 158840 321612 158846
rect 321560 158782 321612 158788
rect 321652 158840 321704 158846
rect 321652 158782 321704 158788
rect 320272 158772 320324 158778
rect 320272 158714 320324 158720
rect 320180 155576 320232 155582
rect 320180 155518 320232 155524
rect 319996 155372 320048 155378
rect 319996 155314 320048 155320
rect 319536 154284 319588 154290
rect 319536 154226 319588 154232
rect 319548 150226 319576 154226
rect 320192 150226 320220 155518
rect 320284 152794 320312 158714
rect 321468 153128 321520 153134
rect 321468 153070 321520 153076
rect 320272 152788 320324 152794
rect 320272 152730 320324 152736
rect 320824 152312 320876 152318
rect 320824 152254 320876 152260
rect 320836 150226 320864 152254
rect 321480 150226 321508 153070
rect 321572 151910 321600 158782
rect 321744 155644 321796 155650
rect 321744 155586 321796 155592
rect 321560 151904 321612 151910
rect 321560 151846 321612 151852
rect 311176 150198 311250 150226
rect 311820 150198 311894 150226
rect 312464 150198 312538 150226
rect 313108 150198 313182 150226
rect 313752 150198 313826 150226
rect 314396 150198 314470 150226
rect 315040 150198 315114 150226
rect 315684 150198 315758 150226
rect 316328 150198 316402 150226
rect 316972 150198 317046 150226
rect 317616 150198 317690 150226
rect 318260 150198 318334 150226
rect 318904 150198 318978 150226
rect 319548 150198 319622 150226
rect 320192 150198 320266 150226
rect 320836 150198 320910 150226
rect 321480 150198 321554 150226
rect 321756 150210 321784 155586
rect 323320 154086 323348 163200
rect 324044 159928 324096 159934
rect 324044 159870 324096 159876
rect 323308 154080 323360 154086
rect 323308 154022 323360 154028
rect 322204 153468 322256 153474
rect 322204 153410 322256 153416
rect 322216 150226 322244 153410
rect 323124 152788 323176 152794
rect 323124 152730 323176 152736
rect 323136 151814 323164 152730
rect 323136 151786 323440 151814
rect 310578 149940 310606 150198
rect 311222 149940 311250 150198
rect 311866 149940 311894 150198
rect 312510 149940 312538 150198
rect 313154 149940 313182 150198
rect 313798 149940 313826 150198
rect 314442 149940 314470 150198
rect 315086 149940 315114 150198
rect 315730 149940 315758 150198
rect 316374 149940 316402 150198
rect 317018 149940 317046 150198
rect 317662 149940 317690 150198
rect 318306 149940 318334 150198
rect 318950 149940 318978 150198
rect 319594 149940 319622 150198
rect 320238 149940 320266 150198
rect 320882 149940 320910 150198
rect 321526 149940 321554 150198
rect 321744 150204 321796 150210
rect 321744 150146 321796 150152
rect 322170 150198 322244 150226
rect 323412 150226 323440 151786
rect 324056 150226 324084 159870
rect 324240 152794 324268 163200
rect 324332 153134 324360 163254
rect 324976 163146 325004 163254
rect 325054 163200 325110 164400
rect 325882 163200 325938 164400
rect 326710 163200 326766 164400
rect 327538 163200 327594 164400
rect 328366 163200 328422 164400
rect 329194 163200 329250 164400
rect 330114 163200 330170 164400
rect 330942 163200 330998 164400
rect 331232 163254 331720 163282
rect 325068 163146 325096 163200
rect 324976 163118 325096 163146
rect 325332 155712 325384 155718
rect 325332 155654 325384 155660
rect 324688 153332 324740 153338
rect 324688 153274 324740 153280
rect 324320 153128 324372 153134
rect 324320 153070 324372 153076
rect 324228 152788 324280 152794
rect 324228 152730 324280 152736
rect 324700 150226 324728 153274
rect 325344 150226 325372 155654
rect 325896 152318 325924 163200
rect 326724 154154 326752 163200
rect 327552 158778 327580 163200
rect 328380 159934 328408 163200
rect 329208 160002 329236 163200
rect 328460 159996 328512 160002
rect 328460 159938 328512 159944
rect 329196 159996 329248 160002
rect 329196 159938 329248 159944
rect 328368 159928 328420 159934
rect 328368 159870 328420 159876
rect 327540 158772 327592 158778
rect 327540 158714 327592 158720
rect 327908 157072 327960 157078
rect 327908 157014 327960 157020
rect 326712 154148 326764 154154
rect 326712 154090 326764 154096
rect 327264 153264 327316 153270
rect 327264 153206 327316 153212
rect 326620 153060 326672 153066
rect 326620 153002 326672 153008
rect 325884 152312 325936 152318
rect 325884 152254 325936 152260
rect 325976 151972 326028 151978
rect 325976 151914 326028 151920
rect 325988 150226 326016 151914
rect 326632 150226 326660 153002
rect 327276 150226 327304 153206
rect 327920 150226 327948 157014
rect 322802 150204 322854 150210
rect 322170 149940 322198 150198
rect 323412 150198 323486 150226
rect 324056 150198 324130 150226
rect 324700 150198 324774 150226
rect 325344 150198 325418 150226
rect 325988 150198 326062 150226
rect 326632 150198 326706 150226
rect 327276 150198 327350 150226
rect 327920 150198 327994 150226
rect 328472 150210 328500 159938
rect 328550 159488 328606 159497
rect 328550 159423 328606 159432
rect 328564 150226 328592 159423
rect 330128 155446 330156 163200
rect 330484 157004 330536 157010
rect 330484 156946 330536 156952
rect 330116 155440 330168 155446
rect 330116 155382 330168 155388
rect 329932 154420 329984 154426
rect 329932 154362 329984 154368
rect 329944 150226 329972 154362
rect 322802 150146 322854 150152
rect 322814 149940 322842 150146
rect 323458 149940 323486 150198
rect 324102 149940 324130 150198
rect 324746 149940 324774 150198
rect 325390 149940 325418 150198
rect 326034 149940 326062 150198
rect 326678 149940 326706 150198
rect 327322 149940 327350 150198
rect 327966 149940 327994 150198
rect 328460 150204 328512 150210
rect 328564 150198 328638 150226
rect 328460 150146 328512 150152
rect 328610 149940 328638 150198
rect 329242 150204 329294 150210
rect 329242 150146 329294 150152
rect 329898 150198 329972 150226
rect 330496 150226 330524 156946
rect 330956 153066 330984 163200
rect 330944 153060 330996 153066
rect 330944 153002 330996 153008
rect 331128 152176 331180 152182
rect 331128 152118 331180 152124
rect 331140 150226 331168 152118
rect 331232 151978 331260 163254
rect 331692 163146 331720 163254
rect 331770 163200 331826 164400
rect 332598 163200 332654 164400
rect 333426 163200 333482 164400
rect 334254 163200 334310 164400
rect 335082 163200 335138 164400
rect 335372 163254 335952 163282
rect 331784 163146 331812 163200
rect 331692 163118 331812 163146
rect 332416 154352 332468 154358
rect 332416 154294 332468 154300
rect 331772 152924 331824 152930
rect 331772 152866 331824 152872
rect 331220 151972 331272 151978
rect 331220 151914 331272 151920
rect 331784 150226 331812 152866
rect 332428 150226 332456 154294
rect 332612 152182 332640 163200
rect 332692 160064 332744 160070
rect 332692 160006 332744 160012
rect 332600 152176 332652 152182
rect 332600 152118 332652 152124
rect 330496 150198 330570 150226
rect 331140 150198 331214 150226
rect 331784 150198 331858 150226
rect 332428 150198 332502 150226
rect 332704 150210 332732 160006
rect 333060 157140 333112 157146
rect 333060 157082 333112 157088
rect 333072 150226 333100 157082
rect 333440 155514 333468 163200
rect 334268 160070 334296 163200
rect 334256 160064 334308 160070
rect 334256 160006 334308 160012
rect 335096 159322 335124 163200
rect 334348 159316 334400 159322
rect 334348 159258 334400 159264
rect 335084 159316 335136 159322
rect 335084 159258 335136 159264
rect 333428 155508 333480 155514
rect 333428 155450 333480 155456
rect 334360 150226 334388 159258
rect 334900 154488 334952 154494
rect 334900 154430 334952 154436
rect 334912 150226 334940 154430
rect 335372 152930 335400 163254
rect 335924 163146 335952 163254
rect 336002 163200 336058 164400
rect 336830 163200 336886 164400
rect 337658 163200 337714 164400
rect 338486 163200 338542 164400
rect 339314 163200 339370 164400
rect 339512 163254 340092 163282
rect 336016 163146 336044 163200
rect 335924 163118 336044 163146
rect 335544 157276 335596 157282
rect 335544 157218 335596 157224
rect 335360 152924 335412 152930
rect 335360 152866 335412 152872
rect 335556 150226 335584 157218
rect 336844 154222 336872 163200
rect 337672 155582 337700 163200
rect 338500 159186 338528 163200
rect 339328 159254 339356 163200
rect 338764 159248 338816 159254
rect 338764 159190 338816 159196
rect 339316 159248 339368 159254
rect 339316 159190 339368 159196
rect 338396 159180 338448 159186
rect 338396 159122 338448 159128
rect 338488 159180 338540 159186
rect 338488 159122 338540 159128
rect 338120 156732 338172 156738
rect 338120 156674 338172 156680
rect 337660 155576 337712 155582
rect 337660 155518 337712 155524
rect 337476 154556 337528 154562
rect 337476 154498 337528 154504
rect 336832 154216 336884 154222
rect 336832 154158 336884 154164
rect 336832 153196 336884 153202
rect 336832 153138 336884 153144
rect 336188 152244 336240 152250
rect 336188 152186 336240 152192
rect 336200 150226 336228 152186
rect 336844 150226 336872 153138
rect 337488 150226 337516 154498
rect 338132 150226 338160 156674
rect 329254 149940 329282 150146
rect 329898 149940 329926 150198
rect 330542 149940 330570 150198
rect 331186 149940 331214 150198
rect 331830 149940 331858 150198
rect 332474 149940 332502 150198
rect 332692 150204 332744 150210
rect 333072 150198 333146 150226
rect 332692 150146 332744 150152
rect 333118 149940 333146 150198
rect 333750 150204 333802 150210
rect 334360 150198 334434 150226
rect 334912 150198 334986 150226
rect 335556 150198 335630 150226
rect 336200 150198 336274 150226
rect 336844 150198 336918 150226
rect 337488 150198 337562 150226
rect 338132 150198 338206 150226
rect 338408 150210 338436 159122
rect 338776 150226 338804 159190
rect 339512 154290 339540 163254
rect 340064 163146 340092 163254
rect 340142 163200 340198 164400
rect 340970 163200 341026 164400
rect 341890 163200 341946 164400
rect 342718 163200 342774 164400
rect 342824 163254 343496 163282
rect 340156 163146 340184 163200
rect 340064 163118 340184 163146
rect 339684 159180 339736 159186
rect 339684 159122 339736 159128
rect 339592 155780 339644 155786
rect 339592 155722 339644 155728
rect 339500 154284 339552 154290
rect 339500 154226 339552 154232
rect 339604 151814 339632 155722
rect 339696 153202 339724 159122
rect 340052 156868 340104 156874
rect 340052 156810 340104 156816
rect 339684 153196 339736 153202
rect 339684 153138 339736 153144
rect 340064 151814 340092 156810
rect 340984 155650 341012 163200
rect 341904 159186 341932 163200
rect 342444 159520 342496 159526
rect 342444 159462 342496 159468
rect 342260 159384 342312 159390
rect 342260 159326 342312 159332
rect 341892 159180 341944 159186
rect 341892 159122 341944 159128
rect 340972 155644 341024 155650
rect 340972 155586 341024 155592
rect 342272 152998 342300 159326
rect 342352 155848 342404 155854
rect 342352 155790 342404 155796
rect 341340 152992 341392 152998
rect 341340 152934 341392 152940
rect 342260 152992 342312 152998
rect 342260 152934 342312 152940
rect 339604 151786 340000 151814
rect 340064 151786 340736 151814
rect 339972 150226 340000 151786
rect 340708 150226 340736 151786
rect 341352 150226 341380 152934
rect 341984 152380 342036 152386
rect 341984 152322 342036 152328
rect 341996 150226 342024 152322
rect 342364 151814 342392 155790
rect 342456 152250 342484 159462
rect 342732 159390 342760 163200
rect 342720 159384 342772 159390
rect 342720 159326 342772 159332
rect 342720 156936 342772 156942
rect 342720 156878 342772 156884
rect 342444 152244 342496 152250
rect 342444 152186 342496 152192
rect 342732 151814 342760 156878
rect 342824 154358 342852 163254
rect 343468 163146 343496 163254
rect 343546 163200 343602 164400
rect 344374 163200 344430 164400
rect 345202 163200 345258 164400
rect 346030 163200 346086 164400
rect 346412 163254 346808 163282
rect 343560 163146 343588 163200
rect 343468 163118 343588 163146
rect 343640 159384 343692 159390
rect 343640 159326 343692 159332
rect 342812 154352 342864 154358
rect 342812 154294 342864 154300
rect 343652 152386 343680 159326
rect 344388 155718 344416 163200
rect 345216 161474 345244 163200
rect 345216 161446 345336 161474
rect 345112 156800 345164 156806
rect 345112 156742 345164 156748
rect 344376 155712 344428 155718
rect 344376 155654 344428 155660
rect 343916 152992 343968 152998
rect 343916 152934 343968 152940
rect 343640 152380 343692 152386
rect 343640 152322 343692 152328
rect 342364 151786 342668 151814
rect 342732 151786 343312 151814
rect 342640 150226 342668 151786
rect 343284 150226 343312 151786
rect 343928 150226 343956 152934
rect 344560 152244 344612 152250
rect 344560 152186 344612 152192
rect 344572 150226 344600 152186
rect 333750 150146 333802 150152
rect 333762 149940 333790 150146
rect 334406 149940 334434 150198
rect 334958 149940 334986 150198
rect 335602 149940 335630 150198
rect 336246 149940 336274 150198
rect 336890 149940 336918 150198
rect 337534 149940 337562 150198
rect 338178 149940 338206 150198
rect 338396 150204 338448 150210
rect 338776 150198 338850 150226
rect 338396 150146 338448 150152
rect 338822 149940 338850 150198
rect 339454 150204 339506 150210
rect 339972 150198 340138 150226
rect 340708 150198 340782 150226
rect 341352 150198 341426 150226
rect 341996 150198 342070 150226
rect 342640 150198 342714 150226
rect 343284 150198 343358 150226
rect 343928 150198 344002 150226
rect 344572 150198 344646 150226
rect 345124 150210 345152 156742
rect 345204 155916 345256 155922
rect 345204 155858 345256 155864
rect 345216 150226 345244 155858
rect 345308 152998 345336 161446
rect 346044 159390 346072 163200
rect 346032 159384 346084 159390
rect 346032 159326 346084 159332
rect 346412 154426 346440 163254
rect 346780 163146 346808 163254
rect 346858 163200 346914 164400
rect 347778 163200 347834 164400
rect 347976 163254 348556 163282
rect 346872 163146 346900 163200
rect 346780 163118 346900 163146
rect 347688 159520 347740 159526
rect 347688 159462 347740 159468
rect 347700 158982 347728 159462
rect 347792 158982 347820 163200
rect 347688 158976 347740 158982
rect 347688 158918 347740 158924
rect 347780 158976 347832 158982
rect 347780 158918 347832 158924
rect 347872 155236 347924 155242
rect 347872 155178 347924 155184
rect 346400 154420 346452 154426
rect 346400 154362 346452 154368
rect 345296 152992 345348 152998
rect 345296 152934 345348 152940
rect 347136 152516 347188 152522
rect 347136 152458 347188 152464
rect 346492 151836 346544 151842
rect 346492 151778 346544 151784
rect 346504 150226 346532 151778
rect 347148 150226 347176 152458
rect 347884 150226 347912 155178
rect 347976 152522 348004 163254
rect 348528 163146 348556 163254
rect 348606 163200 348662 164400
rect 349172 163254 349384 163282
rect 348620 163146 348648 163200
rect 348528 163118 348648 163146
rect 349068 159452 349120 159458
rect 349068 159394 349120 159400
rect 348056 157208 348108 157214
rect 348056 157150 348108 157156
rect 347964 152516 348016 152522
rect 347964 152458 348016 152464
rect 348068 151814 348096 157150
rect 348068 151786 348464 151814
rect 339454 150146 339506 150152
rect 339466 149940 339494 150146
rect 340110 149940 340138 150198
rect 340754 149940 340782 150198
rect 341398 149940 341426 150198
rect 342042 149940 342070 150198
rect 342686 149940 342714 150198
rect 343330 149940 343358 150198
rect 343974 149940 344002 150198
rect 344618 149940 344646 150198
rect 345112 150204 345164 150210
rect 345216 150198 345290 150226
rect 345112 150146 345164 150152
rect 345262 149940 345290 150198
rect 345894 150204 345946 150210
rect 346504 150198 346578 150226
rect 347148 150198 347222 150226
rect 345894 150146 345946 150152
rect 345906 149940 345934 150146
rect 346550 149940 346578 150198
rect 347194 149940 347222 150198
rect 347838 150198 347912 150226
rect 348436 150226 348464 151786
rect 349080 150226 349108 159394
rect 349172 152250 349200 163254
rect 349356 163146 349384 163254
rect 349434 163200 349490 164400
rect 349540 163254 350212 163282
rect 349448 163146 349476 163200
rect 349356 163118 349476 163146
rect 349252 159656 349304 159662
rect 349252 159598 349304 159604
rect 349160 152244 349212 152250
rect 349160 152186 349212 152192
rect 349264 151814 349292 159598
rect 349540 154494 349568 163254
rect 350184 163146 350212 163254
rect 350262 163200 350318 164400
rect 351090 163200 351146 164400
rect 351918 163200 351974 164400
rect 352024 163254 352696 163282
rect 350276 163146 350304 163200
rect 350184 163118 350304 163146
rect 349804 159452 349856 159458
rect 349804 159394 349856 159400
rect 349816 159118 349844 159394
rect 349804 159112 349856 159118
rect 349804 159054 349856 159060
rect 351104 159050 351132 163200
rect 351932 159662 351960 163200
rect 351920 159656 351972 159662
rect 351920 159598 351972 159604
rect 351092 159044 351144 159050
rect 351092 158986 351144 158992
rect 350356 155168 350408 155174
rect 350356 155110 350408 155116
rect 349528 154488 349580 154494
rect 349528 154430 349580 154436
rect 349804 152380 349856 152386
rect 349804 152322 349856 152328
rect 349896 152380 349948 152386
rect 349896 152322 349948 152328
rect 349816 151842 349844 152322
rect 349908 152250 349936 152322
rect 349896 152244 349948 152250
rect 349896 152186 349948 152192
rect 349804 151836 349856 151842
rect 349264 151786 349752 151814
rect 349724 150226 349752 151786
rect 349804 151778 349856 151784
rect 350368 150226 350396 155110
rect 352024 152590 352052 163254
rect 352668 163146 352696 163254
rect 352746 163200 352802 164400
rect 353666 163200 353722 164400
rect 354494 163200 354550 164400
rect 354692 163254 355272 163282
rect 352760 163146 352788 163200
rect 352668 163118 352788 163146
rect 353208 159112 353260 159118
rect 353208 159054 353260 159060
rect 352472 155304 352524 155310
rect 352472 155246 352524 155252
rect 351644 152584 351696 152590
rect 351644 152526 351696 152532
rect 352012 152584 352064 152590
rect 352012 152526 352064 152532
rect 351000 152108 351052 152114
rect 351000 152050 351052 152056
rect 351012 150226 351040 152050
rect 351656 150226 351684 152526
rect 352288 152040 352340 152046
rect 352288 151982 352340 151988
rect 352300 150226 352328 151982
rect 352484 151814 352512 155246
rect 353220 151814 353248 159054
rect 353680 154562 353708 163200
rect 354220 159520 354272 159526
rect 354220 159462 354272 159468
rect 353668 154556 353720 154562
rect 353668 154498 353720 154504
rect 352484 151786 352972 151814
rect 353220 151786 353616 151814
rect 352944 150226 352972 151786
rect 353588 150226 353616 151786
rect 354232 150226 354260 159462
rect 354508 152250 354536 163200
rect 354496 152244 354548 152250
rect 354496 152186 354548 152192
rect 354692 152114 354720 163254
rect 355244 163146 355272 163254
rect 355322 163200 355378 164400
rect 356150 163200 356206 164400
rect 356256 163254 356928 163282
rect 355336 163146 355364 163200
rect 355244 163118 355364 163146
rect 356164 159526 356192 163200
rect 356152 159520 356204 159526
rect 356152 159462 356204 159468
rect 354864 159452 354916 159458
rect 354864 159394 354916 159400
rect 354680 152108 354732 152114
rect 354680 152050 354732 152056
rect 354876 150226 354904 159394
rect 356256 153882 356284 163254
rect 356900 163146 356928 163254
rect 356978 163200 357034 164400
rect 357806 163200 357862 164400
rect 358634 163200 358690 164400
rect 358832 163254 359504 163282
rect 356992 163146 357020 163200
rect 356900 163118 357020 163146
rect 357820 159118 357848 163200
rect 357992 159724 358044 159730
rect 357992 159666 358044 159672
rect 357808 159112 357860 159118
rect 357808 159054 357860 159060
rect 357440 158908 357492 158914
rect 357440 158850 357492 158856
rect 355508 153876 355560 153882
rect 355508 153818 355560 153824
rect 356244 153876 356296 153882
rect 356244 153818 356296 153824
rect 355520 150226 355548 153818
rect 357452 152862 357480 158850
rect 357900 154012 357952 154018
rect 357900 153954 357952 153960
rect 356152 152856 356204 152862
rect 356152 152798 356204 152804
rect 357440 152856 357492 152862
rect 357440 152798 357492 152804
rect 356164 150226 356192 152798
rect 356796 152652 356848 152658
rect 356796 152594 356848 152600
rect 356808 150226 356836 152594
rect 357438 152416 357494 152425
rect 357438 152351 357494 152360
rect 357452 150226 357480 152351
rect 357912 150498 357940 153954
rect 358004 151814 358032 159666
rect 358648 159458 358676 163200
rect 358636 159452 358688 159458
rect 358636 159394 358688 159400
rect 358832 152658 358860 163254
rect 359476 163146 359504 163254
rect 359554 163200 359610 164400
rect 360382 163200 360438 164400
rect 361210 163200 361266 164400
rect 361592 163254 361988 163282
rect 359568 163146 359596 163200
rect 359476 163118 359596 163146
rect 358912 159588 358964 159594
rect 358912 159530 358964 159536
rect 358820 152652 358872 152658
rect 358820 152594 358872 152600
rect 358004 151786 358768 151814
rect 357912 150470 358124 150498
rect 358096 150226 358124 150470
rect 358740 150226 358768 151786
rect 348436 150198 348510 150226
rect 349080 150198 349154 150226
rect 349724 150198 349798 150226
rect 350368 150198 350442 150226
rect 351012 150198 351086 150226
rect 351656 150198 351730 150226
rect 352300 150198 352374 150226
rect 352944 150198 353018 150226
rect 353588 150198 353662 150226
rect 354232 150198 354306 150226
rect 354876 150198 354950 150226
rect 355520 150198 355594 150226
rect 356164 150198 356238 150226
rect 356808 150198 356882 150226
rect 357452 150198 357526 150226
rect 358096 150198 358170 150226
rect 358740 150198 358814 150226
rect 358924 150210 358952 159530
rect 360396 153814 360424 163200
rect 361224 158914 361252 163200
rect 361212 158908 361264 158914
rect 361212 158850 361264 158856
rect 360660 153944 360712 153950
rect 360660 153886 360712 153892
rect 360384 153808 360436 153814
rect 360384 153750 360436 153756
rect 359372 152856 359424 152862
rect 359372 152798 359424 152804
rect 359384 150226 359412 152798
rect 360672 150226 360700 153886
rect 361592 152862 361620 163254
rect 361960 163146 361988 163254
rect 362038 163200 362094 164400
rect 362866 163200 362922 164400
rect 363064 163254 363644 163282
rect 362052 163146 362080 163200
rect 361960 163118 362080 163146
rect 362880 159594 362908 163200
rect 362960 159860 363012 159866
rect 362960 159802 363012 159808
rect 362868 159588 362920 159594
rect 362868 159530 362920 159536
rect 361580 152856 361632 152862
rect 361580 152798 361632 152804
rect 361948 152720 362000 152726
rect 361948 152662 362000 152668
rect 361304 152448 361356 152454
rect 361304 152390 361356 152396
rect 361316 150226 361344 152390
rect 361960 150226 361988 152662
rect 362592 151904 362644 151910
rect 362592 151846 362644 151852
rect 362604 150226 362632 151846
rect 347838 149940 347866 150198
rect 348482 149940 348510 150198
rect 349126 149940 349154 150198
rect 349770 149940 349798 150198
rect 350414 149940 350442 150198
rect 351058 149940 351086 150198
rect 351702 149940 351730 150198
rect 352346 149940 352374 150198
rect 352990 149940 353018 150198
rect 353634 149940 353662 150198
rect 354278 149940 354306 150198
rect 354922 149940 354950 150198
rect 355566 149940 355594 150198
rect 356210 149940 356238 150198
rect 356854 149940 356882 150198
rect 357498 149940 357526 150198
rect 358142 149940 358170 150198
rect 358786 149940 358814 150198
rect 358912 150204 358964 150210
rect 359384 150198 359458 150226
rect 358912 150146 358964 150152
rect 359430 149940 359458 150198
rect 360062 150204 360114 150210
rect 360672 150198 360746 150226
rect 361316 150198 361390 150226
rect 361960 150198 362034 150226
rect 362604 150198 362678 150226
rect 362972 150210 363000 159802
rect 363064 153950 363092 163254
rect 363616 163146 363644 163254
rect 363694 163200 363750 164400
rect 364522 163200 364578 164400
rect 365442 163200 365498 164400
rect 365732 163254 366220 163282
rect 363708 163146 363736 163200
rect 363616 163118 363736 163146
rect 363144 158840 363196 158846
rect 363144 158782 363196 158788
rect 363052 153944 363104 153950
rect 363052 153886 363104 153892
rect 363156 151910 363184 158782
rect 363236 155372 363288 155378
rect 363236 155314 363288 155320
rect 363144 151904 363196 151910
rect 363144 151846 363196 151852
rect 363248 150226 363276 155314
rect 364536 152046 364564 163200
rect 365456 159798 365484 163200
rect 365168 159792 365220 159798
rect 365168 159734 365220 159740
rect 365444 159792 365496 159798
rect 365444 159734 365496 159740
rect 364524 152040 364576 152046
rect 364524 151982 364576 151988
rect 364524 151904 364576 151910
rect 364524 151846 364576 151852
rect 364536 150226 364564 151846
rect 365180 150226 365208 159734
rect 365732 152454 365760 163254
rect 366192 163146 366220 163254
rect 366270 163200 366326 164400
rect 367098 163200 367154 164400
rect 367926 163200 367982 164400
rect 368492 163254 368704 163282
rect 366284 163146 366312 163200
rect 366192 163118 366312 163146
rect 365812 154080 365864 154086
rect 365812 154022 365864 154028
rect 365720 152448 365772 152454
rect 365720 152390 365772 152396
rect 365824 150226 365852 154022
rect 367112 154018 367140 163200
rect 367940 158846 367968 163200
rect 367928 158840 367980 158846
rect 367928 158782 367980 158788
rect 367192 158772 367244 158778
rect 367192 158714 367244 158720
rect 367100 154012 367152 154018
rect 367100 153954 367152 153960
rect 367204 153134 367232 158714
rect 368296 154148 368348 154154
rect 368296 154090 368348 154096
rect 367008 153128 367060 153134
rect 367008 153070 367060 153076
rect 367192 153128 367244 153134
rect 367192 153070 367244 153076
rect 366364 152788 366416 152794
rect 366364 152730 366416 152736
rect 360062 150146 360114 150152
rect 360074 149940 360102 150146
rect 360718 149940 360746 150198
rect 361362 149940 361390 150198
rect 362006 149940 362034 150198
rect 362650 149940 362678 150198
rect 362960 150204 363012 150210
rect 363248 150198 363322 150226
rect 362960 150146 363012 150152
rect 363294 149940 363322 150198
rect 363926 150204 363978 150210
rect 364536 150198 364610 150226
rect 365180 150198 365254 150226
rect 363926 150146 363978 150152
rect 363938 149940 363966 150146
rect 364582 149940 364610 150198
rect 365226 149940 365254 150198
rect 365778 150198 365852 150226
rect 366376 150226 366404 152730
rect 367020 150226 367048 153070
rect 367652 152312 367704 152318
rect 367652 152254 367704 152260
rect 367664 150226 367692 152254
rect 368308 150226 368336 154090
rect 368492 152726 368520 163254
rect 368676 163146 368704 163254
rect 368754 163200 368810 164400
rect 369582 163200 369638 164400
rect 370410 163200 370466 164400
rect 371330 163200 371386 164400
rect 372158 163200 372214 164400
rect 372632 163254 372936 163282
rect 368768 163146 368796 163200
rect 368676 163118 368796 163146
rect 369492 159928 369544 159934
rect 369492 159870 369544 159876
rect 368940 153128 368992 153134
rect 368940 153070 368992 153076
rect 368480 152720 368532 152726
rect 368480 152662 368532 152668
rect 368952 150226 368980 153070
rect 369504 151814 369532 159870
rect 369596 159730 369624 163200
rect 369952 159996 370004 160002
rect 369952 159938 370004 159944
rect 369584 159724 369636 159730
rect 369584 159666 369636 159672
rect 369964 151814 369992 159938
rect 370424 155242 370452 163200
rect 370872 155440 370924 155446
rect 370872 155382 370924 155388
rect 370412 155236 370464 155242
rect 370412 155178 370464 155184
rect 369504 151786 369624 151814
rect 369964 151786 370268 151814
rect 369596 150226 369624 151786
rect 370240 150226 370268 151786
rect 370884 150226 370912 155382
rect 371344 152318 371372 163200
rect 372172 160002 372200 163200
rect 372160 159996 372212 160002
rect 372160 159938 372212 159944
rect 371516 153060 371568 153066
rect 371516 153002 371568 153008
rect 371332 152312 371384 152318
rect 371332 152254 371384 152260
rect 371528 150226 371556 153002
rect 372632 152794 372660 163254
rect 372908 163146 372936 163254
rect 372986 163200 373042 164400
rect 373814 163200 373870 164400
rect 374642 163200 374698 164400
rect 375470 163200 375526 164400
rect 376298 163200 376354 164400
rect 376864 163254 377168 163282
rect 373000 163146 373028 163200
rect 372908 163118 373028 163146
rect 373448 155508 373500 155514
rect 373448 155450 373500 155456
rect 372620 152788 372672 152794
rect 372620 152730 372672 152736
rect 372804 152176 372856 152182
rect 372804 152118 372856 152124
rect 372160 151972 372212 151978
rect 372160 151914 372212 151920
rect 372172 150226 372200 151914
rect 372816 150226 372844 152118
rect 373460 150226 373488 155450
rect 373828 155310 373856 163200
rect 374092 160064 374144 160070
rect 374092 160006 374144 160012
rect 373816 155304 373868 155310
rect 373816 155246 373868 155252
rect 374104 150226 374132 160006
rect 374656 158778 374684 163200
rect 374736 159316 374788 159322
rect 374736 159258 374788 159264
rect 374644 158772 374696 158778
rect 374644 158714 374696 158720
rect 374748 150226 374776 159258
rect 375484 153066 375512 163200
rect 376312 159866 376340 163200
rect 376300 159860 376352 159866
rect 376300 159802 376352 159808
rect 375564 155576 375616 155582
rect 375564 155518 375616 155524
rect 375472 153060 375524 153066
rect 375472 153002 375524 153008
rect 375380 152924 375432 152930
rect 375380 152866 375432 152872
rect 375392 150226 375420 152866
rect 366376 150198 366450 150226
rect 367020 150198 367094 150226
rect 367664 150198 367738 150226
rect 368308 150198 368382 150226
rect 368952 150198 369026 150226
rect 369596 150198 369670 150226
rect 370240 150198 370314 150226
rect 370884 150198 370958 150226
rect 371528 150198 371602 150226
rect 372172 150198 372246 150226
rect 372816 150198 372890 150226
rect 373460 150198 373534 150226
rect 374104 150198 374178 150226
rect 374748 150198 374822 150226
rect 375392 150198 375466 150226
rect 375576 150210 375604 155518
rect 376024 154216 376076 154222
rect 376024 154158 376076 154164
rect 376036 150226 376064 154158
rect 376864 154154 376892 163254
rect 377140 163146 377168 163254
rect 377218 163200 377274 164400
rect 378046 163200 378102 164400
rect 378874 163200 378930 164400
rect 379702 163200 379758 164400
rect 380176 163254 380480 163282
rect 377232 163146 377260 163200
rect 377140 163118 377260 163146
rect 378060 159322 378088 163200
rect 378888 160070 378916 163200
rect 378876 160064 378928 160070
rect 378876 160006 378928 160012
rect 379716 159934 379744 163200
rect 379704 159928 379756 159934
rect 379704 159870 379756 159876
rect 378048 159316 378100 159322
rect 378048 159258 378100 159264
rect 377956 159248 378008 159254
rect 377956 159190 378008 159196
rect 376852 154148 376904 154154
rect 376852 154090 376904 154096
rect 377312 153196 377364 153202
rect 377312 153138 377364 153144
rect 377324 150226 377352 153138
rect 377968 150226 377996 159190
rect 378232 159180 378284 159186
rect 378232 159122 378284 159128
rect 378140 155644 378192 155650
rect 378140 155586 378192 155592
rect 365778 149940 365806 150198
rect 366422 149940 366450 150198
rect 367066 149940 367094 150198
rect 367710 149940 367738 150198
rect 368354 149940 368382 150198
rect 368998 149940 369026 150198
rect 369642 149940 369670 150198
rect 370286 149940 370314 150198
rect 370930 149940 370958 150198
rect 371574 149940 371602 150198
rect 372218 149940 372246 150198
rect 372862 149940 372890 150198
rect 373506 149940 373534 150198
rect 374150 149940 374178 150198
rect 374794 149940 374822 150198
rect 375438 149940 375466 150198
rect 375564 150204 375616 150210
rect 376036 150198 376110 150226
rect 375564 150146 375616 150152
rect 376082 149940 376110 150198
rect 376714 150204 376766 150210
rect 377324 150198 377398 150226
rect 377968 150198 378042 150226
rect 378152 150210 378180 155586
rect 378244 153202 378272 159122
rect 378784 158976 378836 158982
rect 378784 158918 378836 158924
rect 378600 154284 378652 154290
rect 378600 154226 378652 154232
rect 378232 153196 378284 153202
rect 378232 153138 378284 153144
rect 378612 150226 378640 154226
rect 378796 151978 378824 158918
rect 380176 154086 380204 163254
rect 380452 163146 380480 163254
rect 380530 163200 380586 164400
rect 381004 163254 381308 163282
rect 380544 163146 380572 163200
rect 380452 163118 380572 163146
rect 380164 154080 380216 154086
rect 380164 154022 380216 154028
rect 379888 153196 379940 153202
rect 379888 153138 379940 153144
rect 378784 151972 378836 151978
rect 378784 151914 378836 151920
rect 379900 150226 379928 153138
rect 381004 153134 381032 163254
rect 381280 163146 381308 163254
rect 381358 163200 381414 164400
rect 382186 163200 382242 164400
rect 383106 163200 383162 164400
rect 383672 163254 383884 163282
rect 381372 163146 381400 163200
rect 381280 163118 381400 163146
rect 381820 155712 381872 155718
rect 381820 155654 381872 155660
rect 381176 154352 381228 154358
rect 381176 154294 381228 154300
rect 380992 153128 381044 153134
rect 380992 153070 381044 153076
rect 380532 151836 380584 151842
rect 380532 151778 380584 151784
rect 380544 150226 380572 151778
rect 381188 150226 381216 154294
rect 381832 150226 381860 155654
rect 382200 152930 382228 163200
rect 382832 159384 382884 159390
rect 382832 159326 382884 159332
rect 382556 159044 382608 159050
rect 382556 158986 382608 158992
rect 382568 152998 382596 158986
rect 382464 152992 382516 152998
rect 382464 152934 382516 152940
rect 382556 152992 382608 152998
rect 382556 152934 382608 152940
rect 382188 152924 382240 152930
rect 382188 152866 382240 152872
rect 382476 150226 382504 152934
rect 382844 151814 382872 159326
rect 383120 159186 383148 163200
rect 383108 159180 383160 159186
rect 383108 159122 383160 159128
rect 383672 154222 383700 163254
rect 383856 163146 383884 163254
rect 383934 163200 383990 164400
rect 384762 163200 384818 164400
rect 385590 163200 385646 164400
rect 386418 163200 386474 164400
rect 386524 163254 387196 163282
rect 383948 163146 383976 163200
rect 383856 163118 383976 163146
rect 384776 158982 384804 163200
rect 385604 159254 385632 163200
rect 385776 159656 385828 159662
rect 385776 159598 385828 159604
rect 385592 159248 385644 159254
rect 385592 159190 385644 159196
rect 384948 159112 385000 159118
rect 384948 159054 385000 159060
rect 384764 158976 384816 158982
rect 384764 158918 384816 158924
rect 383752 154420 383804 154426
rect 383752 154362 383804 154368
rect 383660 154216 383712 154222
rect 383660 154158 383712 154164
rect 382844 151786 383148 151814
rect 383120 150226 383148 151786
rect 383764 150226 383792 154362
rect 384960 152182 384988 159054
rect 385040 158840 385092 158846
rect 385040 158782 385092 158788
rect 385052 153202 385080 158782
rect 385040 153196 385092 153202
rect 385040 153138 385092 153144
rect 385040 152516 385092 152522
rect 385040 152458 385092 152464
rect 384948 152176 385000 152182
rect 384948 152118 385000 152124
rect 384396 151972 384448 151978
rect 384396 151914 384448 151920
rect 384408 150226 384436 151914
rect 385052 150226 385080 152458
rect 385788 152386 385816 159598
rect 386328 158908 386380 158914
rect 386328 158850 386380 158856
rect 386236 154488 386288 154494
rect 386236 154430 386288 154436
rect 385684 152380 385736 152386
rect 385684 152322 385736 152328
rect 385776 152380 385828 152386
rect 385776 152322 385828 152328
rect 385696 150226 385724 152322
rect 386248 151814 386276 154430
rect 386340 151910 386368 158850
rect 386432 152522 386460 163200
rect 386524 154290 386552 163254
rect 387168 163146 387196 163254
rect 387246 163200 387302 164400
rect 388074 163200 388130 164400
rect 388994 163200 389050 164400
rect 389822 163200 389878 164400
rect 390650 163200 390706 164400
rect 391478 163200 391534 164400
rect 392306 163200 392362 164400
rect 393134 163200 393190 164400
rect 393332 163254 393912 163282
rect 387260 163146 387288 163200
rect 387168 163118 387288 163146
rect 388088 159662 388116 163200
rect 388076 159656 388128 159662
rect 388076 159598 388128 159604
rect 389008 159322 389036 163200
rect 389836 159662 389864 163200
rect 389088 159656 389140 159662
rect 389088 159598 389140 159604
rect 389824 159656 389876 159662
rect 389824 159598 389876 159604
rect 388352 159316 388404 159322
rect 388352 159258 388404 159264
rect 388996 159316 389048 159322
rect 388996 159258 389048 159264
rect 386512 154284 386564 154290
rect 386512 154226 386564 154232
rect 386972 152992 387024 152998
rect 386972 152934 387024 152940
rect 386420 152516 386472 152522
rect 386420 152458 386472 152464
rect 386328 151904 386380 151910
rect 386328 151846 386380 151852
rect 386248 151786 386368 151814
rect 386340 150226 386368 151786
rect 386984 150226 387012 152934
rect 388364 152590 388392 159258
rect 389100 158846 389128 159598
rect 390560 159520 390612 159526
rect 390560 159462 390612 159468
rect 389088 158840 389140 158846
rect 389088 158782 389140 158788
rect 390376 158840 390428 158846
rect 390376 158782 390428 158788
rect 388444 158772 388496 158778
rect 388444 158714 388496 158720
rect 389180 158772 389232 158778
rect 389180 158714 389232 158720
rect 388260 152584 388312 152590
rect 388260 152526 388312 152532
rect 388352 152584 388404 152590
rect 388352 152526 388404 152532
rect 387616 152380 387668 152386
rect 387616 152322 387668 152328
rect 387628 150226 387656 152322
rect 388272 150226 388300 152526
rect 388456 151978 388484 158714
rect 388904 154556 388956 154562
rect 388904 154498 388956 154504
rect 388444 151972 388496 151978
rect 388444 151914 388496 151920
rect 388916 150226 388944 154498
rect 389192 152386 389220 158714
rect 390388 152998 390416 158782
rect 390376 152992 390428 152998
rect 390376 152934 390428 152940
rect 389180 152380 389232 152386
rect 389180 152322 389232 152328
rect 389548 152244 389600 152250
rect 389548 152186 389600 152192
rect 389560 150226 389588 152186
rect 390192 152108 390244 152114
rect 390192 152050 390244 152056
rect 390204 150226 390232 152050
rect 390572 151814 390600 159462
rect 390664 154494 390692 163200
rect 391492 160070 391520 163200
rect 391388 160064 391440 160070
rect 391388 160006 391440 160012
rect 391480 160064 391532 160070
rect 391480 160006 391532 160012
rect 391400 159526 391428 160006
rect 391388 159520 391440 159526
rect 391388 159462 391440 159468
rect 392320 159186 392348 163200
rect 392768 159452 392820 159458
rect 392768 159394 392820 159400
rect 392308 159180 392360 159186
rect 392308 159122 392360 159128
rect 390652 154488 390704 154494
rect 390652 154430 390704 154436
rect 391480 153876 391532 153882
rect 391480 153818 391532 153824
rect 390572 151786 390876 151814
rect 390848 150226 390876 151786
rect 391492 150226 391520 153818
rect 392216 152584 392268 152590
rect 392216 152526 392268 152532
rect 392228 152182 392256 152526
rect 392124 152176 392176 152182
rect 392124 152118 392176 152124
rect 392216 152176 392268 152182
rect 392216 152118 392268 152124
rect 392136 150226 392164 152118
rect 392780 150226 392808 159394
rect 393148 152590 393176 163200
rect 393332 154358 393360 163254
rect 393884 163146 393912 163254
rect 393962 163200 394018 164400
rect 394882 163200 394938 164400
rect 395710 163200 395766 164400
rect 396538 163200 396594 164400
rect 397366 163200 397422 164400
rect 397472 163254 398144 163282
rect 393976 163146 394004 163200
rect 393884 163118 394004 163146
rect 394608 160064 394660 160070
rect 394608 160006 394660 160012
rect 393320 154352 393372 154358
rect 393320 154294 393372 154300
rect 394056 153808 394108 153814
rect 394056 153750 394108 153756
rect 393412 152652 393464 152658
rect 393412 152594 393464 152600
rect 393136 152584 393188 152590
rect 393136 152526 393188 152532
rect 393424 150226 393452 152594
rect 394068 150226 394096 153750
rect 394620 152250 394648 160006
rect 394896 152658 394924 163200
rect 395528 159792 395580 159798
rect 395528 159734 395580 159740
rect 394976 159588 395028 159594
rect 394976 159530 395028 159536
rect 394884 152652 394936 152658
rect 394884 152594 394936 152600
rect 394608 152244 394660 152250
rect 394608 152186 394660 152192
rect 394700 151904 394752 151910
rect 394700 151846 394752 151852
rect 394712 150226 394740 151846
rect 376714 150146 376766 150152
rect 376726 149940 376754 150146
rect 377370 149940 377398 150198
rect 378014 149940 378042 150198
rect 378140 150204 378192 150210
rect 378612 150198 378686 150226
rect 378140 150146 378192 150152
rect 378658 149940 378686 150198
rect 379290 150204 379342 150210
rect 379900 150198 379974 150226
rect 380544 150198 380618 150226
rect 381188 150198 381262 150226
rect 381832 150198 381906 150226
rect 382476 150198 382550 150226
rect 383120 150198 383194 150226
rect 383764 150198 383838 150226
rect 384408 150198 384482 150226
rect 385052 150198 385126 150226
rect 385696 150198 385770 150226
rect 386340 150198 386414 150226
rect 386984 150198 387058 150226
rect 387628 150198 387702 150226
rect 388272 150198 388346 150226
rect 388916 150198 388990 150226
rect 389560 150198 389634 150226
rect 390204 150198 390278 150226
rect 390848 150198 390922 150226
rect 391492 150198 391566 150226
rect 392136 150198 392210 150226
rect 392780 150198 392854 150226
rect 393424 150198 393498 150226
rect 394068 150198 394142 150226
rect 394712 150198 394786 150226
rect 394988 150210 395016 159530
rect 395160 159316 395212 159322
rect 395160 159258 395212 159264
rect 395172 159050 395200 159258
rect 395160 159044 395212 159050
rect 395160 158986 395212 158992
rect 395540 152862 395568 159734
rect 395724 159118 395752 163200
rect 396172 159996 396224 160002
rect 396172 159938 396224 159944
rect 395712 159112 395764 159118
rect 395712 159054 395764 159060
rect 395252 152856 395304 152862
rect 395252 152798 395304 152804
rect 395528 152856 395580 152862
rect 395528 152798 395580 152804
rect 395264 151814 395292 152798
rect 396184 151910 396212 159938
rect 396552 159798 396580 163200
rect 396540 159792 396592 159798
rect 396540 159734 396592 159740
rect 397380 154426 397408 163200
rect 397368 154420 397420 154426
rect 397368 154362 397420 154368
rect 396540 153944 396592 153950
rect 396540 153886 396592 153892
rect 396172 151904 396224 151910
rect 396172 151846 396224 151852
rect 395264 151786 395384 151814
rect 395356 150226 395384 151786
rect 396552 150226 396580 153886
rect 397472 153882 397500 163254
rect 398116 163146 398144 163254
rect 398194 163200 398250 164400
rect 399022 163200 399078 164400
rect 399128 163254 399800 163282
rect 398208 163146 398236 163200
rect 398116 163118 398236 163146
rect 399036 159594 399064 163200
rect 399024 159588 399076 159594
rect 399024 159530 399076 159536
rect 398564 159520 398616 159526
rect 398564 159462 398616 159468
rect 397460 153876 397512 153882
rect 397460 153818 397512 153824
rect 398104 153060 398156 153066
rect 398104 153002 398156 153008
rect 397828 152856 397880 152862
rect 397828 152798 397880 152804
rect 397184 152040 397236 152046
rect 397184 151982 397236 151988
rect 397196 150226 397224 151982
rect 397840 150226 397868 152798
rect 398116 151842 398144 153002
rect 398576 152454 398604 159462
rect 398840 159248 398892 159254
rect 398840 159190 398892 159196
rect 398472 152448 398524 152454
rect 398472 152390 398524 152396
rect 398564 152448 398616 152454
rect 398564 152390 398616 152396
rect 398104 151836 398156 151842
rect 398104 151778 398156 151784
rect 398484 150226 398512 152390
rect 398852 152114 398880 159190
rect 399128 157334 399156 163254
rect 399772 163146 399800 163254
rect 399850 163200 399906 164400
rect 400770 163200 400826 164400
rect 401598 163200 401654 164400
rect 402426 163200 402482 164400
rect 403254 163200 403310 164400
rect 404082 163200 404138 164400
rect 404372 163254 404860 163282
rect 399864 163146 399892 163200
rect 399772 163118 399892 163146
rect 400784 160070 400812 163200
rect 400772 160064 400824 160070
rect 400772 160006 400824 160012
rect 401048 159724 401100 159730
rect 401048 159666 401100 159672
rect 399128 157306 399248 157334
rect 399116 154012 399168 154018
rect 399116 153954 399168 153960
rect 398840 152108 398892 152114
rect 398840 152050 398892 152056
rect 379290 150146 379342 150152
rect 379302 149940 379330 150146
rect 379946 149940 379974 150198
rect 380590 149940 380618 150198
rect 381234 149940 381262 150198
rect 381878 149940 381906 150198
rect 382522 149940 382550 150198
rect 383166 149940 383194 150198
rect 383810 149940 383838 150198
rect 384454 149940 384482 150198
rect 385098 149940 385126 150198
rect 385742 149940 385770 150198
rect 386386 149940 386414 150198
rect 387030 149940 387058 150198
rect 387674 149940 387702 150198
rect 388318 149940 388346 150198
rect 388962 149940 388990 150198
rect 389606 149940 389634 150198
rect 390250 149940 390278 150198
rect 390894 149940 390922 150198
rect 391538 149940 391566 150198
rect 392182 149940 392210 150198
rect 392826 149940 392854 150198
rect 393470 149940 393498 150198
rect 394114 149940 394142 150198
rect 394758 149940 394786 150198
rect 394976 150204 395028 150210
rect 395356 150198 395430 150226
rect 394976 150146 395028 150152
rect 395402 149940 395430 150198
rect 396034 150204 396086 150210
rect 396552 150198 396626 150226
rect 397196 150198 397270 150226
rect 397840 150198 397914 150226
rect 398484 150198 398558 150226
rect 396034 150146 396086 150152
rect 396046 149940 396074 150146
rect 396598 149940 396626 150198
rect 397242 149940 397270 150198
rect 397886 149940 397914 150198
rect 398530 149940 398558 150198
rect 399128 150090 399156 153954
rect 399220 152862 399248 157306
rect 399760 153196 399812 153202
rect 399760 153138 399812 153144
rect 399208 152856 399260 152862
rect 399208 152798 399260 152804
rect 399772 150090 399800 153138
rect 400404 152720 400456 152726
rect 400404 152662 400456 152668
rect 400416 150090 400444 152662
rect 401060 150226 401088 159666
rect 401612 153950 401640 163200
rect 401692 155236 401744 155242
rect 401692 155178 401744 155184
rect 401600 153944 401652 153950
rect 401600 153886 401652 153892
rect 401060 150198 401134 150226
rect 399128 150062 399202 150090
rect 399772 150062 399846 150090
rect 400416 150062 400490 150090
rect 399174 149940 399202 150062
rect 399818 149940 399846 150062
rect 400462 149940 400490 150062
rect 401106 149940 401134 150198
rect 401704 150090 401732 155178
rect 402440 153202 402468 163200
rect 403268 160002 403296 163200
rect 403256 159996 403308 160002
rect 403256 159938 403308 159944
rect 404096 159458 404124 163200
rect 404084 159452 404136 159458
rect 404084 159394 404136 159400
rect 404268 159180 404320 159186
rect 404268 159122 404320 159128
rect 404176 159044 404228 159050
rect 404176 158986 404228 158992
rect 404084 155304 404136 155310
rect 404084 155246 404136 155252
rect 402428 153196 402480 153202
rect 402428 153138 402480 153144
rect 403624 152788 403676 152794
rect 403624 152730 403676 152736
rect 402336 152312 402388 152318
rect 402336 152254 402388 152260
rect 402348 150090 402376 152254
rect 402980 151904 403032 151910
rect 402980 151846 403032 151852
rect 402992 150226 403020 151846
rect 402992 150198 403066 150226
rect 401704 150062 401778 150090
rect 402348 150062 402422 150090
rect 401750 149940 401778 150062
rect 402394 149940 402422 150062
rect 403038 149940 403066 150198
rect 403636 150090 403664 152730
rect 404096 150226 404124 155246
rect 404188 151910 404216 158986
rect 404280 152318 404308 159122
rect 404372 152726 404400 163254
rect 404832 163146 404860 163254
rect 404910 163200 404966 164400
rect 405738 163200 405794 164400
rect 406658 163200 406714 164400
rect 407486 163200 407542 164400
rect 407592 163254 408264 163282
rect 404924 163146 404952 163200
rect 404832 163118 404952 163146
rect 405648 159112 405700 159118
rect 405648 159054 405700 159060
rect 404360 152720 404412 152726
rect 404360 152662 404412 152668
rect 404268 152312 404320 152318
rect 404268 152254 404320 152260
rect 405096 152312 405148 152318
rect 405096 152254 405148 152260
rect 405108 152046 405136 152254
rect 405660 152114 405688 159054
rect 405752 158778 405780 163200
rect 405832 159928 405884 159934
rect 405832 159870 405884 159876
rect 405740 158772 405792 158778
rect 405740 158714 405792 158720
rect 405844 153066 405872 159870
rect 406200 159860 406252 159866
rect 406200 159802 406252 159808
rect 405832 153060 405884 153066
rect 405832 153002 405884 153008
rect 405648 152108 405700 152114
rect 405648 152050 405700 152056
rect 405096 152040 405148 152046
rect 405096 151982 405148 151988
rect 404912 151972 404964 151978
rect 404912 151914 404964 151920
rect 404176 151904 404228 151910
rect 404176 151846 404228 151852
rect 404096 150198 404354 150226
rect 403636 150062 403710 150090
rect 403682 149940 403710 150062
rect 404326 149940 404354 150198
rect 404924 150090 404952 151914
rect 405556 151836 405608 151842
rect 405556 151778 405608 151784
rect 405568 150226 405596 151778
rect 406212 150226 406240 159802
rect 406672 152794 406700 163200
rect 407500 159730 407528 163200
rect 407488 159724 407540 159730
rect 407488 159666 407540 159672
rect 406844 154148 406896 154154
rect 406844 154090 406896 154096
rect 406660 152788 406712 152794
rect 406660 152730 406712 152736
rect 405568 150198 405642 150226
rect 406212 150198 406286 150226
rect 404924 150062 404998 150090
rect 404970 149940 404998 150062
rect 405614 149940 405642 150198
rect 406258 149940 406286 150198
rect 406856 150090 406884 154090
rect 407592 152425 407620 163254
rect 408236 163146 408264 163254
rect 408314 163200 408370 164400
rect 409142 163200 409198 164400
rect 409970 163200 410026 164400
rect 410798 163200 410854 164400
rect 411272 163254 411576 163282
rect 408328 163146 408356 163200
rect 408236 163118 408356 163146
rect 408500 159588 408552 159594
rect 408500 159530 408552 159536
rect 408132 152448 408184 152454
rect 407578 152416 407634 152425
rect 408132 152390 408184 152396
rect 407578 152351 407634 152360
rect 407488 152176 407540 152182
rect 407488 152118 407540 152124
rect 407500 150090 407528 152118
rect 408144 150090 408172 152390
rect 408512 152182 408540 159530
rect 409156 158846 409184 163200
rect 409984 159866 410012 163200
rect 409972 159860 410024 159866
rect 409972 159802 410024 159808
rect 410812 159594 410840 163200
rect 410800 159588 410852 159594
rect 410800 159530 410852 159536
rect 409144 158840 409196 158846
rect 409144 158782 409196 158788
rect 410708 158840 410760 158846
rect 410708 158782 410760 158788
rect 409236 158772 409288 158778
rect 409236 158714 409288 158720
rect 408776 153060 408828 153066
rect 408776 153002 408828 153008
rect 408500 152176 408552 152182
rect 408500 152118 408552 152124
rect 408788 150226 408816 153002
rect 409248 152318 409276 158714
rect 409420 154080 409472 154086
rect 409420 154022 409472 154028
rect 409236 152312 409288 152318
rect 409236 152254 409288 152260
rect 409432 150226 409460 154022
rect 410720 153134 410748 158782
rect 410064 153128 410116 153134
rect 410064 153070 410116 153076
rect 410708 153128 410760 153134
rect 410708 153070 410760 153076
rect 410076 150226 410104 153070
rect 411272 152930 411300 163254
rect 411548 163146 411576 163254
rect 411626 163200 411682 164400
rect 412546 163200 412602 164400
rect 413374 163200 413430 164400
rect 414202 163200 414258 164400
rect 414400 163254 414980 163282
rect 411640 163146 411668 163200
rect 411548 163118 411668 163146
rect 411352 158976 411404 158982
rect 411352 158918 411404 158924
rect 410708 152924 410760 152930
rect 410708 152866 410760 152872
rect 411260 152924 411312 152930
rect 411260 152866 411312 152872
rect 410720 150226 410748 152866
rect 411364 150226 411392 158918
rect 412560 158914 412588 163200
rect 413388 159798 413416 163200
rect 413192 159792 413244 159798
rect 413192 159734 413244 159740
rect 413376 159792 413428 159798
rect 413376 159734 413428 159740
rect 412548 158908 412600 158914
rect 412548 158850 412600 158856
rect 412824 158908 412876 158914
rect 412824 158850 412876 158856
rect 411996 154216 412048 154222
rect 411996 154158 412048 154164
rect 412008 150226 412036 154158
rect 412836 152454 412864 158850
rect 412824 152448 412876 152454
rect 412824 152390 412876 152396
rect 412640 152380 412692 152386
rect 412640 152322 412692 152328
rect 412652 150226 412680 152322
rect 413204 151910 413232 159734
rect 413376 159656 413428 159662
rect 413376 159598 413428 159604
rect 413388 153066 413416 159598
rect 414216 159390 414244 163200
rect 414204 159384 414256 159390
rect 414204 159326 414256 159332
rect 413376 153060 413428 153066
rect 413376 153002 413428 153008
rect 414400 152522 414428 163254
rect 414952 163146 414980 163254
rect 415030 163200 415086 164400
rect 415412 163254 415808 163282
rect 415044 163146 415072 163200
rect 414952 163118 415072 163146
rect 414572 154284 414624 154290
rect 414572 154226 414624 154232
rect 413928 152516 413980 152522
rect 413928 152458 413980 152464
rect 414388 152516 414440 152522
rect 414388 152458 414440 152464
rect 413284 151972 413336 151978
rect 413284 151914 413336 151920
rect 413192 151904 413244 151910
rect 413192 151846 413244 151852
rect 413296 150226 413324 151914
rect 413940 150226 413968 152458
rect 414584 150226 414612 154226
rect 415412 152998 415440 163254
rect 415780 163146 415808 163254
rect 415858 163200 415914 164400
rect 416686 163200 416742 164400
rect 417514 163200 417570 164400
rect 418434 163200 418490 164400
rect 419262 163200 419318 164400
rect 420090 163200 420146 164400
rect 420918 163200 420974 164400
rect 421392 163254 421696 163282
rect 415872 163146 415900 163200
rect 415780 163118 415900 163146
rect 415860 159996 415912 160002
rect 415860 159938 415912 159944
rect 415216 152992 415268 152998
rect 415216 152934 415268 152940
rect 415400 152992 415452 152998
rect 415400 152934 415452 152940
rect 415228 150226 415256 152934
rect 415872 152386 415900 159938
rect 416700 158982 416728 163200
rect 417240 159860 417292 159866
rect 417240 159802 417292 159808
rect 416688 158976 416740 158982
rect 416688 158918 416740 158924
rect 417148 154488 417200 154494
rect 417148 154430 417200 154436
rect 416504 153060 416556 153066
rect 416504 153002 416556 153008
rect 415860 152380 415912 152386
rect 415860 152322 415912 152328
rect 415860 151836 415912 151842
rect 415860 151778 415912 151784
rect 415872 150226 415900 151778
rect 416516 150226 416544 153002
rect 417160 150226 417188 154430
rect 417252 151978 417280 159802
rect 417528 159662 417556 163200
rect 417516 159656 417568 159662
rect 417516 159598 417568 159604
rect 418448 157334 418476 163200
rect 418448 157306 418568 157334
rect 417884 152312 417936 152318
rect 417882 152280 417884 152289
rect 417936 152280 417938 152289
rect 417792 152244 417844 152250
rect 417882 152215 417938 152224
rect 417792 152186 417844 152192
rect 417240 151972 417292 151978
rect 417240 151914 417292 151920
rect 417804 150226 417832 152186
rect 418436 152040 418488 152046
rect 418436 151982 418488 151988
rect 408788 150198 408862 150226
rect 409432 150198 409506 150226
rect 410076 150198 410150 150226
rect 410720 150198 410794 150226
rect 411364 150198 411438 150226
rect 412008 150198 412082 150226
rect 412652 150198 412726 150226
rect 413296 150198 413370 150226
rect 413940 150198 414014 150226
rect 414584 150198 414658 150226
rect 415228 150198 415302 150226
rect 415872 150198 415946 150226
rect 416516 150198 416590 150226
rect 417160 150198 417234 150226
rect 417804 150198 417878 150226
rect 406856 150062 406930 150090
rect 407500 150062 407574 150090
rect 408144 150062 408218 150090
rect 406902 149940 406930 150062
rect 407546 149940 407574 150062
rect 408190 149940 408218 150062
rect 408834 149940 408862 150198
rect 409478 149940 409506 150198
rect 410122 149940 410150 150198
rect 410766 149940 410794 150198
rect 411410 149940 411438 150198
rect 412054 149940 412082 150198
rect 412698 149940 412726 150198
rect 413342 149940 413370 150198
rect 413986 149940 414014 150198
rect 414630 149940 414658 150198
rect 415274 149940 415302 150198
rect 415918 149940 415946 150198
rect 416562 149940 416590 150198
rect 417206 149940 417234 150198
rect 417850 149940 417878 150198
rect 418448 150090 418476 151982
rect 418540 151910 418568 157306
rect 419276 153066 419304 163200
rect 419632 159792 419684 159798
rect 419632 159734 419684 159740
rect 419540 158976 419592 158982
rect 419540 158918 419592 158924
rect 419264 153060 419316 153066
rect 419264 153002 419316 153008
rect 419552 152590 419580 158918
rect 419080 152584 419132 152590
rect 419080 152526 419132 152532
rect 419540 152584 419592 152590
rect 419540 152526 419592 152532
rect 418528 151904 418580 151910
rect 418528 151846 418580 151852
rect 419092 150090 419120 152526
rect 419644 152046 419672 159734
rect 420104 158982 420132 163200
rect 420932 159798 420960 163200
rect 420920 159792 420972 159798
rect 420920 159734 420972 159740
rect 420092 158976 420144 158982
rect 420092 158918 420144 158924
rect 419724 154352 419776 154358
rect 419724 154294 419776 154300
rect 419632 152040 419684 152046
rect 419632 151982 419684 151988
rect 419736 150090 419764 154294
rect 421012 153128 421064 153134
rect 421012 153070 421064 153076
rect 420368 152652 420420 152658
rect 420368 152594 420420 152600
rect 419816 152584 419868 152590
rect 419816 152526 419868 152532
rect 419828 152250 419856 152526
rect 419908 152312 419960 152318
rect 419906 152280 419908 152289
rect 419960 152280 419962 152289
rect 419816 152244 419868 152250
rect 419906 152215 419962 152224
rect 419816 152186 419868 152192
rect 420380 150090 420408 152594
rect 421024 152590 421052 153070
rect 421392 152658 421420 163254
rect 421668 163146 421696 163254
rect 421746 163200 421802 164400
rect 422574 163200 422630 164400
rect 423402 163200 423458 164400
rect 424322 163200 424378 164400
rect 425150 163200 425206 164400
rect 425256 163254 425928 163282
rect 421760 163146 421788 163200
rect 421668 163118 421788 163146
rect 422300 154420 422352 154426
rect 422300 154362 422352 154368
rect 421380 152652 421432 152658
rect 421380 152594 421432 152600
rect 421012 152584 421064 152590
rect 421012 152526 421064 152532
rect 421748 152244 421800 152250
rect 421748 152186 421800 152192
rect 421012 152108 421064 152114
rect 421012 152050 421064 152056
rect 421024 150090 421052 152050
rect 421760 151842 421788 152186
rect 421656 151836 421708 151842
rect 421656 151778 421708 151784
rect 421748 151836 421800 151842
rect 421748 151778 421800 151784
rect 421668 150090 421696 151778
rect 422312 150090 422340 154362
rect 422588 153134 422616 163200
rect 422852 153876 422904 153882
rect 422852 153818 422904 153824
rect 422576 153128 422628 153134
rect 422576 153070 422628 153076
rect 422864 150226 422892 153818
rect 422944 152788 422996 152794
rect 422944 152730 422996 152736
rect 422956 152250 422984 152730
rect 423416 152590 423444 163200
rect 424336 159526 424364 163200
rect 425164 161474 425192 163200
rect 425072 161446 425192 161474
rect 424876 160064 424928 160070
rect 424876 160006 424928 160012
rect 424324 159520 424376 159526
rect 424324 159462 424376 159468
rect 423588 158976 423640 158982
rect 423588 158918 423640 158924
rect 423600 153202 423628 158918
rect 423496 153196 423548 153202
rect 423496 153138 423548 153144
rect 423588 153196 423640 153202
rect 423588 153138 423640 153144
rect 423508 152794 423536 153138
rect 424232 152856 424284 152862
rect 424232 152798 424284 152804
rect 423496 152788 423548 152794
rect 423496 152730 423548 152736
rect 423312 152584 423364 152590
rect 423312 152526 423364 152532
rect 423404 152584 423456 152590
rect 423404 152526 423456 152532
rect 423324 152402 423352 152526
rect 423324 152374 423720 152402
rect 422944 152244 422996 152250
rect 422944 152186 422996 152192
rect 423692 152182 423720 152374
rect 423588 152176 423640 152182
rect 423588 152118 423640 152124
rect 423680 152176 423732 152182
rect 423680 152118 423732 152124
rect 422864 150198 423030 150226
rect 418448 150062 418522 150090
rect 419092 150062 419166 150090
rect 419736 150062 419810 150090
rect 420380 150062 420454 150090
rect 421024 150062 421098 150090
rect 421668 150062 421742 150090
rect 422312 150062 422386 150090
rect 418494 149940 418522 150062
rect 419138 149940 419166 150062
rect 419782 149940 419810 150062
rect 420426 149940 420454 150062
rect 421070 149940 421098 150062
rect 421714 149940 421742 150062
rect 422358 149940 422386 150062
rect 423002 149940 423030 150198
rect 423600 150090 423628 152118
rect 424244 150090 424272 152798
rect 424888 150226 424916 160006
rect 425072 152046 425100 161446
rect 425256 152794 425284 163254
rect 425900 163146 425928 163254
rect 425978 163200 426034 164400
rect 426452 163254 426756 163282
rect 425992 163146 426020 163200
rect 425900 163118 426020 163146
rect 425520 153944 425572 153950
rect 425520 153886 425572 153892
rect 425244 152788 425296 152794
rect 425244 152730 425296 152736
rect 425060 152040 425112 152046
rect 425060 151982 425112 151988
rect 424888 150198 424962 150226
rect 423600 150062 423674 150090
rect 424244 150062 424318 150090
rect 423646 149940 423674 150062
rect 424290 149940 424318 150062
rect 424934 149940 424962 150198
rect 425532 150090 425560 153886
rect 426452 152862 426480 163254
rect 426728 163146 426756 163254
rect 426806 163200 426862 164400
rect 427634 163200 427690 164400
rect 427832 163254 428412 163282
rect 426820 163146 426848 163200
rect 426728 163118 426848 163146
rect 427648 159458 427676 163200
rect 427360 159452 427412 159458
rect 427360 159394 427412 159400
rect 427636 159452 427688 159458
rect 427636 159394 427688 159400
rect 426164 152856 426216 152862
rect 426164 152798 426216 152804
rect 426440 152856 426492 152862
rect 426440 152798 426492 152804
rect 426176 150090 426204 152798
rect 426808 152380 426860 152386
rect 426808 152322 426860 152328
rect 426900 152380 426952 152386
rect 426900 152322 426952 152328
rect 426820 150090 426848 152322
rect 426912 151910 426940 152322
rect 427084 152176 427136 152182
rect 427084 152118 427136 152124
rect 426900 151904 426952 151910
rect 426900 151846 426952 151852
rect 427096 151842 427124 152118
rect 427084 151836 427136 151842
rect 427084 151778 427136 151784
rect 427372 150226 427400 159394
rect 427832 152182 427860 163254
rect 428384 163146 428412 163254
rect 428462 163200 428518 164400
rect 429290 163200 429346 164400
rect 430210 163200 430266 164400
rect 430592 163254 430988 163282
rect 428476 163146 428504 163200
rect 428384 163118 428504 163146
rect 428004 152720 428056 152726
rect 428004 152662 428056 152668
rect 427820 152176 427872 152182
rect 427820 152118 427872 152124
rect 428016 150226 428044 152662
rect 429304 152318 429332 163200
rect 429936 159724 429988 159730
rect 429936 159666 429988 159672
rect 429476 153128 429528 153134
rect 429476 153070 429528 153076
rect 428648 152312 428700 152318
rect 428648 152254 428700 152260
rect 429292 152312 429344 152318
rect 429292 152254 429344 152260
rect 428660 150226 428688 152254
rect 429488 152250 429516 153070
rect 429384 152244 429436 152250
rect 429384 152186 429436 152192
rect 429476 152244 429528 152250
rect 429476 152186 429528 152192
rect 429396 150226 429424 152186
rect 427372 150198 427446 150226
rect 428016 150198 428090 150226
rect 428660 150198 428734 150226
rect 425532 150062 425606 150090
rect 426176 150062 426250 150090
rect 426820 150062 426894 150090
rect 425578 149940 425606 150062
rect 426222 149940 426250 150062
rect 426866 149940 426894 150062
rect 427418 149940 427446 150198
rect 428062 149940 428090 150198
rect 428706 149940 428734 150198
rect 429350 150198 429424 150226
rect 429948 150226 429976 159666
rect 430224 153202 430252 163200
rect 430212 153196 430264 153202
rect 430212 153138 430264 153144
rect 430592 152726 430620 163254
rect 430960 163146 430988 163254
rect 431038 163200 431094 164400
rect 431236 163254 431816 163282
rect 431052 163146 431080 163200
rect 430960 163118 431080 163146
rect 430580 152720 430632 152726
rect 430580 152662 430632 152668
rect 431236 152561 431264 163254
rect 431788 163146 431816 163254
rect 431866 163200 431922 164400
rect 431972 163254 432644 163282
rect 431880 163146 431908 163200
rect 431788 163118 431908 163146
rect 431972 153134 432000 163254
rect 432616 163146 432644 163254
rect 432694 163200 432750 164400
rect 433522 163200 433578 164400
rect 434350 163200 434406 164400
rect 434732 163254 435128 163282
rect 432708 163146 432736 163200
rect 432616 163118 432736 163146
rect 432512 159588 432564 159594
rect 432512 159530 432564 159536
rect 431868 153128 431920 153134
rect 431868 153070 431920 153076
rect 431960 153128 432012 153134
rect 431960 153070 432012 153076
rect 431222 152552 431278 152561
rect 431222 152487 431278 152496
rect 430578 152416 430634 152425
rect 430578 152351 430634 152360
rect 430592 150226 430620 152351
rect 431880 151978 431908 153070
rect 432052 152380 432104 152386
rect 432052 152322 432104 152328
rect 432064 152250 432092 152322
rect 431960 152244 432012 152250
rect 431960 152186 432012 152192
rect 432052 152244 432104 152250
rect 432052 152186 432104 152192
rect 431776 151972 431828 151978
rect 431776 151914 431828 151920
rect 431868 151972 431920 151978
rect 431868 151914 431920 151920
rect 431224 151836 431276 151842
rect 431788 151814 431816 151914
rect 431972 151842 432000 152186
rect 431960 151836 432012 151842
rect 431788 151786 431908 151814
rect 431224 151778 431276 151784
rect 431236 150226 431264 151778
rect 431880 150226 431908 151786
rect 431960 151778 432012 151784
rect 432524 150226 432552 159530
rect 433536 152930 433564 163200
rect 433156 152924 433208 152930
rect 433156 152866 433208 152872
rect 433524 152924 433576 152930
rect 433524 152866 433576 152872
rect 433168 150226 433196 152866
rect 434364 152794 434392 163200
rect 434732 154358 434760 163254
rect 435100 163146 435128 163254
rect 435178 163200 435234 164400
rect 436098 163200 436154 164400
rect 436926 163200 436982 164400
rect 437492 163254 437704 163282
rect 435192 163146 435220 163200
rect 435100 163118 435220 163146
rect 435088 159384 435140 159390
rect 435088 159326 435140 159332
rect 434720 154352 434772 154358
rect 434720 154294 434772 154300
rect 434628 153060 434680 153066
rect 434628 153002 434680 153008
rect 434260 152788 434312 152794
rect 434260 152730 434312 152736
rect 434352 152788 434404 152794
rect 434352 152730 434404 152736
rect 434272 152658 434300 152730
rect 434260 152652 434312 152658
rect 434260 152594 434312 152600
rect 434640 152386 434668 153002
rect 433800 152380 433852 152386
rect 433800 152322 433852 152328
rect 434536 152380 434588 152386
rect 434536 152322 434588 152328
rect 434628 152380 434680 152386
rect 434628 152322 434680 152328
rect 433812 150226 433840 152322
rect 434548 152266 434576 152322
rect 434548 152238 434760 152266
rect 434732 152114 434760 152238
rect 434444 152108 434496 152114
rect 434444 152050 434496 152056
rect 434720 152108 434772 152114
rect 434720 152050 434772 152056
rect 434456 150226 434484 152050
rect 435100 150226 435128 159326
rect 436112 153066 436140 163200
rect 436940 161474 436968 163200
rect 436940 161446 437152 161474
rect 436100 153060 436152 153066
rect 436100 153002 436152 153008
rect 436376 152992 436428 152998
rect 436376 152934 436428 152940
rect 435732 152108 435784 152114
rect 435732 152050 435784 152056
rect 435744 150226 435772 152050
rect 436388 150226 436416 152934
rect 436928 152652 436980 152658
rect 436928 152594 436980 152600
rect 437020 152652 437072 152658
rect 437020 152594 437072 152600
rect 436836 152176 436888 152182
rect 436836 152118 436888 152124
rect 436848 152046 436876 152118
rect 436940 152046 436968 152594
rect 437032 152386 437060 152594
rect 437020 152380 437072 152386
rect 437020 152322 437072 152328
rect 436836 152040 436888 152046
rect 436836 151982 436888 151988
rect 436928 152040 436980 152046
rect 436928 151982 436980 151988
rect 437124 151910 437152 161446
rect 437492 152998 437520 163254
rect 437676 163146 437704 163254
rect 437754 163200 437810 164400
rect 437860 163254 438532 163282
rect 437768 163146 437796 163200
rect 437676 163118 437796 163146
rect 437664 159656 437716 159662
rect 437664 159598 437716 159604
rect 437480 152992 437532 152998
rect 437480 152934 437532 152940
rect 437020 151904 437072 151910
rect 437020 151846 437072 151852
rect 437112 151904 437164 151910
rect 437112 151846 437164 151852
rect 437032 150226 437060 151846
rect 437676 150226 437704 159598
rect 437860 153066 437888 163254
rect 438504 163146 438532 163254
rect 438582 163200 438638 164400
rect 438872 163254 439360 163282
rect 438596 163146 438624 163200
rect 438504 163118 438624 163146
rect 437756 153060 437808 153066
rect 437756 153002 437808 153008
rect 437848 153060 437900 153066
rect 437848 153002 437900 153008
rect 437768 152386 437796 153002
rect 438872 152386 438900 163254
rect 439332 163146 439360 163254
rect 439410 163200 439466 164400
rect 440238 163200 440294 164400
rect 440344 163254 441016 163282
rect 439424 163146 439452 163200
rect 439332 163118 439452 163146
rect 440252 152862 440280 163200
rect 440148 152856 440200 152862
rect 440148 152798 440200 152804
rect 440240 152856 440292 152862
rect 440240 152798 440292 152804
rect 438952 152652 439004 152658
rect 438952 152594 439004 152600
rect 437756 152380 437808 152386
rect 437756 152322 437808 152328
rect 438860 152380 438912 152386
rect 438860 152322 438912 152328
rect 438400 152312 438452 152318
rect 438584 152312 438636 152318
rect 438452 152260 438584 152266
rect 438400 152254 438636 152260
rect 438308 152244 438360 152250
rect 438412 152238 438624 152254
rect 438308 152186 438360 152192
rect 429948 150198 430022 150226
rect 430592 150198 430666 150226
rect 431236 150198 431310 150226
rect 431880 150198 431954 150226
rect 432524 150198 432598 150226
rect 433168 150198 433242 150226
rect 433812 150198 433886 150226
rect 434456 150198 434530 150226
rect 435100 150198 435174 150226
rect 435744 150198 435818 150226
rect 436388 150198 436462 150226
rect 437032 150198 437106 150226
rect 437676 150198 437750 150226
rect 429350 149940 429378 150198
rect 429994 149940 430022 150198
rect 430638 149940 430666 150198
rect 431282 149940 431310 150198
rect 431926 149940 431954 150198
rect 432570 149940 432598 150198
rect 433214 149940 433242 150198
rect 433858 149940 433886 150198
rect 434502 149940 434530 150198
rect 435146 149940 435174 150198
rect 435790 149940 435818 150198
rect 436434 149940 436462 150198
rect 437078 149940 437106 150198
rect 437722 149940 437750 150198
rect 438320 150090 438348 152186
rect 438964 150090 438992 152594
rect 440160 151978 440188 152798
rect 440344 152658 440372 163254
rect 440988 163146 441016 163254
rect 441066 163200 441122 164400
rect 441632 163254 441936 163282
rect 441080 163146 441108 163200
rect 440988 163118 441108 163146
rect 440424 159792 440476 159798
rect 440424 159734 440476 159740
rect 440332 152652 440384 152658
rect 440332 152594 440384 152600
rect 439596 151972 439648 151978
rect 439596 151914 439648 151920
rect 440148 151972 440200 151978
rect 440148 151914 440200 151920
rect 439608 150090 439636 151914
rect 440436 150226 440464 159734
rect 440884 152584 440936 152590
rect 440884 152526 440936 152532
rect 440298 150198 440464 150226
rect 438320 150062 438394 150090
rect 438964 150062 439038 150090
rect 439608 150062 439682 150090
rect 438366 149940 438394 150062
rect 439010 149940 439038 150062
rect 439654 149940 439682 150062
rect 440298 149940 440326 150198
rect 440896 150090 440924 152526
rect 441632 152250 441660 163254
rect 441908 163146 441936 163254
rect 441986 163200 442042 164400
rect 442092 163254 442764 163282
rect 442000 163146 442028 163200
rect 441908 163118 442028 163146
rect 441988 153128 442040 153134
rect 441988 153070 442040 153076
rect 441896 152992 441948 152998
rect 441894 152960 441896 152969
rect 441948 152960 441950 152969
rect 441894 152895 441950 152904
rect 441436 152244 441488 152250
rect 441436 152186 441488 152192
rect 441620 152244 441672 152250
rect 441620 152186 441672 152192
rect 441448 151706 441476 152186
rect 442000 151842 442028 153070
rect 442092 152590 442120 163254
rect 442736 163146 442764 163254
rect 442814 163200 442870 164400
rect 443012 163254 443592 163282
rect 442828 163146 442856 163200
rect 442736 163118 442856 163146
rect 442816 159520 442868 159526
rect 442816 159462 442868 159468
rect 442172 153128 442224 153134
rect 442172 153070 442224 153076
rect 442184 152946 442212 153070
rect 442540 152992 442592 152998
rect 442538 152960 442540 152969
rect 442592 152960 442594 152969
rect 442184 152918 442488 152946
rect 442460 152862 442488 152918
rect 442538 152895 442594 152904
rect 442448 152856 442500 152862
rect 442448 152798 442500 152804
rect 442080 152584 442132 152590
rect 442080 152526 442132 152532
rect 442172 152448 442224 152454
rect 442172 152390 442224 152396
rect 441528 151836 441580 151842
rect 441528 151778 441580 151784
rect 441988 151836 442040 151842
rect 441988 151778 442040 151784
rect 441436 151700 441488 151706
rect 441436 151642 441488 151648
rect 441540 150090 441568 151778
rect 442184 150090 442212 152390
rect 442828 150226 442856 159462
rect 443012 152930 443040 163254
rect 443564 163146 443592 163254
rect 443642 163200 443698 164400
rect 444470 163200 444526 164400
rect 445298 163200 445354 164400
rect 446126 163200 446182 164400
rect 446324 163254 446904 163282
rect 443656 163146 443684 163200
rect 443564 163118 443684 163146
rect 444288 154352 444340 154358
rect 444288 154294 444340 154300
rect 443000 152924 443052 152930
rect 443000 152866 443052 152872
rect 444196 152380 444248 152386
rect 443840 152340 444196 152368
rect 443460 152176 443512 152182
rect 443460 152118 443512 152124
rect 442828 150198 442902 150226
rect 440896 150062 440970 150090
rect 441540 150062 441614 150090
rect 442184 150062 442258 150090
rect 440942 149940 440970 150062
rect 441586 149940 441614 150062
rect 442230 149940 442258 150062
rect 442874 149940 442902 150198
rect 443472 150090 443500 152118
rect 443840 151910 443868 152340
rect 444196 152322 444248 152328
rect 444104 152040 444156 152046
rect 444104 151982 444156 151988
rect 443828 151904 443880 151910
rect 443828 151846 443880 151852
rect 444116 150226 444144 151982
rect 444300 151978 444328 154294
rect 444380 152856 444432 152862
rect 444380 152798 444432 152804
rect 444392 152386 444420 152798
rect 444380 152380 444432 152386
rect 444380 152322 444432 152328
rect 444380 152108 444432 152114
rect 444380 152050 444432 152056
rect 444288 151972 444340 151978
rect 444288 151914 444340 151920
rect 444392 151842 444420 152050
rect 444484 152046 444512 163200
rect 445312 152182 445340 163200
rect 446140 159866 446168 163200
rect 446128 159860 446180 159866
rect 446128 159802 446180 159808
rect 445392 159452 445444 159458
rect 445392 159394 445444 159400
rect 445208 152176 445260 152182
rect 445208 152118 445260 152124
rect 445300 152176 445352 152182
rect 445300 152118 445352 152124
rect 444472 152040 444524 152046
rect 444472 151982 444524 151988
rect 444472 151904 444524 151910
rect 444472 151846 444524 151852
rect 444380 151836 444432 151842
rect 444380 151778 444432 151784
rect 444484 150226 444512 151846
rect 445220 151842 445248 152118
rect 445208 151836 445260 151842
rect 445208 151778 445260 151784
rect 445404 150226 445432 159394
rect 446324 152862 446352 163254
rect 446876 163146 446904 163254
rect 446954 163200 447010 164400
rect 447874 163200 447930 164400
rect 448702 163200 448758 164400
rect 449530 163200 449586 164400
rect 450358 163200 450414 164400
rect 451186 163200 451242 164400
rect 452014 163200 452070 164400
rect 452842 163200 452898 164400
rect 453762 163200 453818 164400
rect 454590 163200 454646 164400
rect 455418 163200 455474 164400
rect 456246 163200 456302 164400
rect 457074 163200 457130 164400
rect 457902 163200 457958 164400
rect 458730 163200 458786 164400
rect 459650 163200 459706 164400
rect 460478 163200 460534 164400
rect 461306 163200 461362 164400
rect 462134 163200 462190 164400
rect 462962 163200 463018 164400
rect 463790 163200 463846 164400
rect 464618 163200 464674 164400
rect 465538 163200 465594 164400
rect 466366 163200 466422 164400
rect 467194 163200 467250 164400
rect 468022 163200 468078 164400
rect 468850 163200 468906 164400
rect 469678 163200 469734 164400
rect 470506 163200 470562 164400
rect 471426 163200 471482 164400
rect 472254 163200 472310 164400
rect 473082 163200 473138 164400
rect 473910 163200 473966 164400
rect 474738 163200 474794 164400
rect 475566 163200 475622 164400
rect 476394 163200 476450 164400
rect 477314 163200 477370 164400
rect 478142 163200 478198 164400
rect 478970 163200 479026 164400
rect 479798 163200 479854 164400
rect 480626 163200 480682 164400
rect 481454 163200 481510 164400
rect 482282 163200 482338 164400
rect 483202 163200 483258 164400
rect 484030 163200 484086 164400
rect 484412 163254 484808 163282
rect 446968 163146 446996 163200
rect 446876 163118 446996 163146
rect 447888 159526 447916 163200
rect 448716 159798 448744 163200
rect 448704 159792 448756 159798
rect 448704 159734 448756 159740
rect 447876 159520 447928 159526
rect 447876 159462 447928 159468
rect 449544 159458 449572 163200
rect 449532 159452 449584 159458
rect 449532 159394 449584 159400
rect 450372 159390 450400 163200
rect 451200 159730 451228 163200
rect 451188 159724 451240 159730
rect 451188 159666 451240 159672
rect 452028 159594 452056 163200
rect 452016 159588 452068 159594
rect 452016 159530 452068 159536
rect 450360 159384 450412 159390
rect 450360 159326 450412 159332
rect 452856 158778 452884 163200
rect 453776 159662 453804 163200
rect 453764 159656 453816 159662
rect 453764 159598 453816 159604
rect 454604 158914 454632 163200
rect 454592 158908 454644 158914
rect 454592 158850 454644 158856
rect 455432 158846 455460 163200
rect 456260 158982 456288 163200
rect 457088 159934 457116 163200
rect 457076 159928 457128 159934
rect 457076 159870 457128 159876
rect 456800 159860 456852 159866
rect 456800 159802 456852 159808
rect 456248 158976 456300 158982
rect 456248 158918 456300 158924
rect 455420 158840 455472 158846
rect 455420 158782 455472 158788
rect 452844 158772 452896 158778
rect 452844 158714 452896 158720
rect 456812 153202 456840 159802
rect 457916 159118 457944 163200
rect 458744 159866 458772 163200
rect 458732 159860 458784 159866
rect 458732 159802 458784 159808
rect 459664 159254 459692 163200
rect 460112 159520 460164 159526
rect 460112 159462 460164 159468
rect 459652 159248 459704 159254
rect 459652 159190 459704 159196
rect 457904 159112 457956 159118
rect 457904 159054 457956 159060
rect 459560 158772 459612 158778
rect 459560 158714 459612 158720
rect 447324 153196 447376 153202
rect 447324 153138 447376 153144
rect 456800 153196 456852 153202
rect 456800 153138 456852 153144
rect 459468 153196 459520 153202
rect 459468 153138 459520 153144
rect 446312 152856 446364 152862
rect 446312 152798 446364 152804
rect 446680 152312 446732 152318
rect 446680 152254 446732 152260
rect 446036 151836 446088 151842
rect 446036 151778 446088 151784
rect 444116 150198 444190 150226
rect 444484 150198 444834 150226
rect 445404 150198 445478 150226
rect 443472 150062 443546 150090
rect 443518 149940 443546 150062
rect 444162 149940 444190 150198
rect 444806 149940 444834 150198
rect 445450 149940 445478 150198
rect 446048 150090 446076 151778
rect 446692 150090 446720 152254
rect 447336 150226 447364 153138
rect 449900 153128 449952 153134
rect 449900 153070 449952 153076
rect 447968 152720 448020 152726
rect 447968 152662 448020 152668
rect 447980 150226 448008 152662
rect 448610 152552 448666 152561
rect 448610 152487 448666 152496
rect 448624 150226 448652 152487
rect 449256 152108 449308 152114
rect 449256 152050 449308 152056
rect 449268 150226 449296 152050
rect 449912 150226 449940 153070
rect 455052 153060 455104 153066
rect 455052 153002 455104 153008
rect 453120 152992 453172 152998
rect 453120 152934 453172 152940
rect 451188 152924 451240 152930
rect 451188 152866 451240 152872
rect 450544 152788 450596 152794
rect 450544 152730 450596 152736
rect 450556 150226 450584 152730
rect 451200 151978 451228 152866
rect 452476 152448 452528 152454
rect 452476 152390 452528 152396
rect 451096 151972 451148 151978
rect 451096 151914 451148 151920
rect 451188 151972 451240 151978
rect 451188 151914 451240 151920
rect 451108 151814 451136 151914
rect 451832 151904 451884 151910
rect 451832 151846 451884 151852
rect 451108 151786 451228 151814
rect 451200 150226 451228 151786
rect 451844 150226 451872 151846
rect 452488 150226 452516 152390
rect 453132 150226 453160 152934
rect 454408 152516 454460 152522
rect 454408 152458 454460 152464
rect 453764 152380 453816 152386
rect 453764 152322 453816 152328
rect 453776 150226 453804 152322
rect 454420 150226 454448 152458
rect 455064 150226 455092 153002
rect 455696 152652 455748 152658
rect 455696 152594 455748 152600
rect 455708 150226 455736 152594
rect 456984 152584 457036 152590
rect 456984 152526 457036 152532
rect 456340 152244 456392 152250
rect 456340 152186 456392 152192
rect 456352 150226 456380 152186
rect 456996 150226 457024 152526
rect 458824 152176 458876 152182
rect 458824 152118 458876 152124
rect 458180 152040 458232 152046
rect 458180 151982 458232 151988
rect 457628 151972 457680 151978
rect 457628 151914 457680 151920
rect 457640 150226 457668 151914
rect 458192 150226 458220 151982
rect 458836 150226 458864 152118
rect 459480 150226 459508 153138
rect 459572 152590 459600 158714
rect 460020 152856 460072 152862
rect 460020 152798 460072 152804
rect 459560 152584 459612 152590
rect 459560 152526 459612 152532
rect 460032 150498 460060 152798
rect 460124 151814 460152 159462
rect 460492 159050 460520 163200
rect 460940 159792 460992 159798
rect 460940 159734 460992 159740
rect 460480 159044 460532 159050
rect 460480 158986 460532 158992
rect 460952 151814 460980 159734
rect 461320 159526 461348 163200
rect 461308 159520 461360 159526
rect 461308 159462 461360 159468
rect 461492 159452 461544 159458
rect 461492 159394 461544 159400
rect 461504 151814 461532 159394
rect 462148 159322 462176 163200
rect 462320 159724 462372 159730
rect 462320 159666 462372 159672
rect 462136 159316 462188 159322
rect 462136 159258 462188 159264
rect 461676 158908 461728 158914
rect 461676 158850 461728 158856
rect 461688 153202 461716 158850
rect 461676 153196 461728 153202
rect 461676 153138 461728 153144
rect 460124 151786 460796 151814
rect 460952 151786 461440 151814
rect 461504 151786 462084 151814
rect 460032 150470 460152 150498
rect 460124 150226 460152 150470
rect 460768 150226 460796 151786
rect 461412 150226 461440 151786
rect 462056 150226 462084 151786
rect 447336 150198 447410 150226
rect 447980 150198 448054 150226
rect 448624 150198 448698 150226
rect 449268 150198 449342 150226
rect 449912 150198 449986 150226
rect 450556 150198 450630 150226
rect 451200 150198 451274 150226
rect 451844 150198 451918 150226
rect 452488 150198 452562 150226
rect 453132 150198 453206 150226
rect 453776 150198 453850 150226
rect 454420 150198 454494 150226
rect 455064 150198 455138 150226
rect 455708 150198 455782 150226
rect 456352 150198 456426 150226
rect 456996 150198 457070 150226
rect 457640 150198 457714 150226
rect 458192 150198 458266 150226
rect 458836 150198 458910 150226
rect 459480 150198 459554 150226
rect 460124 150198 460198 150226
rect 460768 150198 460842 150226
rect 461412 150198 461486 150226
rect 462056 150198 462130 150226
rect 462332 150210 462360 159666
rect 462688 159384 462740 159390
rect 462688 159326 462740 159332
rect 462700 150226 462728 159326
rect 462976 159186 463004 163200
rect 462964 159180 463016 159186
rect 462964 159122 463016 159128
rect 463148 158976 463200 158982
rect 463148 158918 463200 158924
rect 463160 153066 463188 158918
rect 463608 158840 463660 158846
rect 463608 158782 463660 158788
rect 463620 153134 463648 158782
rect 463804 158778 463832 163200
rect 464344 159928 464396 159934
rect 464344 159870 464396 159876
rect 463976 159588 464028 159594
rect 463976 159530 464028 159536
rect 463792 158772 463844 158778
rect 463792 158714 463844 158720
rect 463608 153128 463660 153134
rect 463608 153070 463660 153076
rect 463148 153060 463200 153066
rect 463148 153002 463200 153008
rect 463988 150226 464016 159530
rect 464356 151910 464384 159870
rect 464528 159112 464580 159118
rect 464528 159054 464580 159060
rect 464540 152998 464568 159054
rect 464632 158846 464660 163200
rect 465080 159860 465132 159866
rect 465080 159802 465132 159808
rect 464620 158840 464672 158846
rect 464620 158782 464672 158788
rect 464528 152992 464580 152998
rect 464528 152934 464580 152940
rect 465092 152930 465120 159802
rect 465264 159656 465316 159662
rect 465264 159598 465316 159604
rect 465080 152924 465132 152930
rect 465080 152866 465132 152872
rect 464620 152584 464672 152590
rect 464620 152526 464672 152532
rect 464344 151904 464396 151910
rect 464344 151846 464396 151852
rect 464632 150226 464660 152526
rect 465276 150226 465304 159598
rect 465552 158914 465580 163200
rect 466380 158982 466408 163200
rect 467208 159594 467236 163200
rect 468036 159730 468064 163200
rect 468024 159724 468076 159730
rect 468024 159666 468076 159672
rect 467196 159588 467248 159594
rect 467196 159530 467248 159536
rect 467932 159520 467984 159526
rect 467932 159462 467984 159468
rect 467840 159316 467892 159322
rect 467840 159258 467892 159264
rect 466644 159248 466696 159254
rect 466644 159190 466696 159196
rect 466460 159044 466512 159050
rect 466460 158986 466512 158992
rect 466368 158976 466420 158982
rect 466368 158918 466420 158924
rect 465540 158908 465592 158914
rect 465540 158850 465592 158856
rect 466472 153202 466500 158986
rect 465908 153196 465960 153202
rect 465908 153138 465960 153144
rect 466460 153196 466512 153202
rect 466460 153138 466512 153144
rect 465920 150226 465948 153138
rect 466656 153134 466684 159190
rect 466552 153128 466604 153134
rect 466552 153070 466604 153076
rect 466644 153128 466696 153134
rect 466644 153070 466696 153076
rect 466564 150226 466592 153070
rect 467196 153060 467248 153066
rect 467196 153002 467248 153008
rect 467208 150226 467236 153002
rect 467852 152046 467880 159258
rect 467840 152040 467892 152046
rect 467840 151982 467892 151988
rect 467944 151910 467972 159462
rect 468864 159458 468892 163200
rect 469692 159798 469720 163200
rect 469680 159792 469732 159798
rect 469680 159734 469732 159740
rect 468852 159452 468904 159458
rect 468852 159394 468904 159400
rect 470520 159390 470548 163200
rect 470508 159384 470560 159390
rect 470508 159326 470560 159332
rect 469220 159180 469272 159186
rect 469220 159122 469272 159128
rect 468392 152992 468444 152998
rect 468392 152934 468444 152940
rect 467840 151904 467892 151910
rect 467840 151846 467892 151852
rect 467932 151904 467984 151910
rect 467932 151846 467984 151852
rect 467852 150226 467880 151846
rect 468404 151814 468432 152934
rect 469128 152924 469180 152930
rect 469128 152866 469180 152872
rect 468404 151786 468524 151814
rect 468496 150226 468524 151786
rect 469140 150226 469168 152866
rect 469232 151978 469260 159122
rect 471440 159118 471468 163200
rect 472268 159866 472296 163200
rect 472256 159860 472308 159866
rect 472256 159802 472308 159808
rect 471428 159112 471480 159118
rect 471428 159054 471480 159060
rect 472348 158976 472400 158982
rect 472348 158918 472400 158924
rect 472164 158908 472216 158914
rect 472164 158850 472216 158856
rect 471428 158840 471480 158846
rect 471428 158782 471480 158788
rect 470416 153196 470468 153202
rect 470416 153138 470468 153144
rect 469772 153128 469824 153134
rect 469772 153070 469824 153076
rect 469220 151972 469272 151978
rect 469220 151914 469272 151920
rect 469784 150226 469812 153070
rect 470428 150226 470456 153138
rect 471440 153134 471468 158782
rect 471796 158772 471848 158778
rect 471796 158714 471848 158720
rect 471808 153202 471836 158714
rect 471796 153196 471848 153202
rect 471796 153138 471848 153144
rect 471428 153128 471480 153134
rect 471428 153070 471480 153076
rect 472176 153066 472204 158850
rect 472164 153060 472216 153066
rect 472164 153002 472216 153008
rect 472360 152998 472388 158918
rect 473096 158778 473124 163200
rect 473360 159588 473412 159594
rect 473360 159530 473412 159536
rect 473084 158772 473136 158778
rect 473084 158714 473136 158720
rect 473372 153202 473400 159530
rect 473924 159050 473952 163200
rect 473912 159044 473964 159050
rect 473912 158986 473964 158992
rect 474752 158914 474780 163200
rect 474832 159452 474884 159458
rect 474832 159394 474884 159400
rect 474740 158908 474792 158914
rect 474740 158850 474792 158856
rect 472992 153196 473044 153202
rect 472992 153138 473044 153144
rect 473360 153196 473412 153202
rect 473360 153138 473412 153144
rect 472348 152992 472400 152998
rect 472348 152934 472400 152940
rect 471704 152040 471756 152046
rect 471704 151982 471756 151988
rect 471060 151904 471112 151910
rect 471060 151846 471112 151852
rect 471072 150226 471100 151846
rect 471716 150226 471744 151982
rect 472348 151972 472400 151978
rect 472348 151914 472400 151920
rect 472360 150226 472388 151914
rect 473004 150226 473032 153138
rect 474844 153134 474872 159394
rect 475580 158982 475608 163200
rect 476028 159724 476080 159730
rect 476028 159666 476080 159672
rect 475568 158976 475620 158982
rect 475568 158918 475620 158924
rect 475568 153196 475620 153202
rect 475568 153138 475620 153144
rect 473636 153128 473688 153134
rect 473636 153070 473688 153076
rect 474832 153128 474884 153134
rect 474832 153070 474884 153076
rect 473648 150226 473676 153070
rect 474280 153060 474332 153066
rect 474280 153002 474332 153008
rect 474292 150226 474320 153002
rect 474924 152992 474976 152998
rect 474924 152934 474976 152940
rect 474936 150226 474964 152934
rect 475580 150226 475608 153138
rect 476040 151814 476068 159666
rect 476120 159384 476172 159390
rect 476120 159326 476172 159332
rect 476132 153202 476160 159326
rect 476408 158846 476436 163200
rect 477328 159458 477356 163200
rect 477408 159792 477460 159798
rect 477408 159734 477460 159740
rect 477316 159452 477368 159458
rect 477316 159394 477368 159400
rect 476396 158840 476448 158846
rect 476396 158782 476448 158788
rect 476120 153196 476172 153202
rect 476120 153138 476172 153144
rect 476856 153128 476908 153134
rect 476856 153070 476908 153076
rect 476040 151786 476252 151814
rect 476224 150226 476252 151786
rect 476868 150226 476896 153070
rect 477420 151814 477448 159734
rect 478156 159390 478184 163200
rect 478984 159798 479012 163200
rect 479432 159860 479484 159866
rect 479432 159802 479484 159808
rect 478972 159792 479024 159798
rect 478972 159734 479024 159740
rect 478144 159384 478196 159390
rect 478144 159326 478196 159332
rect 477684 159112 477736 159118
rect 477684 159054 477736 159060
rect 477420 151786 477540 151814
rect 477512 150226 477540 151786
rect 446048 150062 446122 150090
rect 446692 150062 446766 150090
rect 446094 149940 446122 150062
rect 446738 149940 446766 150062
rect 447382 149940 447410 150198
rect 448026 149940 448054 150198
rect 448670 149940 448698 150198
rect 449314 149940 449342 150198
rect 449958 149940 449986 150198
rect 450602 149940 450630 150198
rect 451246 149940 451274 150198
rect 451890 149940 451918 150198
rect 452534 149940 452562 150198
rect 453178 149940 453206 150198
rect 453822 149940 453850 150198
rect 454466 149940 454494 150198
rect 455110 149940 455138 150198
rect 455754 149940 455782 150198
rect 456398 149940 456426 150198
rect 457042 149940 457070 150198
rect 457686 149940 457714 150198
rect 458238 149940 458266 150198
rect 458882 149940 458910 150198
rect 459526 149940 459554 150198
rect 460170 149940 460198 150198
rect 460814 149940 460842 150198
rect 461458 149940 461486 150198
rect 462102 149940 462130 150198
rect 462320 150204 462372 150210
rect 462700 150198 462774 150226
rect 462320 150146 462372 150152
rect 462746 149940 462774 150198
rect 463378 150204 463430 150210
rect 463988 150198 464062 150226
rect 464632 150198 464706 150226
rect 465276 150198 465350 150226
rect 465920 150198 465994 150226
rect 466564 150198 466638 150226
rect 467208 150198 467282 150226
rect 467852 150198 467926 150226
rect 468496 150198 468570 150226
rect 469140 150198 469214 150226
rect 469784 150198 469858 150226
rect 470428 150198 470502 150226
rect 471072 150198 471146 150226
rect 471716 150198 471790 150226
rect 472360 150198 472434 150226
rect 473004 150198 473078 150226
rect 473648 150198 473722 150226
rect 474292 150198 474366 150226
rect 474936 150198 475010 150226
rect 475580 150198 475654 150226
rect 476224 150198 476298 150226
rect 476868 150198 476942 150226
rect 477512 150198 477586 150226
rect 477696 150210 477724 159054
rect 478972 158772 479024 158778
rect 478972 158714 479024 158720
rect 478144 153196 478196 153202
rect 478144 153138 478196 153144
rect 478156 150226 478184 153138
rect 463378 150146 463430 150152
rect 463390 149940 463418 150146
rect 464034 149940 464062 150198
rect 464678 149940 464706 150198
rect 465322 149940 465350 150198
rect 465966 149940 465994 150198
rect 466610 149940 466638 150198
rect 467254 149940 467282 150198
rect 467898 149940 467926 150198
rect 468542 149940 468570 150198
rect 469186 149940 469214 150198
rect 469830 149940 469858 150198
rect 470474 149940 470502 150198
rect 471118 149940 471146 150198
rect 471762 149940 471790 150198
rect 472406 149940 472434 150198
rect 473050 149940 473078 150198
rect 473694 149940 473722 150198
rect 474338 149940 474366 150198
rect 474982 149940 475010 150198
rect 475626 149940 475654 150198
rect 476270 149940 476298 150198
rect 476914 149940 476942 150198
rect 477558 149940 477586 150198
rect 477684 150204 477736 150210
rect 478156 150198 478230 150226
rect 478984 150210 479012 158714
rect 479444 150226 479472 159802
rect 479812 159730 479840 163200
rect 480640 159934 480668 163200
rect 480628 159928 480680 159934
rect 480628 159870 480680 159876
rect 479800 159724 479852 159730
rect 479800 159666 479852 159672
rect 481468 159526 481496 163200
rect 481456 159520 481508 159526
rect 481456 159462 481508 159468
rect 480260 159044 480312 159050
rect 480260 158986 480312 158992
rect 480272 151814 480300 158986
rect 482008 158976 482060 158982
rect 482008 158918 482060 158924
rect 481364 158908 481416 158914
rect 481364 158850 481416 158856
rect 480272 151786 480760 151814
rect 480732 150226 480760 151786
rect 481376 150226 481404 158850
rect 481640 158840 481692 158846
rect 481640 158782 481692 158788
rect 477684 150146 477736 150152
rect 478202 149940 478230 150198
rect 478834 150204 478886 150210
rect 478834 150146 478886 150152
rect 478972 150204 479024 150210
rect 479444 150198 479518 150226
rect 478972 150146 479024 150152
rect 478846 149940 478874 150146
rect 479490 149940 479518 150198
rect 480122 150204 480174 150210
rect 480732 150198 480806 150226
rect 481376 150198 481450 150226
rect 481652 150210 481680 158782
rect 482020 150226 482048 158918
rect 482296 158778 482324 163200
rect 483216 161474 483244 163200
rect 483124 161446 483244 161474
rect 482284 158772 482336 158778
rect 482284 158714 482336 158720
rect 483124 152998 483152 161446
rect 483296 159452 483348 159458
rect 483296 159394 483348 159400
rect 483204 159384 483256 159390
rect 483204 159326 483256 159332
rect 483112 152992 483164 152998
rect 483112 152934 483164 152940
rect 480122 150146 480174 150152
rect 480134 149940 480162 150146
rect 480778 149940 480806 150198
rect 481422 149940 481450 150198
rect 481640 150204 481692 150210
rect 482020 150198 482094 150226
rect 483216 150210 483244 159326
rect 483308 150226 483336 159394
rect 484044 153202 484072 163200
rect 484032 153196 484084 153202
rect 484032 153138 484084 153144
rect 484412 153066 484440 163254
rect 484780 163146 484808 163254
rect 484858 163200 484914 164400
rect 484964 163254 485636 163282
rect 484872 163146 484900 163200
rect 484780 163118 484900 163146
rect 484676 159792 484728 159798
rect 484676 159734 484728 159740
rect 484400 153060 484452 153066
rect 484400 153002 484452 153008
rect 484688 150226 484716 159734
rect 484964 153134 484992 163254
rect 485608 163146 485636 163254
rect 485686 163200 485742 164400
rect 485792 163254 486464 163282
rect 485700 163146 485728 163200
rect 485608 163118 485728 163146
rect 485228 159724 485280 159730
rect 485228 159666 485280 159672
rect 484952 153128 485004 153134
rect 484952 153070 485004 153076
rect 481640 150146 481692 150152
rect 482066 149940 482094 150198
rect 482698 150204 482750 150210
rect 482698 150146 482750 150152
rect 483204 150204 483256 150210
rect 483308 150198 483382 150226
rect 483204 150146 483256 150152
rect 482710 149940 482738 150146
rect 483354 149940 483382 150198
rect 483986 150204 484038 150210
rect 483986 150146 484038 150152
rect 484642 150198 484716 150226
rect 485240 150226 485268 159666
rect 485792 152046 485820 163254
rect 486436 163146 486464 163254
rect 486514 163200 486570 164400
rect 487342 163200 487398 164400
rect 488170 163200 488226 164400
rect 488552 163254 489040 163282
rect 486528 163146 486556 163200
rect 486436 163118 486556 163146
rect 485964 159928 486016 159934
rect 485964 159870 486016 159876
rect 485780 152040 485832 152046
rect 485780 151982 485832 151988
rect 485976 150226 486004 159870
rect 486516 159520 486568 159526
rect 486516 159462 486568 159468
rect 485240 150198 485314 150226
rect 483998 149940 484026 150146
rect 484642 149940 484670 150198
rect 485286 149940 485314 150198
rect 485930 150198 486004 150226
rect 486528 150226 486556 159462
rect 487252 158772 487304 158778
rect 487252 158714 487304 158720
rect 487264 150226 487292 158714
rect 487356 151978 487384 163200
rect 487804 152992 487856 152998
rect 487804 152934 487856 152940
rect 487344 151972 487396 151978
rect 487344 151914 487396 151920
rect 486528 150198 486602 150226
rect 485930 149940 485958 150198
rect 486574 149940 486602 150198
rect 487218 150198 487292 150226
rect 487816 150226 487844 152934
rect 488184 151842 488212 163200
rect 488448 153196 488500 153202
rect 488448 153138 488500 153144
rect 488172 151836 488224 151842
rect 488172 151778 488224 151784
rect 488460 150226 488488 153138
rect 488552 151910 488580 163254
rect 489012 163146 489040 163254
rect 489090 163200 489146 164400
rect 489918 163200 489974 164400
rect 490024 163254 490696 163282
rect 489104 163146 489132 163200
rect 489012 163118 489132 163146
rect 489932 153202 489960 163200
rect 489920 153196 489972 153202
rect 489920 153138 489972 153144
rect 489644 153128 489696 153134
rect 489644 153070 489696 153076
rect 489000 153060 489052 153066
rect 489000 153002 489052 153008
rect 488540 151904 488592 151910
rect 488540 151846 488592 151852
rect 489012 150226 489040 153002
rect 489656 150226 489684 153070
rect 490024 152930 490052 163254
rect 490668 163146 490696 163254
rect 490746 163200 490802 164400
rect 491312 163254 491524 163282
rect 490760 163146 490788 163200
rect 490668 163118 490788 163146
rect 491312 152998 491340 163254
rect 491496 163146 491524 163254
rect 491574 163200 491630 164400
rect 491680 163254 492352 163282
rect 491588 163146 491616 163200
rect 491496 163118 491616 163146
rect 491680 153134 491708 163254
rect 492324 163146 492352 163254
rect 492402 163200 492458 164400
rect 492692 163254 493180 163282
rect 492416 163146 492444 163200
rect 492324 163118 492444 163146
rect 491668 153128 491720 153134
rect 491668 153070 491720 153076
rect 492692 153066 492720 163254
rect 493152 163146 493180 163254
rect 493230 163200 493286 164400
rect 494058 163200 494114 164400
rect 494978 163200 495034 164400
rect 495544 163254 495756 163282
rect 493244 163146 493272 163200
rect 493152 163118 493272 163146
rect 494072 153202 494100 163200
rect 492864 153196 492916 153202
rect 492864 153138 492916 153144
rect 494060 153196 494112 153202
rect 494060 153138 494112 153144
rect 492680 153060 492732 153066
rect 492680 153002 492732 153008
rect 491300 152992 491352 152998
rect 491300 152934 491352 152940
rect 490012 152924 490064 152930
rect 490012 152866 490064 152872
rect 490288 152040 490340 152046
rect 490288 151982 490340 151988
rect 490300 150226 490328 151982
rect 490932 151972 490984 151978
rect 490932 151914 490984 151920
rect 490944 150226 490972 151914
rect 492220 151904 492272 151910
rect 492220 151846 492272 151852
rect 491576 151836 491628 151842
rect 491576 151778 491628 151784
rect 491588 150226 491616 151778
rect 492232 150226 492260 151846
rect 492876 150226 492904 153138
rect 494992 153134 495020 163200
rect 494796 153128 494848 153134
rect 494796 153070 494848 153076
rect 494980 153128 495032 153134
rect 494980 153070 495032 153076
rect 494152 152992 494204 152998
rect 494152 152934 494204 152940
rect 493508 152924 493560 152930
rect 493508 152866 493560 152872
rect 493520 150226 493548 152866
rect 494164 150226 494192 152934
rect 494808 150226 494836 153070
rect 495544 153066 495572 163254
rect 495728 163146 495756 163254
rect 495806 163200 495862 164400
rect 496634 163200 496690 164400
rect 496832 163254 497412 163282
rect 495820 163146 495848 163200
rect 495728 163118 495848 163146
rect 496648 153202 496676 163200
rect 496084 153196 496136 153202
rect 496084 153138 496136 153144
rect 496636 153196 496688 153202
rect 496636 153138 496688 153144
rect 495440 153060 495492 153066
rect 495440 153002 495492 153008
rect 495532 153060 495584 153066
rect 495532 153002 495584 153008
rect 495452 150226 495480 153002
rect 496096 150226 496124 153138
rect 496832 153134 496860 163254
rect 497384 163146 497412 163254
rect 497462 163200 497518 164400
rect 498290 163200 498346 164400
rect 499118 163200 499174 164400
rect 499946 163200 500002 164400
rect 500052 163254 500632 163282
rect 497476 163146 497504 163200
rect 497384 163118 497504 163146
rect 498304 156670 498332 163200
rect 498292 156664 498344 156670
rect 498292 156606 498344 156612
rect 498016 153196 498068 153202
rect 498016 153138 498068 153144
rect 496728 153128 496780 153134
rect 496728 153070 496780 153076
rect 496820 153128 496872 153134
rect 496820 153070 496872 153076
rect 496740 150226 496768 153070
rect 497372 153060 497424 153066
rect 497372 153002 497424 153008
rect 497384 150226 497412 153002
rect 498028 150226 498056 153138
rect 498660 153128 498712 153134
rect 498660 153070 498712 153076
rect 498672 150226 498700 153070
rect 499132 151842 499160 163200
rect 499960 163146 499988 163200
rect 500052 163146 500080 163254
rect 499960 163118 500080 163146
rect 499304 156664 499356 156670
rect 499304 156606 499356 156612
rect 499120 151836 499172 151842
rect 499120 151778 499172 151784
rect 499316 150226 499344 156606
rect 499948 151836 500000 151842
rect 499948 151778 500000 151784
rect 499960 150226 499988 151778
rect 500604 150226 500632 163254
rect 500866 163200 500922 164400
rect 501694 163200 501750 164400
rect 502522 163200 502578 164400
rect 503350 163200 503406 164400
rect 503824 163254 504128 163282
rect 500880 151814 500908 163200
rect 501708 161474 501736 163200
rect 501708 161446 501920 161474
rect 500880 151786 501276 151814
rect 501248 150226 501276 151786
rect 501892 150226 501920 161446
rect 502536 150226 502564 163200
rect 503364 151814 503392 163200
rect 503272 151786 503392 151814
rect 503272 150226 503300 151786
rect 487816 150198 487890 150226
rect 488460 150198 488534 150226
rect 489012 150198 489086 150226
rect 489656 150198 489730 150226
rect 490300 150198 490374 150226
rect 490944 150198 491018 150226
rect 491588 150198 491662 150226
rect 492232 150198 492306 150226
rect 492876 150198 492950 150226
rect 493520 150198 493594 150226
rect 494164 150198 494238 150226
rect 494808 150198 494882 150226
rect 495452 150198 495526 150226
rect 496096 150198 496170 150226
rect 496740 150198 496814 150226
rect 497384 150198 497458 150226
rect 498028 150198 498102 150226
rect 498672 150198 498746 150226
rect 499316 150198 499390 150226
rect 499960 150198 500034 150226
rect 500604 150198 500678 150226
rect 501248 150198 501322 150226
rect 501892 150198 501966 150226
rect 502536 150198 502610 150226
rect 487218 149940 487246 150198
rect 487862 149940 487890 150198
rect 488506 149940 488534 150198
rect 489058 149940 489086 150198
rect 489702 149940 489730 150198
rect 490346 149940 490374 150198
rect 490990 149940 491018 150198
rect 491634 149940 491662 150198
rect 492278 149940 492306 150198
rect 492922 149940 492950 150198
rect 493566 149940 493594 150198
rect 494210 149940 494238 150198
rect 494854 149940 494882 150198
rect 495498 149940 495526 150198
rect 496142 149940 496170 150198
rect 496786 149940 496814 150198
rect 497430 149940 497458 150198
rect 498074 149940 498102 150198
rect 498718 149940 498746 150198
rect 499362 149940 499390 150198
rect 500006 149940 500034 150198
rect 500650 149940 500678 150198
rect 501294 149940 501322 150198
rect 501938 149940 501966 150198
rect 502582 149940 502610 150198
rect 503226 150198 503300 150226
rect 503824 150226 503852 163254
rect 504100 163146 504128 163254
rect 504178 163200 504234 164400
rect 504468 163254 504956 163282
rect 504192 163146 504220 163200
rect 504100 163118 504220 163146
rect 504468 150226 504496 163254
rect 504928 163146 504956 163254
rect 505006 163200 505062 164400
rect 505112 163254 505784 163282
rect 505020 163146 505048 163200
rect 504928 163118 505048 163146
rect 505112 150226 505140 163254
rect 505756 163146 505784 163254
rect 505834 163200 505890 164400
rect 506754 163200 506810 164400
rect 507582 163200 507638 164400
rect 508410 163200 508466 164400
rect 509238 163200 509294 164400
rect 509344 163254 509556 163282
rect 505848 163146 505876 163200
rect 505756 163118 505876 163146
rect 506388 158840 506440 158846
rect 506388 158782 506440 158788
rect 505284 158772 505336 158778
rect 505284 158714 505336 158720
rect 505296 151814 505324 158714
rect 505296 151786 505784 151814
rect 505756 150226 505784 151786
rect 506400 150226 506428 158782
rect 506768 158778 506796 163200
rect 507596 158846 507624 163200
rect 508320 158908 508372 158914
rect 508320 158850 508372 158856
rect 507584 158840 507636 158846
rect 507584 158782 507636 158788
rect 506756 158772 506808 158778
rect 506756 158714 506808 158720
rect 507032 158772 507084 158778
rect 507032 158714 507084 158720
rect 507044 150226 507072 158714
rect 507768 151904 507820 151910
rect 507768 151846 507820 151852
rect 507780 150226 507808 151846
rect 503824 150198 503898 150226
rect 504468 150198 504542 150226
rect 505112 150198 505186 150226
rect 505756 150198 505830 150226
rect 506400 150198 506474 150226
rect 507044 150198 507118 150226
rect 503226 149940 503254 150198
rect 503870 149940 503898 150198
rect 504514 149940 504542 150198
rect 505158 149940 505186 150198
rect 505802 149940 505830 150198
rect 506446 149940 506474 150198
rect 507090 149940 507118 150198
rect 507734 150198 507808 150226
rect 508332 150226 508360 158850
rect 508424 158778 508452 163200
rect 509252 163146 509280 163200
rect 509344 163146 509372 163254
rect 509252 163118 509372 163146
rect 508412 158772 508464 158778
rect 508412 158714 508464 158720
rect 509424 158772 509476 158778
rect 509424 158714 509476 158720
rect 509056 151972 509108 151978
rect 509056 151914 509108 151920
rect 509068 150226 509096 151914
rect 509436 151814 509464 158714
rect 509528 151910 509556 163254
rect 510066 163200 510122 164400
rect 510894 163200 510950 164400
rect 511722 163200 511778 164400
rect 512012 163254 512592 163282
rect 510080 158914 510108 163200
rect 510068 158908 510120 158914
rect 510068 158850 510120 158856
rect 510344 152856 510396 152862
rect 510344 152798 510396 152804
rect 509516 151904 509568 151910
rect 509516 151846 509568 151852
rect 509436 151786 509648 151814
rect 508332 150198 508406 150226
rect 507734 149940 507762 150198
rect 508378 149940 508406 150198
rect 509022 150198 509096 150226
rect 509620 150226 509648 151786
rect 510356 150226 510384 152798
rect 510908 151978 510936 163200
rect 511736 158778 511764 163200
rect 511724 158772 511776 158778
rect 511724 158714 511776 158720
rect 510988 153196 511040 153202
rect 510988 153138 511040 153144
rect 510896 151972 510948 151978
rect 510896 151914 510948 151920
rect 511000 150226 511028 153138
rect 512012 152862 512040 163254
rect 512564 163146 512592 163254
rect 512642 163200 512698 164400
rect 513470 163200 513526 164400
rect 513576 163254 514248 163282
rect 512656 163146 512684 163200
rect 512564 163118 512684 163146
rect 513484 153202 513512 163200
rect 513472 153196 513524 153202
rect 513472 153138 513524 153144
rect 512920 153128 512972 153134
rect 512920 153070 512972 153076
rect 512276 152992 512328 152998
rect 512276 152934 512328 152940
rect 512000 152856 512052 152862
rect 512000 152798 512052 152804
rect 511632 152380 511684 152386
rect 511632 152322 511684 152328
rect 511644 150226 511672 152322
rect 512288 150226 512316 152934
rect 512932 150226 512960 153070
rect 513576 152386 513604 163254
rect 514220 163146 514248 163254
rect 514298 163200 514354 164400
rect 514772 163254 515076 163282
rect 514312 163146 514340 163200
rect 514220 163118 514340 163146
rect 514208 153196 514260 153202
rect 514208 153138 514260 153144
rect 513564 152380 513616 152386
rect 513564 152322 513616 152328
rect 513564 152244 513616 152250
rect 513564 152186 513616 152192
rect 513576 150226 513604 152186
rect 514220 150226 514248 153138
rect 514772 152998 514800 163254
rect 515048 163146 515076 163254
rect 515126 163200 515182 164400
rect 515232 163254 515904 163282
rect 515140 163146 515168 163200
rect 515048 163118 515168 163146
rect 514944 158772 514996 158778
rect 514944 158714 514996 158720
rect 514760 152992 514812 152998
rect 514760 152934 514812 152940
rect 514956 151814 514984 158714
rect 515232 153134 515260 163254
rect 515876 163146 515904 163254
rect 515954 163200 516010 164400
rect 516152 163254 516732 163282
rect 515968 163146 515996 163200
rect 515876 163118 515996 163146
rect 515220 153128 515272 153134
rect 515220 153070 515272 153076
rect 516152 152250 516180 163254
rect 516704 163146 516732 163254
rect 516782 163200 516838 164400
rect 517610 163200 517666 164400
rect 518530 163200 518586 164400
rect 518912 163254 519308 163282
rect 516796 163146 516824 163200
rect 516704 163118 516824 163146
rect 517624 161474 517652 163200
rect 517532 161446 517652 161474
rect 517532 158794 517560 161446
rect 517440 158766 517560 158794
rect 518544 158778 518572 163200
rect 518808 159520 518860 159526
rect 518808 159462 518860 159468
rect 518716 159384 518768 159390
rect 518716 159326 518768 159332
rect 518532 158772 518584 158778
rect 517440 153202 517468 158766
rect 518532 158714 518584 158720
rect 517428 153196 517480 153202
rect 517428 153138 517480 153144
rect 516140 152244 516192 152250
rect 516140 152186 516192 152192
rect 516692 152040 516744 152046
rect 516692 151982 516744 151988
rect 515496 151972 515548 151978
rect 515496 151914 515548 151920
rect 514864 151786 514984 151814
rect 514864 150226 514892 151786
rect 515508 150226 515536 151914
rect 516048 151904 516100 151910
rect 516048 151846 516100 151852
rect 509620 150198 509694 150226
rect 509022 149940 509050 150198
rect 509666 149940 509694 150198
rect 510310 150198 510384 150226
rect 510954 150198 511028 150226
rect 511598 150198 511672 150226
rect 512242 150198 512316 150226
rect 512886 150198 512960 150226
rect 513530 150198 513604 150226
rect 514174 150198 514248 150226
rect 514818 150198 514892 150226
rect 515462 150198 515536 150226
rect 516060 150226 516088 151846
rect 516704 150226 516732 151982
rect 517428 151836 517480 151842
rect 517428 151778 517480 151784
rect 517440 150226 517468 151778
rect 518728 150226 518756 159326
rect 516060 150198 516134 150226
rect 516704 150198 516778 150226
rect 510310 149940 510338 150198
rect 510954 149940 510982 150198
rect 511598 149940 511626 150198
rect 512242 149940 512270 150198
rect 512886 149940 512914 150198
rect 513530 149940 513558 150198
rect 514174 149940 514202 150198
rect 514818 149940 514846 150198
rect 515462 149940 515490 150198
rect 516106 149940 516134 150198
rect 516750 149940 516778 150198
rect 517394 150198 517468 150226
rect 518026 150204 518078 150210
rect 517394 149940 517422 150198
rect 518026 150146 518078 150152
rect 518682 150198 518756 150226
rect 518820 150210 518848 159462
rect 518912 151978 518940 163254
rect 519280 163146 519308 163254
rect 519358 163200 519414 164400
rect 519464 163254 520136 163282
rect 519372 163146 519400 163200
rect 519280 163118 519400 163146
rect 519358 157176 519414 157185
rect 519358 157111 519414 157120
rect 518900 151972 518952 151978
rect 518900 151914 518952 151920
rect 518808 150204 518860 150210
rect 518038 149940 518066 150146
rect 518682 149940 518710 150198
rect 518808 150146 518860 150152
rect 519372 143857 519400 157111
rect 519464 151910 519492 163254
rect 519726 163160 519782 163169
rect 520108 163146 520136 163254
rect 520186 163200 520242 164400
rect 520292 163254 520964 163282
rect 520200 163146 520228 163200
rect 520108 163118 520228 163146
rect 519726 163095 519782 163104
rect 519542 161664 519598 161673
rect 519542 161599 519598 161608
rect 519452 151904 519504 151910
rect 519452 151846 519504 151852
rect 519556 147937 519584 161599
rect 519634 160168 519690 160177
rect 519634 160103 519690 160112
rect 519542 147928 519598 147937
rect 519542 147863 519598 147872
rect 519648 146577 519676 160103
rect 519740 149297 519768 163095
rect 520002 158672 520058 158681
rect 520002 158607 520058 158616
rect 519818 151192 519874 151201
rect 519818 151127 519874 151136
rect 519726 149288 519782 149297
rect 519726 149223 519782 149232
rect 519726 148200 519782 148209
rect 519726 148135 519782 148144
rect 519634 146568 519690 146577
rect 519634 146503 519690 146512
rect 519634 145072 519690 145081
rect 519634 145007 519690 145016
rect 519358 143848 519414 143857
rect 519358 143783 519414 143792
rect 519542 142216 519598 142225
rect 519542 142151 519598 142160
rect 519450 140584 519506 140593
rect 519450 140519 519506 140528
rect 519266 139088 519322 139097
rect 519266 139023 519322 139032
rect 519280 127537 519308 139023
rect 519358 137592 519414 137601
rect 519358 137527 519414 137536
rect 519266 127528 519322 127537
rect 519266 127463 519322 127472
rect 519372 126177 519400 137527
rect 519464 128897 519492 140519
rect 519556 130257 519584 142151
rect 519648 132977 519676 145007
rect 519740 135697 519768 148135
rect 519832 138417 519860 151127
rect 519910 149696 519966 149705
rect 519910 149631 519966 149640
rect 519818 138408 519874 138417
rect 519818 138343 519874 138352
rect 519924 137057 519952 149631
rect 520016 145217 520044 158607
rect 520094 155680 520150 155689
rect 520094 155615 520150 155624
rect 520002 145208 520058 145217
rect 520002 145143 520058 145152
rect 520108 142497 520136 155615
rect 520186 154184 520242 154193
rect 520186 154119 520242 154128
rect 520094 142488 520150 142497
rect 520094 142423 520150 142432
rect 520200 141137 520228 154119
rect 520292 152046 520320 163254
rect 520936 163146 520964 163254
rect 521014 163200 521070 164400
rect 521842 163200 521898 164400
rect 522670 163200 522726 164400
rect 523498 163200 523554 164400
rect 521028 163146 521056 163200
rect 520936 163118 521056 163146
rect 521856 161474 521884 163200
rect 521672 161446 521884 161474
rect 521672 158794 521700 161446
rect 522684 159526 522712 163200
rect 522672 159520 522724 159526
rect 522672 159462 522724 159468
rect 523512 159390 523540 163200
rect 523500 159384 523552 159390
rect 523500 159326 523552 159332
rect 521580 158766 521700 158794
rect 521106 152688 521162 152697
rect 521106 152623 521162 152632
rect 520280 152040 520332 152046
rect 520280 151982 520332 151988
rect 521014 146704 521070 146713
rect 521014 146639 521070 146648
rect 520922 143712 520978 143721
rect 520922 143647 520978 143656
rect 520186 141128 520242 141137
rect 520186 141063 520242 141072
rect 519910 137048 519966 137057
rect 519910 136983 519966 136992
rect 519910 136096 519966 136105
rect 519910 136031 519966 136040
rect 519726 135688 519782 135697
rect 519726 135623 519782 135632
rect 519726 134600 519782 134609
rect 519726 134535 519782 134544
rect 519634 132968 519690 132977
rect 519634 132903 519690 132912
rect 519542 130248 519598 130257
rect 519542 130183 519598 130192
rect 519450 128888 519506 128897
rect 519450 128823 519506 128832
rect 519542 127120 519598 127129
rect 519542 127055 519598 127064
rect 519358 126168 519414 126177
rect 519358 126103 519414 126112
rect 519266 124128 519322 124137
rect 519266 124063 519322 124072
rect 519174 119640 519230 119649
rect 519174 119575 519230 119584
rect 117228 118040 117280 118046
rect 117228 117982 117280 117988
rect 519188 109857 519216 119575
rect 519280 113937 519308 124063
rect 519450 122632 519506 122641
rect 519450 122567 519506 122576
rect 519358 121136 519414 121145
rect 519358 121071 519414 121080
rect 519266 113928 519322 113937
rect 519266 113863 519322 113872
rect 519372 111217 519400 121071
rect 519464 112577 519492 122567
rect 519556 116657 519584 127055
rect 519634 125624 519690 125633
rect 519634 125559 519690 125568
rect 519542 116648 519598 116657
rect 519542 116583 519598 116592
rect 519648 115297 519676 125559
rect 519740 123457 519768 134535
rect 519818 128616 519874 128625
rect 519818 128551 519874 128560
rect 519726 123448 519782 123457
rect 519726 123383 519782 123392
rect 519832 118017 519860 128551
rect 519924 124817 519952 136031
rect 520002 133104 520058 133113
rect 520002 133039 520058 133048
rect 519910 124808 519966 124817
rect 519910 124743 519966 124752
rect 520016 122097 520044 133039
rect 520936 131753 520964 143647
rect 521028 134337 521056 146639
rect 521120 139777 521148 152623
rect 521580 151842 521608 158766
rect 521568 151836 521620 151842
rect 521568 151778 521620 151784
rect 521106 139768 521162 139777
rect 521106 139703 521162 139712
rect 521014 134328 521070 134337
rect 521014 134263 521070 134272
rect 520922 131744 520978 131753
rect 520922 131679 520978 131688
rect 520094 131608 520150 131617
rect 520094 131543 520150 131552
rect 520002 122088 520058 122097
rect 520002 122023 520058 122032
rect 520108 120737 520136 131543
rect 520186 130112 520242 130121
rect 520186 130047 520242 130056
rect 520094 120728 520150 120737
rect 520094 120663 520150 120672
rect 520200 119377 520228 130047
rect 520186 119368 520242 119377
rect 520186 119303 520242 119312
rect 520002 118144 520058 118153
rect 520002 118079 520058 118088
rect 519818 118008 519874 118017
rect 519818 117943 519874 117952
rect 519910 116512 519966 116521
rect 519910 116447 519966 116456
rect 519634 115288 519690 115297
rect 519634 115223 519690 115232
rect 519818 115016 519874 115025
rect 519818 114951 519874 114960
rect 519726 113520 519782 113529
rect 519726 113455 519782 113464
rect 519450 112568 519506 112577
rect 519450 112503 519506 112512
rect 519634 112024 519690 112033
rect 519634 111959 519690 111968
rect 519358 111208 519414 111217
rect 519358 111143 519414 111152
rect 519542 110528 519598 110537
rect 519542 110463 519598 110472
rect 519174 109848 519230 109857
rect 519174 109783 519230 109792
rect 117134 104816 117190 104825
rect 117134 104751 117190 104760
rect 117042 102912 117098 102921
rect 117042 102847 117098 102856
rect 519556 101697 519584 110463
rect 519648 103057 519676 111959
rect 519740 104417 519768 113455
rect 519832 105777 519860 114951
rect 519924 107137 519952 116447
rect 520016 108497 520044 118079
rect 521106 109032 521162 109041
rect 521106 108967 521162 108976
rect 520002 108488 520058 108497
rect 520002 108423 520058 108432
rect 520830 107536 520886 107545
rect 520830 107471 520886 107480
rect 519910 107128 519966 107137
rect 519910 107063 519966 107072
rect 520278 106040 520334 106049
rect 520278 105975 520334 105984
rect 519818 105768 519874 105777
rect 519818 105703 519874 105712
rect 519726 104408 519782 104417
rect 519726 104343 519782 104352
rect 519634 103048 519690 103057
rect 519634 102983 519690 102992
rect 519542 101688 519598 101697
rect 519542 101623 519598 101632
rect 116950 101008 117006 101017
rect 116950 100943 117006 100952
rect 116858 99104 116914 99113
rect 116858 99039 116914 99048
rect 520292 97617 520320 105975
rect 520738 103048 520794 103057
rect 520738 102983 520794 102992
rect 520278 97608 520334 97617
rect 520278 97543 520334 97552
rect 116766 97200 116822 97209
rect 116766 97135 116822 97144
rect 520278 95568 520334 95577
rect 520278 95503 520334 95512
rect 116674 95296 116730 95305
rect 116674 95231 116730 95240
rect 116582 93392 116638 93401
rect 116582 93327 116638 93336
rect 116124 92472 116176 92478
rect 116124 92414 116176 92420
rect 520186 92440 520242 92449
rect 116136 91361 116164 92414
rect 520186 92375 520242 92384
rect 116122 91352 116178 91361
rect 116122 91287 116178 91296
rect 520094 90944 520150 90953
rect 520094 90879 520150 90888
rect 116124 89684 116176 89690
rect 116124 89626 116176 89632
rect 116136 89457 116164 89626
rect 116122 89448 116178 89457
rect 116122 89383 116178 89392
rect 520002 89448 520058 89457
rect 520002 89383 520058 89392
rect 116032 88324 116084 88330
rect 116032 88266 116084 88272
rect 116044 87553 116072 88266
rect 519818 87952 519874 87961
rect 519818 87887 519874 87896
rect 116030 87544 116086 87553
rect 116030 87479 116086 87488
rect 116492 87236 116544 87242
rect 116492 87178 116544 87184
rect 115202 85640 115258 85649
rect 115202 85575 115258 85584
rect 116216 82816 116268 82822
rect 116216 82758 116268 82764
rect 116228 81841 116256 82758
rect 116214 81832 116270 81841
rect 116214 81767 116270 81776
rect 114100 80028 114152 80034
rect 114100 79970 114152 79976
rect 115940 80028 115992 80034
rect 115940 79970 115992 79976
rect 115952 79937 115980 79970
rect 115938 79928 115994 79937
rect 115938 79863 115994 79872
rect 116504 78033 116532 87178
rect 519634 86456 519690 86465
rect 519634 86391 519690 86400
rect 116584 83972 116636 83978
rect 116584 83914 116636 83920
rect 116596 83745 116624 83914
rect 116582 83736 116638 83745
rect 116582 83671 116638 83680
rect 519266 83464 519322 83473
rect 519266 83399 519322 83408
rect 116490 78024 116546 78033
rect 116490 77959 116546 77968
rect 519280 77217 519308 83399
rect 519542 81968 519598 81977
rect 519542 81903 519598 81912
rect 519450 80472 519506 80481
rect 519450 80407 519506 80416
rect 519266 77208 519322 77217
rect 519266 77143 519322 77152
rect 519464 74633 519492 80407
rect 519556 75993 519584 81903
rect 519648 79937 519676 86391
rect 519726 84960 519782 84969
rect 519726 84895 519782 84904
rect 519634 79928 519690 79937
rect 519634 79863 519690 79872
rect 519740 78577 519768 84895
rect 519832 81297 519860 87887
rect 520016 82657 520044 89383
rect 520108 84017 520136 90879
rect 520200 85377 520228 92375
rect 520292 88097 520320 95503
rect 520752 94897 520780 102983
rect 520844 98977 520872 107471
rect 521014 104544 521070 104553
rect 521014 104479 521070 104488
rect 520830 98968 520886 98977
rect 520830 98903 520886 98912
rect 521028 96257 521056 104479
rect 521120 100337 521148 108967
rect 521474 101552 521530 101561
rect 521474 101487 521530 101496
rect 521106 100328 521162 100337
rect 521106 100263 521162 100272
rect 521382 100056 521438 100065
rect 521382 99991 521438 100000
rect 521290 98560 521346 98569
rect 521290 98495 521346 98504
rect 521106 97064 521162 97073
rect 521106 96999 521162 97008
rect 521014 96248 521070 96257
rect 521014 96183 521070 96192
rect 520738 94888 520794 94897
rect 520738 94823 520794 94832
rect 520922 93936 520978 93945
rect 520922 93871 520978 93880
rect 520278 88088 520334 88097
rect 520278 88023 520334 88032
rect 520936 86737 520964 93871
rect 521120 89593 521148 96999
rect 521304 90817 521332 98495
rect 521396 92177 521424 99991
rect 521488 93537 521516 101487
rect 521474 93528 521530 93537
rect 521474 93463 521530 93472
rect 521382 92168 521438 92177
rect 521382 92103 521438 92112
rect 521290 90808 521346 90817
rect 521290 90743 521346 90752
rect 521106 89584 521162 89593
rect 521106 89519 521162 89528
rect 520922 86728 520978 86737
rect 520922 86663 520978 86672
rect 520186 85368 520242 85377
rect 520186 85303 520242 85312
rect 520094 84008 520150 84017
rect 520094 83943 520150 83952
rect 520002 82648 520058 82657
rect 520002 82583 520058 82592
rect 519818 81288 519874 81297
rect 519818 81223 519874 81232
rect 519910 78976 519966 78985
rect 519910 78911 519966 78920
rect 519726 78568 519782 78577
rect 519726 78503 519782 78512
rect 519818 77480 519874 77489
rect 519818 77415 519874 77424
rect 519542 75984 519598 75993
rect 519542 75919 519598 75928
rect 519726 75984 519782 75993
rect 519726 75919 519782 75928
rect 519450 74624 519506 74633
rect 519450 74559 519506 74568
rect 116674 74080 116730 74089
rect 116674 74015 116730 74024
rect 116582 72176 116638 72185
rect 116582 72111 116638 72120
rect 116596 71806 116624 72111
rect 114192 71800 114244 71806
rect 114192 71742 114244 71748
rect 116584 71800 116636 71806
rect 116584 71742 116636 71748
rect 114100 69080 114152 69086
rect 114100 69022 114152 69028
rect 114008 67652 114060 67658
rect 114008 67594 114060 67600
rect 113916 66292 113968 66298
rect 113916 66234 113968 66240
rect 113824 63572 113876 63578
rect 113824 63514 113876 63520
rect 109684 41472 109736 41478
rect 109684 41414 109736 41420
rect 53654 2680 53710 2689
rect 2516 2650 2714 2666
rect 2504 2644 2714 2650
rect 2556 2638 2714 2644
rect 39330 2650 39436 2666
rect 42642 2650 43024 2666
rect 46046 2650 46152 2666
rect 39330 2644 39448 2650
rect 39330 2638 39396 2644
rect 2504 2586 2556 2592
rect 39396 2586 39448 2592
rect 39764 2644 39816 2650
rect 42642 2644 43036 2650
rect 42642 2638 42984 2644
rect 39764 2586 39816 2592
rect 42984 2586 43036 2592
rect 43536 2644 43588 2650
rect 46046 2644 46164 2650
rect 46046 2638 46112 2644
rect 43536 2586 43588 2592
rect 46112 2586 46164 2592
rect 50620 2644 50672 2650
rect 83002 2680 83058 2689
rect 62698 2650 62896 2666
rect 53654 2615 53656 2624
rect 50620 2586 50672 2592
rect 53708 2615 53710 2624
rect 58716 2644 58768 2650
rect 53656 2586 53708 2592
rect 58716 2586 58768 2592
rect 58808 2644 58860 2650
rect 62698 2644 62908 2650
rect 62698 2638 62856 2644
rect 58808 2586 58860 2592
rect 62856 2586 62908 2592
rect 63316 2644 63368 2650
rect 63316 2586 63368 2592
rect 63500 2644 63552 2650
rect 63500 2586 63552 2592
rect 66996 2644 67048 2650
rect 66996 2586 67048 2592
rect 68008 2644 68060 2650
rect 68008 2586 68060 2592
rect 80152 2644 80204 2650
rect 80152 2586 80204 2592
rect 80244 2644 80296 2650
rect 80244 2586 80296 2592
rect 80336 2644 80388 2650
rect 80336 2586 80388 2592
rect 80428 2644 80480 2650
rect 80428 2586 80480 2592
rect 81532 2644 81584 2650
rect 81532 2586 81584 2592
rect 81624 2644 81676 2650
rect 81624 2586 81676 2592
rect 81808 2644 81860 2650
rect 81808 2586 81860 2592
rect 81900 2644 81952 2650
rect 81900 2586 81952 2592
rect 81992 2644 82044 2650
rect 81992 2586 82044 2592
rect 82452 2644 82504 2650
rect 82452 2586 82504 2592
rect 82728 2644 82780 2650
rect 83002 2615 83004 2624
rect 82728 2586 82780 2592
rect 83056 2615 83058 2624
rect 83096 2644 83148 2650
rect 83004 2586 83056 2592
rect 83096 2586 83148 2592
rect 98368 2644 98420 2650
rect 98368 2586 98420 2592
rect 98460 2644 98512 2650
rect 98460 2586 98512 2592
rect 100024 2644 100076 2650
rect 100024 2586 100076 2592
rect 32772 2508 32824 2514
rect 32772 2450 32824 2456
rect 6012 1426 6040 2108
rect 9324 1465 9352 2108
rect 12636 1601 12664 2108
rect 15948 1737 15976 2108
rect 19352 1873 19380 2108
rect 19338 1864 19394 1873
rect 19338 1799 19394 1808
rect 15934 1728 15990 1737
rect 15934 1663 15990 1672
rect 12622 1592 12678 1601
rect 12622 1527 12678 1536
rect 22664 1494 22692 2108
rect 25976 1562 26004 2108
rect 29288 1630 29316 2108
rect 32692 1698 32720 2108
rect 32680 1692 32732 1698
rect 32680 1634 32732 1640
rect 29276 1624 29328 1630
rect 29276 1566 29328 1572
rect 25964 1556 26016 1562
rect 25964 1498 26016 1504
rect 22652 1488 22704 1494
rect 9310 1456 9366 1465
rect 6000 1420 6052 1426
rect 22652 1430 22704 1436
rect 9310 1391 9366 1400
rect 6000 1362 6052 1368
rect 32784 800 32812 2450
rect 39776 2446 39804 2586
rect 43548 2514 43576 2586
rect 43536 2508 43588 2514
rect 43536 2450 43588 2456
rect 50632 2446 50660 2586
rect 58624 2576 58676 2582
rect 58728 2553 58756 2586
rect 58624 2518 58676 2524
rect 58714 2544 58770 2553
rect 58636 2446 58664 2518
rect 58714 2479 58770 2488
rect 36360 2440 36412 2446
rect 36018 2388 36360 2394
rect 36018 2382 36412 2388
rect 39764 2440 39816 2446
rect 39764 2382 39816 2388
rect 50620 2440 50672 2446
rect 56140 2440 56192 2446
rect 56138 2408 56140 2417
rect 58624 2440 58676 2446
rect 56192 2408 56194 2417
rect 50620 2382 50672 2388
rect 36018 2366 36400 2382
rect 52670 2378 52960 2394
rect 52670 2372 52972 2378
rect 52670 2366 52920 2372
rect 58624 2382 58676 2388
rect 56138 2343 56194 2352
rect 52920 2314 52972 2320
rect 58820 2310 58848 2586
rect 59728 2576 59780 2582
rect 59386 2524 59728 2530
rect 59386 2518 59780 2524
rect 59386 2502 59768 2518
rect 49608 2304 49660 2310
rect 49358 2252 49608 2258
rect 58808 2304 58860 2310
rect 49358 2246 49660 2252
rect 49358 2230 49648 2246
rect 55982 2242 56272 2258
rect 58808 2246 58860 2252
rect 55982 2236 56284 2242
rect 55982 2230 56232 2236
rect 56232 2178 56284 2184
rect 63328 2174 63356 2586
rect 63512 2417 63540 2586
rect 63498 2408 63554 2417
rect 66350 2408 66406 2417
rect 66010 2366 66350 2394
rect 63498 2343 63554 2352
rect 67008 2378 67036 2586
rect 68020 2446 68048 2586
rect 73252 2576 73304 2582
rect 73080 2524 73252 2530
rect 73080 2518 73304 2524
rect 73080 2514 73292 2518
rect 73068 2508 73292 2514
rect 73120 2502 73292 2508
rect 73344 2508 73396 2514
rect 73068 2450 73120 2456
rect 73344 2450 73396 2456
rect 68008 2440 68060 2446
rect 73356 2394 73384 2450
rect 80164 2446 80192 2586
rect 68008 2382 68060 2388
rect 69322 2378 69704 2394
rect 66350 2343 66406 2352
rect 66996 2372 67048 2378
rect 69322 2372 69716 2378
rect 69322 2366 69664 2372
rect 66996 2314 67048 2320
rect 69664 2314 69716 2320
rect 73080 2366 73384 2394
rect 80152 2440 80204 2446
rect 80152 2382 80204 2388
rect 73080 2242 73108 2366
rect 80256 2242 80284 2586
rect 73068 2236 73120 2242
rect 73068 2178 73120 2184
rect 80244 2236 80296 2242
rect 80244 2178 80296 2184
rect 80348 2174 80376 2586
rect 63316 2168 63368 2174
rect 63316 2110 63368 2116
rect 80336 2168 80388 2174
rect 80336 2110 80388 2116
rect 72712 1834 72740 2108
rect 72700 1828 72752 1834
rect 72700 1770 72752 1776
rect 76024 1766 76052 2108
rect 79336 1902 79364 2108
rect 80440 2106 80468 2586
rect 81544 2242 81572 2586
rect 81532 2236 81584 2242
rect 81532 2178 81584 2184
rect 81636 2106 81664 2586
rect 81820 2174 81848 2586
rect 81912 2446 81940 2586
rect 81900 2440 81952 2446
rect 81900 2382 81952 2388
rect 82004 2310 82032 2586
rect 82360 2576 82412 2582
rect 82082 2544 82138 2553
rect 82358 2544 82360 2553
rect 82412 2544 82414 2553
rect 82082 2479 82138 2488
rect 82268 2508 82320 2514
rect 81992 2304 82044 2310
rect 81992 2246 82044 2252
rect 82096 2242 82124 2479
rect 82358 2479 82414 2488
rect 82268 2450 82320 2456
rect 82280 2378 82308 2450
rect 82268 2372 82320 2378
rect 82268 2314 82320 2320
rect 82464 2242 82492 2586
rect 82740 2417 82768 2586
rect 83108 2553 83136 2586
rect 83094 2544 83150 2553
rect 98380 2514 98408 2586
rect 83094 2479 83150 2488
rect 98368 2508 98420 2514
rect 98368 2450 98420 2456
rect 82726 2408 82782 2417
rect 82726 2343 82782 2352
rect 96002 2242 96384 2258
rect 82084 2236 82136 2242
rect 82084 2178 82136 2184
rect 82452 2236 82504 2242
rect 96002 2236 96396 2242
rect 96002 2230 96344 2236
rect 82452 2178 82504 2184
rect 96344 2178 96396 2184
rect 81808 2168 81860 2174
rect 93032 2168 93084 2174
rect 81808 2110 81860 2116
rect 80428 2100 80480 2106
rect 80428 2042 80480 2048
rect 81624 2100 81676 2106
rect 81624 2042 81676 2048
rect 82648 1970 82676 2108
rect 86066 2094 86448 2122
rect 89378 2106 89668 2122
rect 92690 2116 93032 2122
rect 92690 2110 93084 2116
rect 89378 2100 89680 2106
rect 89378 2094 89628 2100
rect 86420 2038 86448 2094
rect 92690 2094 93072 2110
rect 89628 2042 89680 2048
rect 86408 2032 86460 2038
rect 86408 1974 86460 1980
rect 82636 1964 82688 1970
rect 82636 1906 82688 1912
rect 79324 1896 79376 1902
rect 79324 1838 79376 1844
rect 76012 1760 76064 1766
rect 76012 1702 76064 1708
rect 98472 1578 98500 2586
rect 100036 2514 100064 2586
rect 109342 2514 109632 2530
rect 100024 2508 100076 2514
rect 109342 2508 109644 2514
rect 109342 2502 109592 2508
rect 100024 2450 100076 2456
rect 109592 2450 109644 2456
rect 106188 2440 106240 2446
rect 102718 2378 103008 2394
rect 106030 2388 106188 2394
rect 106030 2382 106240 2388
rect 102718 2372 103020 2378
rect 102718 2366 102968 2372
rect 106030 2366 106228 2382
rect 102968 2314 103020 2320
rect 99656 2304 99708 2310
rect 99406 2252 99656 2258
rect 99406 2246 99708 2252
rect 99406 2230 99696 2246
rect 109696 1834 109724 41414
rect 111064 34536 111116 34542
rect 111064 34478 111116 34484
rect 109776 4208 109828 4214
rect 109776 4150 109828 4156
rect 109684 1828 109736 1834
rect 109684 1770 109736 1776
rect 98288 1550 98500 1578
rect 98288 800 98316 1550
rect 109788 1426 109816 4150
rect 111076 3942 111104 34478
rect 112444 33176 112496 33182
rect 112444 33118 112496 33124
rect 111156 23520 111208 23526
rect 111156 23462 111208 23468
rect 111064 3936 111116 3942
rect 111064 3878 111116 3884
rect 111168 3534 111196 23462
rect 111248 22160 111300 22166
rect 111248 22102 111300 22108
rect 111156 3528 111208 3534
rect 111156 3470 111208 3476
rect 111260 3466 111288 22102
rect 112456 3874 112484 33118
rect 112536 31816 112588 31822
rect 112536 31758 112588 31764
rect 112444 3868 112496 3874
rect 112444 3810 112496 3816
rect 112548 3806 112576 31758
rect 112628 29028 112680 29034
rect 112628 28970 112680 28976
rect 112536 3800 112588 3806
rect 112536 3742 112588 3748
rect 112640 3738 112668 28970
rect 112720 27668 112772 27674
rect 112720 27610 112772 27616
rect 112628 3732 112680 3738
rect 112628 3674 112680 3680
rect 112732 3670 112760 27610
rect 112812 24880 112864 24886
rect 112812 24822 112864 24828
rect 112720 3664 112772 3670
rect 112720 3606 112772 3612
rect 112824 3602 112852 24822
rect 113836 7721 113864 63514
rect 113928 19009 113956 66234
rect 114020 30433 114048 67594
rect 114112 41857 114140 69022
rect 114204 53145 114232 71742
rect 116306 70272 116362 70281
rect 116306 70207 116362 70216
rect 116320 69086 116348 70207
rect 116308 69080 116360 69086
rect 116308 69022 116360 69028
rect 116122 68368 116178 68377
rect 116122 68303 116178 68312
rect 116136 67658 116164 68303
rect 116124 67652 116176 67658
rect 116124 67594 116176 67600
rect 116582 66464 116638 66473
rect 116582 66399 116638 66408
rect 116596 66298 116624 66399
rect 116584 66292 116636 66298
rect 116584 66234 116636 66240
rect 116688 64874 116716 74015
rect 519740 70553 519768 75919
rect 519832 71913 519860 77415
rect 519924 73273 519952 78911
rect 521014 74488 521070 74497
rect 521014 74423 521070 74432
rect 519910 73264 519966 73273
rect 519910 73199 519966 73208
rect 520922 72992 520978 73001
rect 520922 72927 520978 72936
rect 519818 71904 519874 71913
rect 519818 71839 519874 71848
rect 519726 70544 519782 70553
rect 519726 70479 519782 70488
rect 520936 67833 520964 72927
rect 521028 69193 521056 74423
rect 521198 71496 521254 71505
rect 521198 71431 521254 71440
rect 521106 69864 521162 69873
rect 521106 69799 521162 69808
rect 521014 69184 521070 69193
rect 521014 69119 521070 69128
rect 521014 68368 521070 68377
rect 521014 68303 521070 68312
rect 520922 67824 520978 67833
rect 520922 67759 520978 67768
rect 520462 66872 520518 66881
rect 520462 66807 520518 66816
rect 520370 65376 520426 65385
rect 520370 65311 520426 65320
rect 116596 64846 116716 64874
rect 116596 64598 116624 64846
rect 114468 64592 114520 64598
rect 114466 64560 114468 64569
rect 116584 64592 116636 64598
rect 114520 64560 114522 64569
rect 114466 64495 114522 64504
rect 116214 64560 116270 64569
rect 116584 64534 116636 64540
rect 116214 64495 116270 64504
rect 116228 63578 116256 64495
rect 116216 63572 116268 63578
rect 116216 63514 116268 63520
rect 116582 62656 116638 62665
rect 116582 62591 116638 62600
rect 114190 53136 114246 53145
rect 114190 53071 114246 53080
rect 116490 47152 116546 47161
rect 116490 47087 116546 47096
rect 116214 45248 116270 45257
rect 116214 45183 116270 45192
rect 114098 41848 114154 41857
rect 114098 41783 114154 41792
rect 116124 41472 116176 41478
rect 116122 41440 116124 41449
rect 116176 41440 116178 41449
rect 116122 41375 116178 41384
rect 114100 38684 114152 38690
rect 114100 38626 114152 38632
rect 114006 30424 114062 30433
rect 114006 30359 114062 30368
rect 113914 19000 113970 19009
rect 113914 18935 113970 18944
rect 113822 7712 113878 7721
rect 113822 7647 113878 7656
rect 112812 3596 112864 3602
rect 112812 3538 112864 3544
rect 111248 3460 111300 3466
rect 111248 3402 111300 3408
rect 114112 3330 114140 38626
rect 116228 38554 116256 45183
rect 116306 43344 116362 43353
rect 116306 43279 116362 43288
rect 116216 38548 116268 38554
rect 116216 38490 116268 38496
rect 116214 37632 116270 37641
rect 116214 37567 116270 37576
rect 116228 37330 116256 37567
rect 114192 37324 114244 37330
rect 114192 37266 114244 37272
rect 116216 37324 116268 37330
rect 116216 37266 116268 37272
rect 114204 3398 114232 37266
rect 116122 35728 116178 35737
rect 116122 35663 116178 35672
rect 116136 34542 116164 35663
rect 116124 34536 116176 34542
rect 116124 34478 116176 34484
rect 116122 33824 116178 33833
rect 116122 33759 116178 33768
rect 116136 33182 116164 33759
rect 116124 33176 116176 33182
rect 116124 33118 116176 33124
rect 116124 31816 116176 31822
rect 116122 31784 116124 31793
rect 116176 31784 116178 31793
rect 116122 31719 116178 31728
rect 116122 29880 116178 29889
rect 116122 29815 116178 29824
rect 116136 29034 116164 29815
rect 116124 29028 116176 29034
rect 116124 28970 116176 28976
rect 116122 27976 116178 27985
rect 116122 27911 116178 27920
rect 116136 27674 116164 27911
rect 116124 27668 116176 27674
rect 116124 27610 116176 27616
rect 116122 26072 116178 26081
rect 116122 26007 116178 26016
rect 116136 24886 116164 26007
rect 116124 24880 116176 24886
rect 116124 24822 116176 24828
rect 116122 24168 116178 24177
rect 116122 24103 116178 24112
rect 116136 23526 116164 24103
rect 116124 23520 116176 23526
rect 116124 23462 116176 23468
rect 116030 22264 116086 22273
rect 116030 22199 116086 22208
rect 116044 22166 116072 22199
rect 116032 22160 116084 22166
rect 116032 22102 116084 22108
rect 116214 20360 116270 20369
rect 116214 20295 116270 20304
rect 116122 18456 116178 18465
rect 116122 18391 116178 18400
rect 116032 16516 116084 16522
rect 116032 16458 116084 16464
rect 115938 14512 115994 14521
rect 115938 14447 115994 14456
rect 115952 5234 115980 14447
rect 115940 5228 115992 5234
rect 115940 5170 115992 5176
rect 115940 5092 115992 5098
rect 115940 5034 115992 5040
rect 114192 3392 114244 3398
rect 114192 3334 114244 3340
rect 114100 3324 114152 3330
rect 114100 3266 114152 3272
rect 112444 3256 112496 3262
rect 112444 3198 112496 3204
rect 112456 2990 112484 3198
rect 112444 2984 112496 2990
rect 112444 2926 112496 2932
rect 115952 1630 115980 5034
rect 116044 1698 116072 16458
rect 116136 5098 116164 18391
rect 116228 16522 116256 20295
rect 116216 16516 116268 16522
rect 116216 16458 116268 16464
rect 116214 16416 116270 16425
rect 116214 16351 116270 16360
rect 116228 11898 116256 16351
rect 116216 11892 116268 11898
rect 116216 11834 116268 11840
rect 116320 11778 116348 43279
rect 116398 39536 116454 39545
rect 116398 39471 116454 39480
rect 116412 38690 116440 39471
rect 116400 38684 116452 38690
rect 116400 38626 116452 38632
rect 116400 38548 116452 38554
rect 116400 38490 116452 38496
rect 116228 11750 116348 11778
rect 116124 5092 116176 5098
rect 116124 5034 116176 5040
rect 116122 4992 116178 5001
rect 116122 4927 116178 4936
rect 116136 4214 116164 4927
rect 116124 4208 116176 4214
rect 116124 4150 116176 4156
rect 116122 3088 116178 3097
rect 116122 3023 116178 3032
rect 116136 2922 116164 3023
rect 116124 2916 116176 2922
rect 116124 2858 116176 2864
rect 116228 1766 116256 11750
rect 116308 11688 116360 11694
rect 116308 11630 116360 11636
rect 116320 5370 116348 11630
rect 116308 5364 116360 5370
rect 116308 5306 116360 5312
rect 116308 5228 116360 5234
rect 116308 5170 116360 5176
rect 116216 1760 116268 1766
rect 116216 1702 116268 1708
rect 116032 1692 116084 1698
rect 116032 1634 116084 1640
rect 115940 1624 115992 1630
rect 115940 1566 115992 1572
rect 116320 1494 116348 5170
rect 116412 1902 116440 38490
rect 116504 1970 116532 47087
rect 116596 2514 116624 62591
rect 520384 61033 520412 65311
rect 520476 62393 520504 66807
rect 520738 63880 520794 63889
rect 520738 63815 520794 63824
rect 520462 62384 520518 62393
rect 520462 62319 520518 62328
rect 520370 61024 520426 61033
rect 520370 60959 520426 60968
rect 116674 60616 116730 60625
rect 116674 60551 116730 60560
rect 116584 2508 116636 2514
rect 116584 2450 116636 2456
rect 116688 2446 116716 60551
rect 520752 59673 520780 63815
rect 521028 63753 521056 68303
rect 521120 65113 521148 69799
rect 521212 66473 521240 71431
rect 521198 66464 521254 66473
rect 521198 66399 521254 66408
rect 521106 65104 521162 65113
rect 521106 65039 521162 65048
rect 521014 63744 521070 63753
rect 521014 63679 521070 63688
rect 521014 62384 521070 62393
rect 521014 62319 521070 62328
rect 520738 59664 520794 59673
rect 520738 59599 520794 59608
rect 520738 59392 520794 59401
rect 520738 59327 520794 59336
rect 116766 58712 116822 58721
rect 116766 58647 116822 58656
rect 116676 2440 116728 2446
rect 116676 2382 116728 2388
rect 116780 2378 116808 58647
rect 519910 57896 519966 57905
rect 519910 57831 519966 57840
rect 116858 56808 116914 56817
rect 116858 56743 116914 56752
rect 116768 2372 116820 2378
rect 116768 2314 116820 2320
rect 116872 2310 116900 56743
rect 519818 56400 519874 56409
rect 519818 56335 519874 56344
rect 116950 54904 117006 54913
rect 116950 54839 117006 54848
rect 519082 54904 519138 54913
rect 519082 54839 519138 54848
rect 116964 11506 116992 54839
rect 117042 53000 117098 53009
rect 117042 52935 117098 52944
rect 117056 11642 117084 52935
rect 519096 51513 519124 54839
rect 519832 52873 519860 56335
rect 519924 54233 519952 57831
rect 520752 55593 520780 59327
rect 521028 58313 521056 62319
rect 521106 60888 521162 60897
rect 521106 60823 521162 60832
rect 521014 58304 521070 58313
rect 521014 58239 521070 58248
rect 521120 56953 521148 60823
rect 521106 56944 521162 56953
rect 521106 56879 521162 56888
rect 520738 55584 520794 55593
rect 520738 55519 520794 55528
rect 519910 54224 519966 54233
rect 519910 54159 519966 54168
rect 520186 53408 520242 53417
rect 520186 53343 520242 53352
rect 519818 52864 519874 52873
rect 519818 52799 519874 52808
rect 520094 51912 520150 51921
rect 520094 51847 520150 51856
rect 519082 51504 519138 51513
rect 519082 51439 519138 51448
rect 117134 51096 117190 51105
rect 117134 51031 117190 51040
rect 117148 11778 117176 51031
rect 519082 50416 519138 50425
rect 519082 50351 519138 50360
rect 117226 49192 117282 49201
rect 117226 49127 117282 49136
rect 117240 11914 117268 49127
rect 519096 47433 519124 50351
rect 520108 48793 520136 51847
rect 520200 50153 520228 53343
rect 520186 50144 520242 50153
rect 520186 50079 520242 50088
rect 520186 48920 520242 48929
rect 520186 48855 520242 48864
rect 520094 48784 520150 48793
rect 520094 48719 520150 48728
rect 519082 47424 519138 47433
rect 519082 47359 519138 47368
rect 519450 47288 519506 47297
rect 519450 47223 519506 47232
rect 519464 44713 519492 47223
rect 520200 46073 520228 48855
rect 520186 46064 520242 46073
rect 520186 45999 520242 46008
rect 519726 45792 519782 45801
rect 519726 45727 519782 45736
rect 519450 44704 519506 44713
rect 519450 44639 519506 44648
rect 519740 43353 519768 45727
rect 520186 44296 520242 44305
rect 520186 44231 520242 44240
rect 519726 43344 519782 43353
rect 519726 43279 519782 43288
rect 520200 41993 520228 44231
rect 520738 42800 520794 42809
rect 520738 42735 520794 42744
rect 520186 41984 520242 41993
rect 520186 41919 520242 41928
rect 520752 41313 520780 42735
rect 520738 41304 520794 41313
rect 520738 41239 520794 41248
rect 520922 41304 520978 41313
rect 520922 41239 520978 41248
rect 520936 39953 520964 41239
rect 520922 39944 520978 39953
rect 520922 39879 520978 39888
rect 520922 39808 520978 39817
rect 520922 39743 520978 39752
rect 520936 37913 520964 39743
rect 521106 38312 521162 38321
rect 521106 38247 521162 38256
rect 520922 37904 520978 37913
rect 520922 37839 520978 37848
rect 521120 37233 521148 38247
rect 521106 37224 521162 37233
rect 521106 37159 521162 37168
rect 521566 36816 521622 36825
rect 521566 36751 521622 36760
rect 521580 36009 521608 36751
rect 521566 36000 521622 36009
rect 521566 35935 521622 35944
rect 520922 35320 520978 35329
rect 520922 35255 520978 35264
rect 520936 34513 520964 35255
rect 520922 34504 520978 34513
rect 520922 34439 520978 34448
rect 521106 33824 521162 33833
rect 521106 33759 521162 33768
rect 521120 33153 521148 33759
rect 521106 33144 521162 33153
rect 521106 33079 521162 33088
rect 521106 32328 521162 32337
rect 521106 32263 521162 32272
rect 521120 31657 521148 32263
rect 521106 31648 521162 31657
rect 521106 31583 521162 31592
rect 520922 29336 520978 29345
rect 520922 29271 520978 29280
rect 520936 28393 520964 29271
rect 520922 28384 520978 28393
rect 520922 28319 520978 28328
rect 521106 24848 521162 24857
rect 521106 24783 521162 24792
rect 521120 23633 521148 24783
rect 521106 23624 521162 23633
rect 521106 23559 521162 23568
rect 520370 23216 520426 23225
rect 520370 23151 520426 23160
rect 520384 22273 520412 23151
rect 520370 22264 520426 22273
rect 520370 22199 520426 22208
rect 520922 21720 520978 21729
rect 520922 21655 520978 21664
rect 520936 20913 520964 21655
rect 520922 20904 520978 20913
rect 520922 20839 520978 20848
rect 521106 20224 521162 20233
rect 521106 20159 521162 20168
rect 521120 19553 521148 20159
rect 521106 19544 521162 19553
rect 521106 19479 521162 19488
rect 117240 11886 117360 11914
rect 117148 11750 117268 11778
rect 117056 11614 117176 11642
rect 116964 11478 117084 11506
rect 116952 11416 117004 11422
rect 116952 11358 117004 11364
rect 116964 5506 116992 11358
rect 116952 5500 117004 5506
rect 116952 5442 117004 5448
rect 116952 5364 117004 5370
rect 116952 5306 117004 5312
rect 116860 2304 116912 2310
rect 116860 2246 116912 2252
rect 116492 1964 116544 1970
rect 116492 1906 116544 1912
rect 116400 1896 116452 1902
rect 116400 1838 116452 1844
rect 116964 1562 116992 5306
rect 117056 2242 117084 11478
rect 117148 5658 117176 11614
rect 117240 5794 117268 11750
rect 117332 11422 117360 11886
rect 117320 11416 117372 11422
rect 117320 11358 117372 11364
rect 117240 5766 117360 5794
rect 117148 5630 117268 5658
rect 117136 5500 117188 5506
rect 117136 5442 117188 5448
rect 117044 2236 117096 2242
rect 117044 2178 117096 2184
rect 117148 2038 117176 5442
rect 117240 2174 117268 5630
rect 117228 2168 117280 2174
rect 117228 2110 117280 2116
rect 117332 2106 117360 5766
rect 117964 3052 118016 3058
rect 117964 2994 118016 3000
rect 117688 2984 117740 2990
rect 117688 2926 117740 2932
rect 117320 2100 117372 2106
rect 117320 2042 117372 2048
rect 117136 2032 117188 2038
rect 117136 1974 117188 1980
rect 116952 1556 117004 1562
rect 116952 1498 117004 1504
rect 117700 1494 117728 2926
rect 116308 1488 116360 1494
rect 116308 1430 116360 1436
rect 117688 1488 117740 1494
rect 117688 1430 117740 1436
rect 117976 1426 118004 2994
rect 443656 2514 443992 2530
rect 294788 2508 294840 2514
rect 294788 2450 294840 2456
rect 425796 2508 425848 2514
rect 425796 2450 425848 2456
rect 443644 2508 443992 2514
rect 443696 2502 443992 2508
rect 443644 2450 443696 2456
rect 143644 2094 143980 2122
rect 193600 2094 193936 2122
rect 243648 2094 243984 2122
rect 293604 2094 293940 2122
rect 143644 1494 143672 2094
rect 143632 1488 143684 1494
rect 143632 1430 143684 1436
rect 163778 1456 163834 1465
rect 109776 1420 109828 1426
rect 109776 1362 109828 1368
rect 117964 1420 118016 1426
rect 193600 1426 193628 2094
rect 229282 1592 229338 1601
rect 229282 1527 229338 1536
rect 163778 1391 163834 1400
rect 193588 1420 193640 1426
rect 117964 1362 118016 1368
rect 163792 800 163820 1391
rect 193588 1362 193640 1368
rect 229296 800 229324 1527
rect 243648 1465 243676 2094
rect 293604 1601 293632 2094
rect 293590 1592 293646 1601
rect 293590 1527 293646 1536
rect 243634 1456 243690 1465
rect 294800 1426 294828 2450
rect 343652 2094 343988 2122
rect 393608 2094 393944 2122
rect 343652 1426 343680 2094
rect 393608 1465 393636 2094
rect 360290 1456 360346 1465
rect 243634 1391 243690 1400
rect 294788 1420 294840 1426
rect 294788 1362 294840 1368
rect 343640 1420 343692 1426
rect 360290 1391 360346 1400
rect 393594 1456 393650 1465
rect 393594 1391 393650 1400
rect 343640 1362 343692 1368
rect 294800 800 294828 1362
rect 360304 800 360332 1391
rect 425808 800 425836 2450
rect 493612 2094 493948 2122
rect 493612 1426 493640 2094
rect 491300 1420 491352 1426
rect 491300 1362 491352 1368
rect 493600 1420 493652 1426
rect 493600 1362 493652 1368
rect 491312 800 491340 1362
rect 32770 -400 32826 800
rect 98274 -400 98330 800
rect 163778 -400 163834 800
rect 229282 -400 229338 800
rect 294786 -400 294842 800
rect 360290 -400 360346 800
rect 425794 -400 425850 800
rect 491298 -400 491354 800
<< via2 >>
rect 2962 153720 3018 153776
rect 16302 159296 16358 159352
rect 16578 153856 16634 153912
rect 19890 153992 19946 154048
rect 23018 159432 23074 159488
rect 28078 156712 28134 156768
rect 29826 159568 29882 159624
rect 31482 156576 31538 156632
rect 30378 154128 30434 154184
rect 33966 157936 34022 157992
rect 40682 158208 40738 158264
rect 44086 158072 44142 158128
rect 57518 158344 57574 158400
rect 55862 156848 55918 156904
rect 54298 154264 54354 154320
rect 62578 155488 62634 155544
rect 65982 155352 66038 155408
rect 12438 152496 12494 152552
rect 72698 156984 72754 157040
rect 76010 155760 76066 155816
rect 68466 155216 68522 155272
rect 8850 152360 8906 152416
rect 78586 155624 78642 155680
rect 85302 155896 85358 155952
rect 85578 154400 85634 154456
rect 104622 158480 104678 158536
rect 115570 157120 115626 157176
rect 113822 144200 113878 144256
rect 116122 148996 116124 149016
rect 116124 148996 116176 149016
rect 116176 148996 116178 149016
rect 116122 148960 116178 148996
rect 116122 147056 116178 147112
rect 116214 145152 116270 145208
rect 116030 143248 116086 143304
rect 116398 141344 116454 141400
rect 116122 139440 116178 139496
rect 116490 137536 116546 137592
rect 116122 135496 116178 135552
rect 116030 133592 116086 133648
rect 114190 132776 114246 132832
rect 113914 121352 113970 121408
rect 114006 110064 114062 110120
rect 114098 98640 114154 98696
rect 114466 87236 114522 87272
rect 114466 87216 114468 87236
rect 114468 87216 114520 87236
rect 114520 87216 114522 87236
rect 116122 131688 116178 131744
rect 116122 129784 116178 129840
rect 116122 127880 116178 127936
rect 116030 125976 116086 126032
rect 116122 124108 116124 124128
rect 116124 124108 116176 124128
rect 116176 124108 116178 124128
rect 116122 124072 116178 124108
rect 115938 122168 115994 122224
rect 116122 120128 116178 120184
rect 116122 118224 116178 118280
rect 116122 116320 116178 116376
rect 116122 114452 116124 114472
rect 116124 114452 116176 114472
rect 116176 114452 116178 114472
rect 116122 114416 116178 114452
rect 115938 112512 115994 112568
rect 116122 110608 116178 110664
rect 116122 108704 116178 108760
rect 116490 106800 116546 106856
rect 121734 153720 121790 153776
rect 121918 153720 121974 153776
rect 126242 152360 126298 152416
rect 126610 152360 126666 152416
rect 131026 159296 131082 159352
rect 128818 152496 128874 152552
rect 133602 159432 133658 159488
rect 132038 153856 132094 153912
rect 133602 153040 133658 153096
rect 134614 153992 134670 154048
rect 136546 153040 136602 153096
rect 138018 159568 138074 159624
rect 138386 153584 138442 153640
rect 140410 156712 140466 156768
rect 143170 156576 143226 156632
rect 142342 154128 142398 154184
rect 142618 153992 142674 154048
rect 142526 153856 142582 153912
rect 143262 153992 143318 154048
rect 143354 153876 143410 153912
rect 143354 153856 143356 153876
rect 143356 153856 143408 153876
rect 143408 153856 143410 153876
rect 143538 153584 143594 153640
rect 145102 157936 145158 157992
rect 143630 152360 143686 152416
rect 149610 158208 149666 158264
rect 152554 158072 152610 158128
rect 152186 153856 152242 153912
rect 152646 153856 152702 153912
rect 161662 156848 161718 156904
rect 160926 154264 160982 154320
rect 162858 158344 162914 158400
rect 164882 157836 164884 157856
rect 164884 157836 164936 157856
rect 164936 157836 164938 157856
rect 164882 157800 164938 157836
rect 166722 155488 166778 155544
rect 168378 155352 168434 155408
rect 170494 157836 170496 157856
rect 170496 157836 170548 157856
rect 170548 157836 170550 157856
rect 170494 157800 170550 157836
rect 171230 155216 171286 155272
rect 174450 156984 174506 157040
rect 177026 155760 177082 155816
rect 178958 155624 179014 155680
rect 184018 155896 184074 155952
rect 184662 154400 184718 154456
rect 186318 155080 186374 155136
rect 187238 155080 187294 155136
rect 192390 153720 192446 153776
rect 198738 158480 198794 158536
rect 204718 159296 204774 159352
rect 207202 157120 207258 157176
rect 211526 153720 211582 153776
rect 227442 152360 227498 152416
rect 274546 159432 274602 159488
rect 275190 159296 275246 159352
rect 280986 153720 281042 153776
rect 292578 152360 292634 152416
rect 313646 152360 313702 152416
rect 328550 159432 328606 159488
rect 357438 152360 357494 152416
rect 407578 152360 407634 152416
rect 417882 152260 417884 152280
rect 417884 152260 417936 152280
rect 417936 152260 417938 152280
rect 417882 152224 417938 152260
rect 419906 152260 419908 152280
rect 419908 152260 419960 152280
rect 419960 152260 419962 152280
rect 419906 152224 419962 152260
rect 431222 152496 431278 152552
rect 430578 152360 430634 152416
rect 441894 152940 441896 152960
rect 441896 152940 441948 152960
rect 441948 152940 441950 152960
rect 441894 152904 441950 152940
rect 442538 152940 442540 152960
rect 442540 152940 442592 152960
rect 442592 152940 442594 152960
rect 442538 152904 442594 152940
rect 448610 152496 448666 152552
rect 519358 157120 519414 157176
rect 519726 163104 519782 163160
rect 519542 161608 519598 161664
rect 519634 160112 519690 160168
rect 519542 147872 519598 147928
rect 520002 158616 520058 158672
rect 519818 151136 519874 151192
rect 519726 149232 519782 149288
rect 519726 148144 519782 148200
rect 519634 146512 519690 146568
rect 519634 145016 519690 145072
rect 519358 143792 519414 143848
rect 519542 142160 519598 142216
rect 519450 140528 519506 140584
rect 519266 139032 519322 139088
rect 519358 137536 519414 137592
rect 519266 127472 519322 127528
rect 519910 149640 519966 149696
rect 519818 138352 519874 138408
rect 520094 155624 520150 155680
rect 520002 145152 520058 145208
rect 520186 154128 520242 154184
rect 520094 142432 520150 142488
rect 521106 152632 521162 152688
rect 521014 146648 521070 146704
rect 520922 143656 520978 143712
rect 520186 141072 520242 141128
rect 519910 136992 519966 137048
rect 519910 136040 519966 136096
rect 519726 135632 519782 135688
rect 519726 134544 519782 134600
rect 519634 132912 519690 132968
rect 519542 130192 519598 130248
rect 519450 128832 519506 128888
rect 519542 127064 519598 127120
rect 519358 126112 519414 126168
rect 519266 124072 519322 124128
rect 519174 119584 519230 119640
rect 519450 122576 519506 122632
rect 519358 121080 519414 121136
rect 519266 113872 519322 113928
rect 519634 125568 519690 125624
rect 519542 116592 519598 116648
rect 519818 128560 519874 128616
rect 519726 123392 519782 123448
rect 520002 133048 520058 133104
rect 519910 124752 519966 124808
rect 521106 139712 521162 139768
rect 521014 134272 521070 134328
rect 520922 131688 520978 131744
rect 520094 131552 520150 131608
rect 520002 122032 520058 122088
rect 520186 130056 520242 130112
rect 520094 120672 520150 120728
rect 520186 119312 520242 119368
rect 520002 118088 520058 118144
rect 519818 117952 519874 118008
rect 519910 116456 519966 116512
rect 519634 115232 519690 115288
rect 519818 114960 519874 115016
rect 519726 113464 519782 113520
rect 519450 112512 519506 112568
rect 519634 111968 519690 112024
rect 519358 111152 519414 111208
rect 519542 110472 519598 110528
rect 519174 109792 519230 109848
rect 117134 104760 117190 104816
rect 117042 102856 117098 102912
rect 521106 108976 521162 109032
rect 520002 108432 520058 108488
rect 520830 107480 520886 107536
rect 519910 107072 519966 107128
rect 520278 105984 520334 106040
rect 519818 105712 519874 105768
rect 519726 104352 519782 104408
rect 519634 102992 519690 103048
rect 519542 101632 519598 101688
rect 116950 100952 117006 101008
rect 116858 99048 116914 99104
rect 520738 102992 520794 103048
rect 520278 97552 520334 97608
rect 116766 97144 116822 97200
rect 520278 95512 520334 95568
rect 116674 95240 116730 95296
rect 116582 93336 116638 93392
rect 520186 92384 520242 92440
rect 116122 91296 116178 91352
rect 520094 90888 520150 90944
rect 116122 89392 116178 89448
rect 520002 89392 520058 89448
rect 519818 87896 519874 87952
rect 116030 87488 116086 87544
rect 115202 85584 115258 85640
rect 116214 81776 116270 81832
rect 115938 79872 115994 79928
rect 519634 86400 519690 86456
rect 116582 83680 116638 83736
rect 519266 83408 519322 83464
rect 116490 77968 116546 78024
rect 519542 81912 519598 81968
rect 519450 80416 519506 80472
rect 519266 77152 519322 77208
rect 519726 84904 519782 84960
rect 519634 79872 519690 79928
rect 521014 104488 521070 104544
rect 520830 98912 520886 98968
rect 521474 101496 521530 101552
rect 521106 100272 521162 100328
rect 521382 100000 521438 100056
rect 521290 98504 521346 98560
rect 521106 97008 521162 97064
rect 521014 96192 521070 96248
rect 520738 94832 520794 94888
rect 520922 93880 520978 93936
rect 520278 88032 520334 88088
rect 521474 93472 521530 93528
rect 521382 92112 521438 92168
rect 521290 90752 521346 90808
rect 521106 89528 521162 89584
rect 520922 86672 520978 86728
rect 520186 85312 520242 85368
rect 520094 83952 520150 84008
rect 520002 82592 520058 82648
rect 519818 81232 519874 81288
rect 519910 78920 519966 78976
rect 519726 78512 519782 78568
rect 519818 77424 519874 77480
rect 519542 75928 519598 75984
rect 519726 75928 519782 75984
rect 519450 74568 519506 74624
rect 116674 74024 116730 74080
rect 116582 72120 116638 72176
rect 53654 2644 53710 2680
rect 53654 2624 53656 2644
rect 53656 2624 53708 2644
rect 53708 2624 53710 2644
rect 83002 2644 83058 2680
rect 83002 2624 83004 2644
rect 83004 2624 83056 2644
rect 83056 2624 83058 2644
rect 19338 1808 19394 1864
rect 15934 1672 15990 1728
rect 12622 1536 12678 1592
rect 9310 1400 9366 1456
rect 58714 2488 58770 2544
rect 56138 2388 56140 2408
rect 56140 2388 56192 2408
rect 56192 2388 56194 2408
rect 56138 2352 56194 2388
rect 63498 2352 63554 2408
rect 66350 2352 66406 2408
rect 82082 2488 82138 2544
rect 82358 2524 82360 2544
rect 82360 2524 82412 2544
rect 82412 2524 82414 2544
rect 82358 2488 82414 2524
rect 83094 2488 83150 2544
rect 82726 2352 82782 2408
rect 116306 70216 116362 70272
rect 116122 68312 116178 68368
rect 116582 66408 116638 66464
rect 521014 74432 521070 74488
rect 519910 73208 519966 73264
rect 520922 72936 520978 72992
rect 519818 71848 519874 71904
rect 519726 70488 519782 70544
rect 521198 71440 521254 71496
rect 521106 69808 521162 69864
rect 521014 69128 521070 69184
rect 521014 68312 521070 68368
rect 520922 67768 520978 67824
rect 520462 66816 520518 66872
rect 520370 65320 520426 65376
rect 114466 64540 114468 64560
rect 114468 64540 114520 64560
rect 114520 64540 114522 64560
rect 114466 64504 114522 64540
rect 116214 64504 116270 64560
rect 116582 62600 116638 62656
rect 114190 53080 114246 53136
rect 116490 47096 116546 47152
rect 116214 45192 116270 45248
rect 114098 41792 114154 41848
rect 116122 41420 116124 41440
rect 116124 41420 116176 41440
rect 116176 41420 116178 41440
rect 116122 41384 116178 41420
rect 114006 30368 114062 30424
rect 113914 18944 113970 19000
rect 113822 7656 113878 7712
rect 116306 43288 116362 43344
rect 116214 37576 116270 37632
rect 116122 35672 116178 35728
rect 116122 33768 116178 33824
rect 116122 31764 116124 31784
rect 116124 31764 116176 31784
rect 116176 31764 116178 31784
rect 116122 31728 116178 31764
rect 116122 29824 116178 29880
rect 116122 27920 116178 27976
rect 116122 26016 116178 26072
rect 116122 24112 116178 24168
rect 116030 22208 116086 22264
rect 116214 20304 116270 20360
rect 116122 18400 116178 18456
rect 115938 14456 115994 14512
rect 116214 16360 116270 16416
rect 116398 39480 116454 39536
rect 116122 4936 116178 4992
rect 116122 3032 116178 3088
rect 520738 63824 520794 63880
rect 520462 62328 520518 62384
rect 520370 60968 520426 61024
rect 116674 60560 116730 60616
rect 521198 66408 521254 66464
rect 521106 65048 521162 65104
rect 521014 63688 521070 63744
rect 521014 62328 521070 62384
rect 520738 59608 520794 59664
rect 520738 59336 520794 59392
rect 116766 58656 116822 58712
rect 519910 57840 519966 57896
rect 116858 56752 116914 56808
rect 519818 56344 519874 56400
rect 116950 54848 117006 54904
rect 519082 54848 519138 54904
rect 117042 52944 117098 53000
rect 521106 60832 521162 60888
rect 521014 58248 521070 58304
rect 521106 56888 521162 56944
rect 520738 55528 520794 55584
rect 519910 54168 519966 54224
rect 520186 53352 520242 53408
rect 519818 52808 519874 52864
rect 520094 51856 520150 51912
rect 519082 51448 519138 51504
rect 117134 51040 117190 51096
rect 519082 50360 519138 50416
rect 117226 49136 117282 49192
rect 520186 50088 520242 50144
rect 520186 48864 520242 48920
rect 520094 48728 520150 48784
rect 519082 47368 519138 47424
rect 519450 47232 519506 47288
rect 520186 46008 520242 46064
rect 519726 45736 519782 45792
rect 519450 44648 519506 44704
rect 520186 44240 520242 44296
rect 519726 43288 519782 43344
rect 520738 42744 520794 42800
rect 520186 41928 520242 41984
rect 520738 41248 520794 41304
rect 520922 41248 520978 41304
rect 520922 39888 520978 39944
rect 520922 39752 520978 39808
rect 521106 38256 521162 38312
rect 520922 37848 520978 37904
rect 521106 37168 521162 37224
rect 521566 36760 521622 36816
rect 521566 35944 521622 36000
rect 520922 35264 520978 35320
rect 520922 34448 520978 34504
rect 521106 33768 521162 33824
rect 521106 33088 521162 33144
rect 521106 32272 521162 32328
rect 521106 31592 521162 31648
rect 520922 29280 520978 29336
rect 520922 28328 520978 28384
rect 521106 24792 521162 24848
rect 521106 23568 521162 23624
rect 520370 23160 520426 23216
rect 520370 22208 520426 22264
rect 520922 21664 520978 21720
rect 520922 20848 520978 20904
rect 521106 20168 521162 20224
rect 521106 19488 521162 19544
rect 163778 1400 163834 1456
rect 229282 1536 229338 1592
rect 293590 1536 293646 1592
rect 243634 1400 243690 1456
rect 360290 1400 360346 1456
rect 393594 1400 393650 1456
<< metal3 >>
rect 519721 163162 519787 163165
rect 523200 163162 524400 163192
rect 519721 163160 524400 163162
rect 519721 163104 519726 163160
rect 519782 163104 524400 163160
rect 519721 163102 524400 163104
rect 519721 163099 519787 163102
rect 523200 163072 524400 163102
rect 519537 161666 519603 161669
rect 523200 161666 524400 161696
rect 519537 161664 524400 161666
rect 519537 161608 519542 161664
rect 519598 161608 524400 161664
rect 519537 161606 524400 161608
rect 519537 161603 519603 161606
rect 523200 161576 524400 161606
rect 519629 160170 519695 160173
rect 523200 160170 524400 160200
rect 519629 160168 524400 160170
rect 519629 160112 519634 160168
rect 519690 160112 524400 160168
rect 519629 160110 524400 160112
rect 519629 160107 519695 160110
rect 523200 160080 524400 160110
rect 29821 159626 29887 159629
rect 138013 159626 138079 159629
rect 29821 159624 138079 159626
rect 29821 159568 29826 159624
rect 29882 159568 138018 159624
rect 138074 159568 138079 159624
rect 29821 159566 138079 159568
rect 29821 159563 29887 159566
rect 138013 159563 138079 159566
rect 23013 159490 23079 159493
rect 133597 159490 133663 159493
rect 23013 159488 133663 159490
rect 23013 159432 23018 159488
rect 23074 159432 133602 159488
rect 133658 159432 133663 159488
rect 23013 159430 133663 159432
rect 23013 159427 23079 159430
rect 133597 159427 133663 159430
rect 274541 159490 274607 159493
rect 328545 159490 328611 159493
rect 274541 159488 328611 159490
rect 274541 159432 274546 159488
rect 274602 159432 328550 159488
rect 328606 159432 328611 159488
rect 274541 159430 328611 159432
rect 274541 159427 274607 159430
rect 328545 159427 328611 159430
rect 16297 159354 16363 159357
rect 131021 159354 131087 159357
rect 16297 159352 131087 159354
rect 16297 159296 16302 159352
rect 16358 159296 131026 159352
rect 131082 159296 131087 159352
rect 16297 159294 131087 159296
rect 16297 159291 16363 159294
rect 131021 159291 131087 159294
rect 204713 159354 204779 159357
rect 275185 159354 275251 159357
rect 204713 159352 275251 159354
rect 204713 159296 204718 159352
rect 204774 159296 275190 159352
rect 275246 159296 275251 159352
rect 204713 159294 275251 159296
rect 204713 159291 204779 159294
rect 275185 159291 275251 159294
rect 519997 158674 520063 158677
rect 523200 158674 524400 158704
rect 519997 158672 524400 158674
rect 519997 158616 520002 158672
rect 520058 158616 524400 158672
rect 519997 158614 524400 158616
rect 519997 158611 520063 158614
rect 523200 158584 524400 158614
rect 104617 158538 104683 158541
rect 198733 158538 198799 158541
rect 104617 158536 198799 158538
rect 104617 158480 104622 158536
rect 104678 158480 198738 158536
rect 198794 158480 198799 158536
rect 104617 158478 198799 158480
rect 104617 158475 104683 158478
rect 198733 158475 198799 158478
rect 57513 158402 57579 158405
rect 162853 158402 162919 158405
rect 57513 158400 162919 158402
rect 57513 158344 57518 158400
rect 57574 158344 162858 158400
rect 162914 158344 162919 158400
rect 57513 158342 162919 158344
rect 57513 158339 57579 158342
rect 162853 158339 162919 158342
rect 40677 158266 40743 158269
rect 149605 158266 149671 158269
rect 40677 158264 149671 158266
rect 40677 158208 40682 158264
rect 40738 158208 149610 158264
rect 149666 158208 149671 158264
rect 40677 158206 149671 158208
rect 40677 158203 40743 158206
rect 149605 158203 149671 158206
rect 44081 158130 44147 158133
rect 152549 158130 152615 158133
rect 44081 158128 152615 158130
rect 44081 158072 44086 158128
rect 44142 158072 152554 158128
rect 152610 158072 152615 158128
rect 44081 158070 152615 158072
rect 44081 158067 44147 158070
rect 152549 158067 152615 158070
rect 33961 157994 34027 157997
rect 145097 157994 145163 157997
rect 33961 157992 145163 157994
rect 33961 157936 33966 157992
rect 34022 157936 145102 157992
rect 145158 157936 145163 157992
rect 33961 157934 145163 157936
rect 33961 157931 34027 157934
rect 145097 157931 145163 157934
rect 164877 157858 164943 157861
rect 170489 157858 170555 157861
rect 164877 157856 170555 157858
rect 164877 157800 164882 157856
rect 164938 157800 170494 157856
rect 170550 157800 170555 157856
rect 164877 157798 170555 157800
rect 164877 157795 164943 157798
rect 170489 157795 170555 157798
rect 115565 157178 115631 157181
rect 207197 157178 207263 157181
rect 115565 157176 207263 157178
rect 115565 157120 115570 157176
rect 115626 157120 207202 157176
rect 207258 157120 207263 157176
rect 115565 157118 207263 157120
rect 115565 157115 115631 157118
rect 207197 157115 207263 157118
rect 519353 157178 519419 157181
rect 523200 157178 524400 157208
rect 519353 157176 524400 157178
rect 519353 157120 519358 157176
rect 519414 157120 524400 157176
rect 519353 157118 524400 157120
rect 519353 157115 519419 157118
rect 523200 157088 524400 157118
rect 72693 157042 72759 157045
rect 174445 157042 174511 157045
rect 72693 157040 174511 157042
rect 72693 156984 72698 157040
rect 72754 156984 174450 157040
rect 174506 156984 174511 157040
rect 72693 156982 174511 156984
rect 72693 156979 72759 156982
rect 174445 156979 174511 156982
rect 55857 156906 55923 156909
rect 161657 156906 161723 156909
rect 55857 156904 161723 156906
rect 55857 156848 55862 156904
rect 55918 156848 161662 156904
rect 161718 156848 161723 156904
rect 55857 156846 161723 156848
rect 55857 156843 55923 156846
rect 161657 156843 161723 156846
rect 28073 156770 28139 156773
rect 140405 156770 140471 156773
rect 28073 156768 140471 156770
rect 28073 156712 28078 156768
rect 28134 156712 140410 156768
rect 140466 156712 140471 156768
rect 28073 156710 140471 156712
rect 28073 156707 28139 156710
rect 140405 156707 140471 156710
rect 31477 156634 31543 156637
rect 143165 156634 143231 156637
rect 31477 156632 143231 156634
rect 31477 156576 31482 156632
rect 31538 156576 143170 156632
rect 143226 156576 143231 156632
rect 31477 156574 143231 156576
rect 31477 156571 31543 156574
rect 143165 156571 143231 156574
rect 85297 155954 85363 155957
rect 184013 155954 184079 155957
rect 85297 155952 184079 155954
rect 85297 155896 85302 155952
rect 85358 155896 184018 155952
rect 184074 155896 184079 155952
rect 85297 155894 184079 155896
rect 85297 155891 85363 155894
rect 184013 155891 184079 155894
rect 76005 155818 76071 155821
rect 177021 155818 177087 155821
rect 76005 155816 177087 155818
rect 76005 155760 76010 155816
rect 76066 155760 177026 155816
rect 177082 155760 177087 155816
rect 76005 155758 177087 155760
rect 76005 155755 76071 155758
rect 177021 155755 177087 155758
rect 78581 155682 78647 155685
rect 178953 155682 179019 155685
rect 78581 155680 179019 155682
rect 78581 155624 78586 155680
rect 78642 155624 178958 155680
rect 179014 155624 179019 155680
rect 78581 155622 179019 155624
rect 78581 155619 78647 155622
rect 178953 155619 179019 155622
rect 520089 155682 520155 155685
rect 523200 155682 524400 155712
rect 520089 155680 524400 155682
rect 520089 155624 520094 155680
rect 520150 155624 524400 155680
rect 520089 155622 524400 155624
rect 520089 155619 520155 155622
rect 523200 155592 524400 155622
rect 62573 155546 62639 155549
rect 166717 155546 166783 155549
rect 62573 155544 166783 155546
rect 62573 155488 62578 155544
rect 62634 155488 166722 155544
rect 166778 155488 166783 155544
rect 62573 155486 166783 155488
rect 62573 155483 62639 155486
rect 166717 155483 166783 155486
rect 65977 155410 66043 155413
rect 168373 155410 168439 155413
rect 65977 155408 168439 155410
rect 65977 155352 65982 155408
rect 66038 155352 168378 155408
rect 168434 155352 168439 155408
rect 65977 155350 168439 155352
rect 65977 155347 66043 155350
rect 168373 155347 168439 155350
rect 68461 155274 68527 155277
rect 171225 155274 171291 155277
rect 68461 155272 171291 155274
rect 68461 155216 68466 155272
rect 68522 155216 171230 155272
rect 171286 155216 171291 155272
rect 68461 155214 171291 155216
rect 68461 155211 68527 155214
rect 171225 155211 171291 155214
rect 186313 155138 186379 155141
rect 187233 155138 187299 155141
rect 186313 155136 187299 155138
rect 186313 155080 186318 155136
rect 186374 155080 187238 155136
rect 187294 155080 187299 155136
rect 186313 155078 187299 155080
rect 186313 155075 186379 155078
rect 187233 155075 187299 155078
rect 85573 154458 85639 154461
rect 184657 154458 184723 154461
rect 85573 154456 184723 154458
rect 85573 154400 85578 154456
rect 85634 154400 184662 154456
rect 184718 154400 184723 154456
rect 85573 154398 184723 154400
rect 85573 154395 85639 154398
rect 184657 154395 184723 154398
rect 54293 154322 54359 154325
rect 160921 154322 160987 154325
rect 54293 154320 160987 154322
rect 54293 154264 54298 154320
rect 54354 154264 160926 154320
rect 160982 154264 160987 154320
rect 54293 154262 160987 154264
rect 54293 154259 54359 154262
rect 160921 154259 160987 154262
rect 30373 154186 30439 154189
rect 142337 154186 142403 154189
rect 30373 154184 142403 154186
rect 30373 154128 30378 154184
rect 30434 154128 142342 154184
rect 142398 154128 142403 154184
rect 30373 154126 142403 154128
rect 30373 154123 30439 154126
rect 142337 154123 142403 154126
rect 520181 154186 520247 154189
rect 523200 154186 524400 154216
rect 520181 154184 524400 154186
rect 520181 154128 520186 154184
rect 520242 154128 524400 154184
rect 520181 154126 524400 154128
rect 520181 154123 520247 154126
rect 523200 154096 524400 154126
rect 19885 154050 19951 154053
rect 134609 154050 134675 154053
rect 19885 154048 134675 154050
rect 19885 153992 19890 154048
rect 19946 153992 134614 154048
rect 134670 153992 134675 154048
rect 19885 153990 134675 153992
rect 19885 153987 19951 153990
rect 134609 153987 134675 153990
rect 142613 154050 142679 154053
rect 143257 154050 143323 154053
rect 142613 154048 143323 154050
rect 142613 153992 142618 154048
rect 142674 153992 143262 154048
rect 143318 153992 143323 154048
rect 142613 153990 143323 153992
rect 142613 153987 142679 153990
rect 143257 153987 143323 153990
rect 16573 153914 16639 153917
rect 132033 153914 132099 153917
rect 16573 153912 132099 153914
rect 16573 153856 16578 153912
rect 16634 153856 132038 153912
rect 132094 153856 132099 153912
rect 16573 153854 132099 153856
rect 16573 153851 16639 153854
rect 132033 153851 132099 153854
rect 142521 153914 142587 153917
rect 143349 153914 143415 153917
rect 142521 153912 143415 153914
rect 142521 153856 142526 153912
rect 142582 153856 143354 153912
rect 143410 153856 143415 153912
rect 142521 153854 143415 153856
rect 142521 153851 142587 153854
rect 143349 153851 143415 153854
rect 152181 153914 152247 153917
rect 152641 153914 152707 153917
rect 152181 153912 152707 153914
rect 152181 153856 152186 153912
rect 152242 153856 152646 153912
rect 152702 153856 152707 153912
rect 152181 153854 152707 153856
rect 152181 153851 152247 153854
rect 152641 153851 152707 153854
rect 2957 153778 3023 153781
rect 121729 153778 121795 153781
rect 2957 153776 121795 153778
rect 2957 153720 2962 153776
rect 3018 153720 121734 153776
rect 121790 153720 121795 153776
rect 2957 153718 121795 153720
rect 2957 153715 3023 153718
rect 121729 153715 121795 153718
rect 121913 153778 121979 153781
rect 192385 153778 192451 153781
rect 121913 153776 192451 153778
rect 121913 153720 121918 153776
rect 121974 153720 192390 153776
rect 192446 153720 192451 153776
rect 121913 153718 192451 153720
rect 121913 153715 121979 153718
rect 192385 153715 192451 153718
rect 211521 153778 211587 153781
rect 280981 153778 281047 153781
rect 211521 153776 281047 153778
rect 211521 153720 211526 153776
rect 211582 153720 280986 153776
rect 281042 153720 281047 153776
rect 211521 153718 281047 153720
rect 211521 153715 211587 153718
rect 280981 153715 281047 153718
rect 138381 153642 138447 153645
rect 143533 153642 143599 153645
rect 138381 153640 143599 153642
rect 138381 153584 138386 153640
rect 138442 153584 143538 153640
rect 143594 153584 143599 153640
rect 138381 153582 143599 153584
rect 138381 153579 138447 153582
rect 143533 153579 143599 153582
rect 133597 153098 133663 153101
rect 136541 153098 136607 153101
rect 133597 153096 136607 153098
rect 133597 153040 133602 153096
rect 133658 153040 136546 153096
rect 136602 153040 136607 153096
rect 133597 153038 136607 153040
rect 133597 153035 133663 153038
rect 136541 153035 136607 153038
rect 441889 152962 441955 152965
rect 442533 152962 442599 152965
rect 441889 152960 442599 152962
rect 441889 152904 441894 152960
rect 441950 152904 442538 152960
rect 442594 152904 442599 152960
rect 441889 152902 442599 152904
rect 441889 152899 441955 152902
rect 442533 152899 442599 152902
rect 521101 152690 521167 152693
rect 523200 152690 524400 152720
rect 521101 152688 524400 152690
rect 521101 152632 521106 152688
rect 521162 152632 524400 152688
rect 521101 152630 524400 152632
rect 521101 152627 521167 152630
rect 523200 152600 524400 152630
rect 12433 152554 12499 152557
rect 128813 152554 128879 152557
rect 12433 152552 128879 152554
rect 12433 152496 12438 152552
rect 12494 152496 128818 152552
rect 128874 152496 128879 152552
rect 12433 152494 128879 152496
rect 12433 152491 12499 152494
rect 128813 152491 128879 152494
rect 431217 152554 431283 152557
rect 448605 152554 448671 152557
rect 431217 152552 448671 152554
rect 431217 152496 431222 152552
rect 431278 152496 448610 152552
rect 448666 152496 448671 152552
rect 431217 152494 448671 152496
rect 431217 152491 431283 152494
rect 448605 152491 448671 152494
rect 8845 152418 8911 152421
rect 126237 152418 126303 152421
rect 8845 152416 126303 152418
rect 8845 152360 8850 152416
rect 8906 152360 126242 152416
rect 126298 152360 126303 152416
rect 8845 152358 126303 152360
rect 8845 152355 8911 152358
rect 126237 152355 126303 152358
rect 126605 152418 126671 152421
rect 143625 152418 143691 152421
rect 126605 152416 143691 152418
rect 126605 152360 126610 152416
rect 126666 152360 143630 152416
rect 143686 152360 143691 152416
rect 126605 152358 143691 152360
rect 126605 152355 126671 152358
rect 143625 152355 143691 152358
rect 227437 152418 227503 152421
rect 292573 152418 292639 152421
rect 227437 152416 292639 152418
rect 227437 152360 227442 152416
rect 227498 152360 292578 152416
rect 292634 152360 292639 152416
rect 227437 152358 292639 152360
rect 227437 152355 227503 152358
rect 292573 152355 292639 152358
rect 313641 152418 313707 152421
rect 357433 152418 357499 152421
rect 313641 152416 357499 152418
rect 313641 152360 313646 152416
rect 313702 152360 357438 152416
rect 357494 152360 357499 152416
rect 313641 152358 357499 152360
rect 313641 152355 313707 152358
rect 357433 152355 357499 152358
rect 407573 152418 407639 152421
rect 430573 152418 430639 152421
rect 407573 152416 430639 152418
rect 407573 152360 407578 152416
rect 407634 152360 430578 152416
rect 430634 152360 430639 152416
rect 407573 152358 430639 152360
rect 407573 152355 407639 152358
rect 430573 152355 430639 152358
rect 417877 152282 417943 152285
rect 419901 152282 419967 152285
rect 417877 152280 419967 152282
rect 417877 152224 417882 152280
rect 417938 152224 419906 152280
rect 419962 152224 419967 152280
rect 417877 152222 419967 152224
rect 417877 152219 417943 152222
rect 419901 152219 419967 152222
rect 519813 151194 519879 151197
rect 523200 151194 524400 151224
rect 519813 151192 524400 151194
rect 519813 151136 519818 151192
rect 519874 151136 524400 151192
rect 519813 151134 524400 151136
rect 519813 151131 519879 151134
rect 523200 151104 524400 151134
rect 519905 149698 519971 149701
rect 523200 149698 524400 149728
rect 519905 149696 524400 149698
rect 519905 149640 519910 149696
rect 519966 149640 524400 149696
rect 519905 149638 524400 149640
rect 519905 149635 519971 149638
rect 523200 149608 524400 149638
rect 519721 149290 519787 149293
rect 518788 149288 519787 149290
rect 518788 149232 519726 149288
rect 519782 149232 519787 149288
rect 518788 149230 519787 149232
rect 519721 149227 519787 149230
rect 116117 149018 116183 149021
rect 116117 149016 119140 149018
rect 116117 148960 116122 149016
rect 116178 148960 119140 149016
rect 116117 148958 119140 148960
rect 116117 148955 116183 148958
rect 519721 148202 519787 148205
rect 523200 148202 524400 148232
rect 519721 148200 524400 148202
rect 519721 148144 519726 148200
rect 519782 148144 524400 148200
rect 519721 148142 524400 148144
rect 519721 148139 519787 148142
rect 523200 148112 524400 148142
rect 519537 147930 519603 147933
rect 518788 147928 519603 147930
rect 518788 147872 519542 147928
rect 519598 147872 519603 147928
rect 518788 147870 519603 147872
rect 519537 147867 519603 147870
rect 116117 147114 116183 147117
rect 116117 147112 119140 147114
rect 116117 147056 116122 147112
rect 116178 147056 119140 147112
rect 116117 147054 119140 147056
rect 116117 147051 116183 147054
rect 521009 146706 521075 146709
rect 523200 146706 524400 146736
rect 521009 146704 524400 146706
rect 521009 146648 521014 146704
rect 521070 146648 524400 146704
rect 521009 146646 524400 146648
rect 521009 146643 521075 146646
rect 523200 146616 524400 146646
rect 519629 146570 519695 146573
rect 518788 146568 519695 146570
rect 518788 146512 519634 146568
rect 519690 146512 519695 146568
rect 518788 146510 519695 146512
rect 519629 146507 519695 146510
rect 116209 145210 116275 145213
rect 519997 145210 520063 145213
rect 523200 145210 524400 145240
rect 116209 145208 119140 145210
rect 116209 145152 116214 145208
rect 116270 145152 119140 145208
rect 116209 145150 119140 145152
rect 518788 145208 520063 145210
rect 518788 145152 520002 145208
rect 520058 145152 520063 145208
rect 518788 145150 520063 145152
rect 116209 145147 116275 145150
rect 519997 145147 520063 145150
rect 520230 145150 524400 145210
rect 519629 145074 519695 145077
rect 520230 145074 520290 145150
rect 523200 145120 524400 145150
rect 519629 145072 520290 145074
rect 519629 145016 519634 145072
rect 519690 145016 520290 145072
rect 519629 145014 520290 145016
rect 519629 145011 519695 145014
rect 113817 144258 113883 144261
rect 110860 144256 113883 144258
rect 110860 144200 113822 144256
rect 113878 144200 113883 144256
rect 110860 144198 113883 144200
rect 113817 144195 113883 144198
rect 519353 143850 519419 143853
rect 518788 143848 519419 143850
rect 518788 143792 519358 143848
rect 519414 143792 519419 143848
rect 518788 143790 519419 143792
rect 519353 143787 519419 143790
rect 520917 143714 520983 143717
rect 523200 143714 524400 143744
rect 520917 143712 524400 143714
rect 520917 143656 520922 143712
rect 520978 143656 524400 143712
rect 520917 143654 524400 143656
rect 520917 143651 520983 143654
rect 523200 143624 524400 143654
rect 116025 143306 116091 143309
rect 116025 143304 119140 143306
rect 116025 143248 116030 143304
rect 116086 143248 119140 143304
rect 116025 143246 119140 143248
rect 116025 143243 116091 143246
rect 520089 142490 520155 142493
rect 518788 142488 520155 142490
rect 518788 142432 520094 142488
rect 520150 142432 520155 142488
rect 518788 142430 520155 142432
rect 520089 142427 520155 142430
rect 519537 142218 519603 142221
rect 523200 142218 524400 142248
rect 519537 142216 524400 142218
rect 519537 142160 519542 142216
rect 519598 142160 524400 142216
rect 519537 142158 524400 142160
rect 519537 142155 519603 142158
rect 523200 142128 524400 142158
rect 116393 141402 116459 141405
rect 116393 141400 119140 141402
rect 116393 141344 116398 141400
rect 116454 141344 119140 141400
rect 116393 141342 119140 141344
rect 116393 141339 116459 141342
rect 520181 141130 520247 141133
rect 518788 141128 520247 141130
rect 518788 141072 520186 141128
rect 520242 141072 520247 141128
rect 518788 141070 520247 141072
rect 520181 141067 520247 141070
rect 519445 140586 519511 140589
rect 523200 140586 524400 140616
rect 519445 140584 524400 140586
rect 519445 140528 519450 140584
rect 519506 140528 524400 140584
rect 519445 140526 524400 140528
rect 519445 140523 519511 140526
rect 523200 140496 524400 140526
rect 521101 139770 521167 139773
rect 518788 139768 521167 139770
rect 518788 139712 521106 139768
rect 521162 139712 521167 139768
rect 518788 139710 521167 139712
rect 521101 139707 521167 139710
rect 116117 139498 116183 139501
rect 116117 139496 119140 139498
rect 116117 139440 116122 139496
rect 116178 139440 119140 139496
rect 116117 139438 119140 139440
rect 116117 139435 116183 139438
rect 519261 139090 519327 139093
rect 523200 139090 524400 139120
rect 519261 139088 524400 139090
rect 519261 139032 519266 139088
rect 519322 139032 524400 139088
rect 519261 139030 524400 139032
rect 519261 139027 519327 139030
rect 523200 139000 524400 139030
rect 519813 138410 519879 138413
rect 518788 138408 519879 138410
rect 518788 138352 519818 138408
rect 519874 138352 519879 138408
rect 518788 138350 519879 138352
rect 519813 138347 519879 138350
rect 116485 137594 116551 137597
rect 519353 137594 519419 137597
rect 523200 137594 524400 137624
rect 116485 137592 119140 137594
rect 116485 137536 116490 137592
rect 116546 137536 119140 137592
rect 116485 137534 119140 137536
rect 519353 137592 524400 137594
rect 519353 137536 519358 137592
rect 519414 137536 524400 137592
rect 519353 137534 524400 137536
rect 116485 137531 116551 137534
rect 519353 137531 519419 137534
rect 523200 137504 524400 137534
rect 519905 137050 519971 137053
rect 518788 137048 519971 137050
rect 518788 136992 519910 137048
rect 519966 136992 519971 137048
rect 518788 136990 519971 136992
rect 519905 136987 519971 136990
rect 519905 136098 519971 136101
rect 523200 136098 524400 136128
rect 519905 136096 524400 136098
rect 519905 136040 519910 136096
rect 519966 136040 524400 136096
rect 519905 136038 524400 136040
rect 519905 136035 519971 136038
rect 523200 136008 524400 136038
rect 519721 135690 519787 135693
rect 518788 135688 519787 135690
rect 518788 135632 519726 135688
rect 519782 135632 519787 135688
rect 518788 135630 519787 135632
rect 519721 135627 519787 135630
rect 116117 135554 116183 135557
rect 116117 135552 119140 135554
rect 116117 135496 116122 135552
rect 116178 135496 119140 135552
rect 116117 135494 119140 135496
rect 116117 135491 116183 135494
rect 519721 134602 519787 134605
rect 523200 134602 524400 134632
rect 519721 134600 524400 134602
rect 519721 134544 519726 134600
rect 519782 134544 524400 134600
rect 519721 134542 524400 134544
rect 519721 134539 519787 134542
rect 523200 134512 524400 134542
rect 521009 134330 521075 134333
rect 518788 134328 521075 134330
rect 518788 134272 521014 134328
rect 521070 134272 521075 134328
rect 518788 134270 521075 134272
rect 521009 134267 521075 134270
rect 116025 133650 116091 133653
rect 116025 133648 119140 133650
rect 116025 133592 116030 133648
rect 116086 133592 119140 133648
rect 116025 133590 119140 133592
rect 116025 133587 116091 133590
rect 519997 133106 520063 133109
rect 523200 133106 524400 133136
rect 519997 133104 524400 133106
rect 519997 133048 520002 133104
rect 520058 133048 524400 133104
rect 519997 133046 524400 133048
rect 519997 133043 520063 133046
rect 523200 133016 524400 133046
rect 519629 132970 519695 132973
rect 518788 132968 519695 132970
rect 518788 132912 519634 132968
rect 519690 132912 519695 132968
rect 518788 132910 519695 132912
rect 519629 132907 519695 132910
rect 114185 132834 114251 132837
rect 110860 132832 114251 132834
rect 110860 132776 114190 132832
rect 114246 132776 114251 132832
rect 110860 132774 114251 132776
rect 114185 132771 114251 132774
rect 116117 131746 116183 131749
rect 520917 131746 520983 131749
rect 116117 131744 119140 131746
rect 116117 131688 116122 131744
rect 116178 131688 119140 131744
rect 116117 131686 119140 131688
rect 518758 131744 520983 131746
rect 518758 131688 520922 131744
rect 520978 131688 520983 131744
rect 518758 131686 520983 131688
rect 116117 131683 116183 131686
rect 518758 131580 518818 131686
rect 520917 131683 520983 131686
rect 520089 131610 520155 131613
rect 523200 131610 524400 131640
rect 520089 131608 524400 131610
rect 520089 131552 520094 131608
rect 520150 131552 524400 131608
rect 520089 131550 524400 131552
rect 520089 131547 520155 131550
rect 523200 131520 524400 131550
rect 519537 130250 519603 130253
rect 518788 130248 519603 130250
rect 518788 130192 519542 130248
rect 519598 130192 519603 130248
rect 518788 130190 519603 130192
rect 519537 130187 519603 130190
rect 520181 130114 520247 130117
rect 523200 130114 524400 130144
rect 520181 130112 524400 130114
rect 520181 130056 520186 130112
rect 520242 130056 524400 130112
rect 520181 130054 524400 130056
rect 520181 130051 520247 130054
rect 523200 130024 524400 130054
rect 116117 129842 116183 129845
rect 116117 129840 119140 129842
rect 116117 129784 116122 129840
rect 116178 129784 119140 129840
rect 116117 129782 119140 129784
rect 116117 129779 116183 129782
rect 519445 128890 519511 128893
rect 518788 128888 519511 128890
rect 518788 128832 519450 128888
rect 519506 128832 519511 128888
rect 518788 128830 519511 128832
rect 519445 128827 519511 128830
rect 519813 128618 519879 128621
rect 523200 128618 524400 128648
rect 519813 128616 524400 128618
rect 519813 128560 519818 128616
rect 519874 128560 524400 128616
rect 519813 128558 524400 128560
rect 519813 128555 519879 128558
rect 523200 128528 524400 128558
rect 116117 127938 116183 127941
rect 116117 127936 119140 127938
rect 116117 127880 116122 127936
rect 116178 127880 119140 127936
rect 116117 127878 119140 127880
rect 116117 127875 116183 127878
rect 519261 127530 519327 127533
rect 518788 127528 519327 127530
rect 518788 127472 519266 127528
rect 519322 127472 519327 127528
rect 518788 127470 519327 127472
rect 519261 127467 519327 127470
rect 519537 127122 519603 127125
rect 523200 127122 524400 127152
rect 519537 127120 524400 127122
rect 519537 127064 519542 127120
rect 519598 127064 524400 127120
rect 519537 127062 524400 127064
rect 519537 127059 519603 127062
rect 523200 127032 524400 127062
rect 519353 126170 519419 126173
rect 518788 126168 519419 126170
rect 518788 126112 519358 126168
rect 519414 126112 519419 126168
rect 518788 126110 519419 126112
rect 519353 126107 519419 126110
rect 116025 126034 116091 126037
rect 116025 126032 119140 126034
rect 116025 125976 116030 126032
rect 116086 125976 119140 126032
rect 116025 125974 119140 125976
rect 116025 125971 116091 125974
rect 519629 125626 519695 125629
rect 523200 125626 524400 125656
rect 519629 125624 524400 125626
rect 519629 125568 519634 125624
rect 519690 125568 524400 125624
rect 519629 125566 524400 125568
rect 519629 125563 519695 125566
rect 523200 125536 524400 125566
rect 519905 124810 519971 124813
rect 518788 124808 519971 124810
rect 518788 124752 519910 124808
rect 519966 124752 519971 124808
rect 518788 124750 519971 124752
rect 519905 124747 519971 124750
rect 116117 124130 116183 124133
rect 519261 124130 519327 124133
rect 523200 124130 524400 124160
rect 116117 124128 119140 124130
rect 116117 124072 116122 124128
rect 116178 124072 119140 124128
rect 116117 124070 119140 124072
rect 519261 124128 524400 124130
rect 519261 124072 519266 124128
rect 519322 124072 524400 124128
rect 519261 124070 524400 124072
rect 116117 124067 116183 124070
rect 519261 124067 519327 124070
rect 523200 124040 524400 124070
rect 519721 123450 519787 123453
rect 518788 123448 519787 123450
rect 518788 123392 519726 123448
rect 519782 123392 519787 123448
rect 518788 123390 519787 123392
rect 519721 123387 519787 123390
rect 519445 122634 519511 122637
rect 523200 122634 524400 122664
rect 519445 122632 524400 122634
rect 519445 122576 519450 122632
rect 519506 122576 524400 122632
rect 519445 122574 524400 122576
rect 519445 122571 519511 122574
rect 523200 122544 524400 122574
rect 115933 122226 115999 122229
rect 115933 122224 119140 122226
rect 115933 122168 115938 122224
rect 115994 122168 119140 122224
rect 115933 122166 119140 122168
rect 115933 122163 115999 122166
rect 519997 122090 520063 122093
rect 518788 122088 520063 122090
rect 518788 122032 520002 122088
rect 520058 122032 520063 122088
rect 518788 122030 520063 122032
rect 519997 122027 520063 122030
rect 113909 121410 113975 121413
rect 110860 121408 113975 121410
rect 110860 121352 113914 121408
rect 113970 121352 113975 121408
rect 110860 121350 113975 121352
rect 113909 121347 113975 121350
rect 519353 121138 519419 121141
rect 523200 121138 524400 121168
rect 519353 121136 524400 121138
rect 519353 121080 519358 121136
rect 519414 121080 524400 121136
rect 519353 121078 524400 121080
rect 519353 121075 519419 121078
rect 523200 121048 524400 121078
rect 520089 120730 520155 120733
rect 518788 120728 520155 120730
rect 518788 120672 520094 120728
rect 520150 120672 520155 120728
rect 518788 120670 520155 120672
rect 520089 120667 520155 120670
rect 116117 120186 116183 120189
rect 116117 120184 119140 120186
rect 116117 120128 116122 120184
rect 116178 120128 119140 120184
rect 116117 120126 119140 120128
rect 116117 120123 116183 120126
rect 519169 119642 519235 119645
rect 523200 119642 524400 119672
rect 519169 119640 524400 119642
rect 519169 119584 519174 119640
rect 519230 119584 524400 119640
rect 519169 119582 524400 119584
rect 519169 119579 519235 119582
rect 523200 119552 524400 119582
rect 520181 119370 520247 119373
rect 518788 119368 520247 119370
rect 518788 119312 520186 119368
rect 520242 119312 520247 119368
rect 518788 119310 520247 119312
rect 520181 119307 520247 119310
rect 116117 118282 116183 118285
rect 116117 118280 119140 118282
rect 116117 118224 116122 118280
rect 116178 118224 119140 118280
rect 116117 118222 119140 118224
rect 116117 118219 116183 118222
rect 519997 118146 520063 118149
rect 523200 118146 524400 118176
rect 519997 118144 524400 118146
rect 519997 118088 520002 118144
rect 520058 118088 524400 118144
rect 519997 118086 524400 118088
rect 519997 118083 520063 118086
rect 523200 118056 524400 118086
rect 519813 118010 519879 118013
rect 518788 118008 519879 118010
rect 518788 117952 519818 118008
rect 519874 117952 519879 118008
rect 518788 117950 519879 117952
rect 519813 117947 519879 117950
rect 519537 116650 519603 116653
rect 518788 116648 519603 116650
rect 518788 116592 519542 116648
rect 519598 116592 519603 116648
rect 518788 116590 519603 116592
rect 519537 116587 519603 116590
rect 519905 116514 519971 116517
rect 523200 116514 524400 116544
rect 519905 116512 524400 116514
rect 519905 116456 519910 116512
rect 519966 116456 524400 116512
rect 519905 116454 524400 116456
rect 519905 116451 519971 116454
rect 523200 116424 524400 116454
rect 116117 116378 116183 116381
rect 116117 116376 119140 116378
rect 116117 116320 116122 116376
rect 116178 116320 119140 116376
rect 116117 116318 119140 116320
rect 116117 116315 116183 116318
rect 519629 115290 519695 115293
rect 518788 115288 519695 115290
rect 518788 115232 519634 115288
rect 519690 115232 519695 115288
rect 518788 115230 519695 115232
rect 519629 115227 519695 115230
rect 519813 115018 519879 115021
rect 523200 115018 524400 115048
rect 519813 115016 524400 115018
rect 519813 114960 519818 115016
rect 519874 114960 524400 115016
rect 519813 114958 524400 114960
rect 519813 114955 519879 114958
rect 523200 114928 524400 114958
rect 116117 114474 116183 114477
rect 116117 114472 119140 114474
rect 116117 114416 116122 114472
rect 116178 114416 119140 114472
rect 116117 114414 119140 114416
rect 116117 114411 116183 114414
rect 519261 113930 519327 113933
rect 518788 113928 519327 113930
rect 518788 113872 519266 113928
rect 519322 113872 519327 113928
rect 518788 113870 519327 113872
rect 519261 113867 519327 113870
rect 519721 113522 519787 113525
rect 523200 113522 524400 113552
rect 519721 113520 524400 113522
rect 519721 113464 519726 113520
rect 519782 113464 524400 113520
rect 519721 113462 524400 113464
rect 519721 113459 519787 113462
rect 523200 113432 524400 113462
rect 115933 112570 115999 112573
rect 519445 112570 519511 112573
rect 115933 112568 119140 112570
rect 115933 112512 115938 112568
rect 115994 112512 119140 112568
rect 115933 112510 119140 112512
rect 518788 112568 519511 112570
rect 518788 112512 519450 112568
rect 519506 112512 519511 112568
rect 518788 112510 519511 112512
rect 115933 112507 115999 112510
rect 519445 112507 519511 112510
rect 519629 112026 519695 112029
rect 523200 112026 524400 112056
rect 519629 112024 524400 112026
rect 519629 111968 519634 112024
rect 519690 111968 524400 112024
rect 519629 111966 524400 111968
rect 519629 111963 519695 111966
rect 523200 111936 524400 111966
rect 519353 111210 519419 111213
rect 518788 111208 519419 111210
rect 518788 111152 519358 111208
rect 519414 111152 519419 111208
rect 518788 111150 519419 111152
rect 519353 111147 519419 111150
rect 116117 110666 116183 110669
rect 116117 110664 119140 110666
rect 116117 110608 116122 110664
rect 116178 110608 119140 110664
rect 116117 110606 119140 110608
rect 116117 110603 116183 110606
rect 519537 110530 519603 110533
rect 523200 110530 524400 110560
rect 519537 110528 524400 110530
rect 519537 110472 519542 110528
rect 519598 110472 524400 110528
rect 519537 110470 524400 110472
rect 519537 110467 519603 110470
rect 523200 110440 524400 110470
rect 114001 110122 114067 110125
rect 110860 110120 114067 110122
rect 110860 110064 114006 110120
rect 114062 110064 114067 110120
rect 110860 110062 114067 110064
rect 114001 110059 114067 110062
rect 519169 109850 519235 109853
rect 518788 109848 519235 109850
rect 518788 109792 519174 109848
rect 519230 109792 519235 109848
rect 518788 109790 519235 109792
rect 519169 109787 519235 109790
rect 521101 109034 521167 109037
rect 523200 109034 524400 109064
rect 521101 109032 524400 109034
rect 521101 108976 521106 109032
rect 521162 108976 524400 109032
rect 521101 108974 524400 108976
rect 521101 108971 521167 108974
rect 523200 108944 524400 108974
rect 116117 108762 116183 108765
rect 116117 108760 119140 108762
rect 116117 108704 116122 108760
rect 116178 108704 119140 108760
rect 116117 108702 119140 108704
rect 116117 108699 116183 108702
rect 519997 108490 520063 108493
rect 518788 108488 520063 108490
rect 518788 108432 520002 108488
rect 520058 108432 520063 108488
rect 518788 108430 520063 108432
rect 519997 108427 520063 108430
rect 520825 107538 520891 107541
rect 523200 107538 524400 107568
rect 520825 107536 524400 107538
rect 520825 107480 520830 107536
rect 520886 107480 524400 107536
rect 520825 107478 524400 107480
rect 520825 107475 520891 107478
rect 523200 107448 524400 107478
rect 519905 107130 519971 107133
rect 518788 107128 519971 107130
rect 518788 107072 519910 107128
rect 519966 107072 519971 107128
rect 518788 107070 519971 107072
rect 519905 107067 519971 107070
rect 116485 106858 116551 106861
rect 116485 106856 119140 106858
rect 116485 106800 116490 106856
rect 116546 106800 119140 106856
rect 116485 106798 119140 106800
rect 116485 106795 116551 106798
rect 520273 106042 520339 106045
rect 523200 106042 524400 106072
rect 520273 106040 524400 106042
rect 520273 105984 520278 106040
rect 520334 105984 524400 106040
rect 520273 105982 524400 105984
rect 520273 105979 520339 105982
rect 523200 105952 524400 105982
rect 519813 105770 519879 105773
rect 518788 105768 519879 105770
rect 518788 105712 519818 105768
rect 519874 105712 519879 105768
rect 518788 105710 519879 105712
rect 519813 105707 519879 105710
rect 117129 104818 117195 104821
rect 117129 104816 119140 104818
rect 117129 104760 117134 104816
rect 117190 104760 119140 104816
rect 117129 104758 119140 104760
rect 117129 104755 117195 104758
rect 521009 104546 521075 104549
rect 523200 104546 524400 104576
rect 521009 104544 524400 104546
rect 521009 104488 521014 104544
rect 521070 104488 524400 104544
rect 521009 104486 524400 104488
rect 521009 104483 521075 104486
rect 523200 104456 524400 104486
rect 519721 104410 519787 104413
rect 518788 104408 519787 104410
rect 518788 104352 519726 104408
rect 519782 104352 519787 104408
rect 518788 104350 519787 104352
rect 519721 104347 519787 104350
rect 519629 103050 519695 103053
rect 518788 103048 519695 103050
rect 518788 102992 519634 103048
rect 519690 102992 519695 103048
rect 518788 102990 519695 102992
rect 519629 102987 519695 102990
rect 520733 103050 520799 103053
rect 523200 103050 524400 103080
rect 520733 103048 524400 103050
rect 520733 102992 520738 103048
rect 520794 102992 524400 103048
rect 520733 102990 524400 102992
rect 520733 102987 520799 102990
rect 523200 102960 524400 102990
rect 117037 102914 117103 102917
rect 117037 102912 119140 102914
rect 117037 102856 117042 102912
rect 117098 102856 119140 102912
rect 117037 102854 119140 102856
rect 117037 102851 117103 102854
rect 519537 101690 519603 101693
rect 518788 101688 519603 101690
rect 518788 101632 519542 101688
rect 519598 101632 519603 101688
rect 518788 101630 519603 101632
rect 519537 101627 519603 101630
rect 521469 101554 521535 101557
rect 523200 101554 524400 101584
rect 521469 101552 524400 101554
rect 521469 101496 521474 101552
rect 521530 101496 524400 101552
rect 521469 101494 524400 101496
rect 521469 101491 521535 101494
rect 523200 101464 524400 101494
rect 116945 101010 117011 101013
rect 116945 101008 119140 101010
rect 116945 100952 116950 101008
rect 117006 100952 119140 101008
rect 116945 100950 119140 100952
rect 116945 100947 117011 100950
rect 521101 100330 521167 100333
rect 518788 100328 521167 100330
rect 518788 100272 521106 100328
rect 521162 100272 521167 100328
rect 518788 100270 521167 100272
rect 521101 100267 521167 100270
rect 521377 100058 521443 100061
rect 523200 100058 524400 100088
rect 521377 100056 524400 100058
rect 521377 100000 521382 100056
rect 521438 100000 524400 100056
rect 521377 99998 524400 100000
rect 521377 99995 521443 99998
rect 523200 99968 524400 99998
rect 116853 99106 116919 99109
rect 116853 99104 119140 99106
rect 116853 99048 116858 99104
rect 116914 99048 119140 99104
rect 116853 99046 119140 99048
rect 116853 99043 116919 99046
rect 520825 98970 520891 98973
rect 518788 98968 520891 98970
rect 518788 98912 520830 98968
rect 520886 98912 520891 98968
rect 518788 98910 520891 98912
rect 520825 98907 520891 98910
rect 114093 98698 114159 98701
rect 110860 98696 114159 98698
rect 110860 98640 114098 98696
rect 114154 98640 114159 98696
rect 110860 98638 114159 98640
rect 114093 98635 114159 98638
rect 521285 98562 521351 98565
rect 523200 98562 524400 98592
rect 521285 98560 524400 98562
rect 521285 98504 521290 98560
rect 521346 98504 524400 98560
rect 521285 98502 524400 98504
rect 521285 98499 521351 98502
rect 523200 98472 524400 98502
rect 520273 97610 520339 97613
rect 518788 97608 520339 97610
rect 518788 97552 520278 97608
rect 520334 97552 520339 97608
rect 518788 97550 520339 97552
rect 520273 97547 520339 97550
rect 116761 97202 116827 97205
rect 116761 97200 119140 97202
rect 116761 97144 116766 97200
rect 116822 97144 119140 97200
rect 116761 97142 119140 97144
rect 116761 97139 116827 97142
rect 521101 97066 521167 97069
rect 523200 97066 524400 97096
rect 521101 97064 524400 97066
rect 521101 97008 521106 97064
rect 521162 97008 524400 97064
rect 521101 97006 524400 97008
rect 521101 97003 521167 97006
rect 523200 96976 524400 97006
rect 521009 96250 521075 96253
rect 518788 96248 521075 96250
rect 518788 96192 521014 96248
rect 521070 96192 521075 96248
rect 518788 96190 521075 96192
rect 521009 96187 521075 96190
rect 520273 95570 520339 95573
rect 523200 95570 524400 95600
rect 520273 95568 524400 95570
rect 520273 95512 520278 95568
rect 520334 95512 524400 95568
rect 520273 95510 524400 95512
rect 520273 95507 520339 95510
rect 523200 95480 524400 95510
rect 116669 95298 116735 95301
rect 116669 95296 119140 95298
rect 116669 95240 116674 95296
rect 116730 95240 119140 95296
rect 116669 95238 119140 95240
rect 116669 95235 116735 95238
rect 520733 94890 520799 94893
rect 518788 94888 520799 94890
rect 518788 94832 520738 94888
rect 520794 94832 520799 94888
rect 518788 94830 520799 94832
rect 520733 94827 520799 94830
rect 520917 93938 520983 93941
rect 523200 93938 524400 93968
rect 520917 93936 524400 93938
rect 520917 93880 520922 93936
rect 520978 93880 524400 93936
rect 520917 93878 524400 93880
rect 520917 93875 520983 93878
rect 523200 93848 524400 93878
rect 521469 93530 521535 93533
rect 518788 93528 521535 93530
rect 518788 93472 521474 93528
rect 521530 93472 521535 93528
rect 518788 93470 521535 93472
rect 521469 93467 521535 93470
rect 116577 93394 116643 93397
rect 116577 93392 119140 93394
rect 116577 93336 116582 93392
rect 116638 93336 119140 93392
rect 116577 93334 119140 93336
rect 116577 93331 116643 93334
rect 520181 92442 520247 92445
rect 523200 92442 524400 92472
rect 520181 92440 524400 92442
rect 520181 92384 520186 92440
rect 520242 92384 524400 92440
rect 520181 92382 524400 92384
rect 520181 92379 520247 92382
rect 523200 92352 524400 92382
rect 521377 92170 521443 92173
rect 518788 92168 521443 92170
rect 518788 92112 521382 92168
rect 521438 92112 521443 92168
rect 518788 92110 521443 92112
rect 521377 92107 521443 92110
rect 116117 91354 116183 91357
rect 116117 91352 119140 91354
rect 116117 91296 116122 91352
rect 116178 91296 119140 91352
rect 116117 91294 119140 91296
rect 116117 91291 116183 91294
rect 520089 90946 520155 90949
rect 523200 90946 524400 90976
rect 520089 90944 524400 90946
rect 520089 90888 520094 90944
rect 520150 90888 524400 90944
rect 520089 90886 524400 90888
rect 520089 90883 520155 90886
rect 523200 90856 524400 90886
rect 521285 90810 521351 90813
rect 518788 90808 521351 90810
rect 518788 90752 521290 90808
rect 521346 90752 521351 90808
rect 518788 90750 521351 90752
rect 521285 90747 521351 90750
rect 521101 89586 521167 89589
rect 518758 89584 521167 89586
rect 518758 89528 521106 89584
rect 521162 89528 521167 89584
rect 518758 89526 521167 89528
rect 116117 89450 116183 89453
rect 116117 89448 119140 89450
rect 116117 89392 116122 89448
rect 116178 89392 119140 89448
rect 518758 89420 518818 89526
rect 521101 89523 521167 89526
rect 519997 89450 520063 89453
rect 523200 89450 524400 89480
rect 519997 89448 524400 89450
rect 116117 89390 119140 89392
rect 519997 89392 520002 89448
rect 520058 89392 524400 89448
rect 519997 89390 524400 89392
rect 116117 89387 116183 89390
rect 519997 89387 520063 89390
rect 523200 89360 524400 89390
rect 520273 88090 520339 88093
rect 518788 88088 520339 88090
rect 518788 88032 520278 88088
rect 520334 88032 520339 88088
rect 518788 88030 520339 88032
rect 520273 88027 520339 88030
rect 519813 87954 519879 87957
rect 523200 87954 524400 87984
rect 519813 87952 524400 87954
rect 519813 87896 519818 87952
rect 519874 87896 524400 87952
rect 519813 87894 524400 87896
rect 519813 87891 519879 87894
rect 523200 87864 524400 87894
rect 116025 87546 116091 87549
rect 116025 87544 119140 87546
rect 116025 87488 116030 87544
rect 116086 87488 119140 87544
rect 116025 87486 119140 87488
rect 116025 87483 116091 87486
rect 114461 87274 114527 87277
rect 110860 87272 114527 87274
rect 110860 87216 114466 87272
rect 114522 87216 114527 87272
rect 110860 87214 114527 87216
rect 114461 87211 114527 87214
rect 520917 86730 520983 86733
rect 518788 86728 520983 86730
rect 518788 86672 520922 86728
rect 520978 86672 520983 86728
rect 518788 86670 520983 86672
rect 520917 86667 520983 86670
rect 519629 86458 519695 86461
rect 523200 86458 524400 86488
rect 519629 86456 524400 86458
rect 519629 86400 519634 86456
rect 519690 86400 524400 86456
rect 519629 86398 524400 86400
rect 519629 86395 519695 86398
rect 523200 86368 524400 86398
rect 115197 85642 115263 85645
rect 115197 85640 119140 85642
rect 115197 85584 115202 85640
rect 115258 85584 119140 85640
rect 115197 85582 119140 85584
rect 115197 85579 115263 85582
rect 520181 85370 520247 85373
rect 518788 85368 520247 85370
rect 518788 85312 520186 85368
rect 520242 85312 520247 85368
rect 518788 85310 520247 85312
rect 520181 85307 520247 85310
rect 519721 84962 519787 84965
rect 523200 84962 524400 84992
rect 519721 84960 524400 84962
rect 519721 84904 519726 84960
rect 519782 84904 524400 84960
rect 519721 84902 524400 84904
rect 519721 84899 519787 84902
rect 523200 84872 524400 84902
rect 520089 84010 520155 84013
rect 518788 84008 520155 84010
rect 518788 83952 520094 84008
rect 520150 83952 520155 84008
rect 518788 83950 520155 83952
rect 520089 83947 520155 83950
rect 116577 83738 116643 83741
rect 116577 83736 119140 83738
rect 116577 83680 116582 83736
rect 116638 83680 119140 83736
rect 116577 83678 119140 83680
rect 116577 83675 116643 83678
rect 519261 83466 519327 83469
rect 523200 83466 524400 83496
rect 519261 83464 524400 83466
rect 519261 83408 519266 83464
rect 519322 83408 524400 83464
rect 519261 83406 524400 83408
rect 519261 83403 519327 83406
rect 523200 83376 524400 83406
rect 519997 82650 520063 82653
rect 518788 82648 520063 82650
rect 518788 82592 520002 82648
rect 520058 82592 520063 82648
rect 518788 82590 520063 82592
rect 519997 82587 520063 82590
rect 519537 81970 519603 81973
rect 523200 81970 524400 82000
rect 519537 81968 524400 81970
rect 519537 81912 519542 81968
rect 519598 81912 524400 81968
rect 519537 81910 524400 81912
rect 519537 81907 519603 81910
rect 523200 81880 524400 81910
rect 116209 81834 116275 81837
rect 116209 81832 119140 81834
rect 116209 81776 116214 81832
rect 116270 81776 119140 81832
rect 116209 81774 119140 81776
rect 116209 81771 116275 81774
rect 519813 81290 519879 81293
rect 518788 81288 519879 81290
rect 518788 81232 519818 81288
rect 519874 81232 519879 81288
rect 518788 81230 519879 81232
rect 519813 81227 519879 81230
rect 519445 80474 519511 80477
rect 523200 80474 524400 80504
rect 519445 80472 524400 80474
rect 519445 80416 519450 80472
rect 519506 80416 524400 80472
rect 519445 80414 524400 80416
rect 519445 80411 519511 80414
rect 523200 80384 524400 80414
rect 115933 79930 115999 79933
rect 519629 79930 519695 79933
rect 115933 79928 119140 79930
rect 115933 79872 115938 79928
rect 115994 79872 119140 79928
rect 115933 79870 119140 79872
rect 518788 79928 519695 79930
rect 518788 79872 519634 79928
rect 519690 79872 519695 79928
rect 518788 79870 519695 79872
rect 115933 79867 115999 79870
rect 519629 79867 519695 79870
rect 519905 78978 519971 78981
rect 523200 78978 524400 79008
rect 519905 78976 524400 78978
rect 519905 78920 519910 78976
rect 519966 78920 524400 78976
rect 519905 78918 524400 78920
rect 519905 78915 519971 78918
rect 523200 78888 524400 78918
rect 519721 78570 519787 78573
rect 518788 78568 519787 78570
rect 518788 78512 519726 78568
rect 519782 78512 519787 78568
rect 518788 78510 519787 78512
rect 519721 78507 519787 78510
rect 116485 78026 116551 78029
rect 116485 78024 119140 78026
rect 116485 77968 116490 78024
rect 116546 77968 119140 78024
rect 116485 77966 119140 77968
rect 116485 77963 116551 77966
rect 519813 77482 519879 77485
rect 523200 77482 524400 77512
rect 519813 77480 524400 77482
rect 519813 77424 519818 77480
rect 519874 77424 524400 77480
rect 519813 77422 524400 77424
rect 519813 77419 519879 77422
rect 523200 77392 524400 77422
rect 519261 77210 519327 77213
rect 518788 77208 519327 77210
rect 518788 77152 519266 77208
rect 519322 77152 519327 77208
rect 518788 77150 519327 77152
rect 519261 77147 519327 77150
rect 519537 75986 519603 75989
rect 110860 75926 119140 75986
rect 518788 75984 519603 75986
rect 518788 75928 519542 75984
rect 519598 75928 519603 75984
rect 518788 75926 519603 75928
rect 519537 75923 519603 75926
rect 519721 75986 519787 75989
rect 523200 75986 524400 76016
rect 519721 75984 524400 75986
rect 519721 75928 519726 75984
rect 519782 75928 524400 75984
rect 519721 75926 524400 75928
rect 519721 75923 519787 75926
rect 523200 75896 524400 75926
rect 519445 74626 519511 74629
rect 518788 74624 519511 74626
rect 518788 74568 519450 74624
rect 519506 74568 519511 74624
rect 518788 74566 519511 74568
rect 519445 74563 519511 74566
rect 521009 74490 521075 74493
rect 523200 74490 524400 74520
rect 521009 74488 524400 74490
rect 521009 74432 521014 74488
rect 521070 74432 524400 74488
rect 521009 74430 524400 74432
rect 521009 74427 521075 74430
rect 523200 74400 524400 74430
rect 116669 74082 116735 74085
rect 116669 74080 119140 74082
rect 116669 74024 116674 74080
rect 116730 74024 119140 74080
rect 116669 74022 119140 74024
rect 116669 74019 116735 74022
rect 519905 73266 519971 73269
rect 518788 73264 519971 73266
rect 518788 73208 519910 73264
rect 519966 73208 519971 73264
rect 518788 73206 519971 73208
rect 519905 73203 519971 73206
rect 520917 72994 520983 72997
rect 523200 72994 524400 73024
rect 520917 72992 524400 72994
rect 520917 72936 520922 72992
rect 520978 72936 524400 72992
rect 520917 72934 524400 72936
rect 520917 72931 520983 72934
rect 523200 72904 524400 72934
rect 116577 72178 116643 72181
rect 116577 72176 119140 72178
rect 116577 72120 116582 72176
rect 116638 72120 119140 72176
rect 116577 72118 119140 72120
rect 116577 72115 116643 72118
rect 519813 71906 519879 71909
rect 518788 71904 519879 71906
rect 518788 71848 519818 71904
rect 519874 71848 519879 71904
rect 518788 71846 519879 71848
rect 519813 71843 519879 71846
rect 521193 71498 521259 71501
rect 523200 71498 524400 71528
rect 521193 71496 524400 71498
rect 521193 71440 521198 71496
rect 521254 71440 524400 71496
rect 521193 71438 524400 71440
rect 521193 71435 521259 71438
rect 523200 71408 524400 71438
rect 519721 70546 519787 70549
rect 518788 70544 519787 70546
rect 518788 70488 519726 70544
rect 519782 70488 519787 70544
rect 518788 70486 519787 70488
rect 519721 70483 519787 70486
rect 116301 70274 116367 70277
rect 116301 70272 119140 70274
rect 116301 70216 116306 70272
rect 116362 70216 119140 70272
rect 116301 70214 119140 70216
rect 116301 70211 116367 70214
rect 521101 69866 521167 69869
rect 523200 69866 524400 69896
rect 521101 69864 524400 69866
rect 521101 69808 521106 69864
rect 521162 69808 524400 69864
rect 521101 69806 524400 69808
rect 521101 69803 521167 69806
rect 523200 69776 524400 69806
rect 521009 69186 521075 69189
rect 518788 69184 521075 69186
rect 518788 69128 521014 69184
rect 521070 69128 521075 69184
rect 518788 69126 521075 69128
rect 521009 69123 521075 69126
rect 116117 68370 116183 68373
rect 521009 68370 521075 68373
rect 523200 68370 524400 68400
rect 116117 68368 119140 68370
rect 116117 68312 116122 68368
rect 116178 68312 119140 68368
rect 116117 68310 119140 68312
rect 521009 68368 524400 68370
rect 521009 68312 521014 68368
rect 521070 68312 524400 68368
rect 521009 68310 524400 68312
rect 116117 68307 116183 68310
rect 521009 68307 521075 68310
rect 523200 68280 524400 68310
rect 520917 67826 520983 67829
rect 518788 67824 520983 67826
rect 518788 67768 520922 67824
rect 520978 67768 520983 67824
rect 518788 67766 520983 67768
rect 520917 67763 520983 67766
rect 520457 66874 520523 66877
rect 523200 66874 524400 66904
rect 520457 66872 524400 66874
rect 520457 66816 520462 66872
rect 520518 66816 524400 66872
rect 520457 66814 524400 66816
rect 520457 66811 520523 66814
rect 523200 66784 524400 66814
rect 116577 66466 116643 66469
rect 521193 66466 521259 66469
rect 116577 66464 119140 66466
rect 116577 66408 116582 66464
rect 116638 66408 119140 66464
rect 116577 66406 119140 66408
rect 518788 66464 521259 66466
rect 518788 66408 521198 66464
rect 521254 66408 521259 66464
rect 518788 66406 521259 66408
rect 116577 66403 116643 66406
rect 521193 66403 521259 66406
rect 520365 65378 520431 65381
rect 523200 65378 524400 65408
rect 520365 65376 524400 65378
rect 520365 65320 520370 65376
rect 520426 65320 524400 65376
rect 520365 65318 524400 65320
rect 520365 65315 520431 65318
rect 523200 65288 524400 65318
rect 521101 65106 521167 65109
rect 518788 65104 521167 65106
rect 518788 65048 521106 65104
rect 521162 65048 521167 65104
rect 518788 65046 521167 65048
rect 521101 65043 521167 65046
rect 114461 64562 114527 64565
rect 110860 64560 114527 64562
rect 110860 64504 114466 64560
rect 114522 64504 114527 64560
rect 110860 64502 114527 64504
rect 114461 64499 114527 64502
rect 116209 64562 116275 64565
rect 116209 64560 119140 64562
rect 116209 64504 116214 64560
rect 116270 64504 119140 64560
rect 116209 64502 119140 64504
rect 116209 64499 116275 64502
rect 520733 63882 520799 63885
rect 523200 63882 524400 63912
rect 520733 63880 524400 63882
rect 520733 63824 520738 63880
rect 520794 63824 524400 63880
rect 520733 63822 524400 63824
rect 520733 63819 520799 63822
rect 523200 63792 524400 63822
rect 521009 63746 521075 63749
rect 518788 63744 521075 63746
rect 518788 63688 521014 63744
rect 521070 63688 521075 63744
rect 518788 63686 521075 63688
rect 521009 63683 521075 63686
rect 116577 62658 116643 62661
rect 116577 62656 119140 62658
rect 116577 62600 116582 62656
rect 116638 62600 119140 62656
rect 116577 62598 119140 62600
rect 116577 62595 116643 62598
rect 520457 62386 520523 62389
rect 518788 62384 520523 62386
rect 518788 62328 520462 62384
rect 520518 62328 520523 62384
rect 518788 62326 520523 62328
rect 520457 62323 520523 62326
rect 521009 62386 521075 62389
rect 523200 62386 524400 62416
rect 521009 62384 524400 62386
rect 521009 62328 521014 62384
rect 521070 62328 524400 62384
rect 521009 62326 524400 62328
rect 521009 62323 521075 62326
rect 523200 62296 524400 62326
rect 520365 61026 520431 61029
rect 518788 61024 520431 61026
rect 518788 60968 520370 61024
rect 520426 60968 520431 61024
rect 518788 60966 520431 60968
rect 520365 60963 520431 60966
rect 521101 60890 521167 60893
rect 523200 60890 524400 60920
rect 521101 60888 524400 60890
rect 521101 60832 521106 60888
rect 521162 60832 524400 60888
rect 521101 60830 524400 60832
rect 521101 60827 521167 60830
rect 523200 60800 524400 60830
rect 116669 60618 116735 60621
rect 116669 60616 119140 60618
rect 116669 60560 116674 60616
rect 116730 60560 119140 60616
rect 116669 60558 119140 60560
rect 116669 60555 116735 60558
rect 520733 59666 520799 59669
rect 518788 59664 520799 59666
rect 518788 59608 520738 59664
rect 520794 59608 520799 59664
rect 518788 59606 520799 59608
rect 520733 59603 520799 59606
rect 520733 59394 520799 59397
rect 523200 59394 524400 59424
rect 520733 59392 524400 59394
rect 520733 59336 520738 59392
rect 520794 59336 524400 59392
rect 520733 59334 524400 59336
rect 520733 59331 520799 59334
rect 523200 59304 524400 59334
rect 116761 58714 116827 58717
rect 116761 58712 119140 58714
rect 116761 58656 116766 58712
rect 116822 58656 119140 58712
rect 116761 58654 119140 58656
rect 116761 58651 116827 58654
rect 521009 58306 521075 58309
rect 518788 58304 521075 58306
rect 518788 58248 521014 58304
rect 521070 58248 521075 58304
rect 518788 58246 521075 58248
rect 521009 58243 521075 58246
rect 519905 57898 519971 57901
rect 523200 57898 524400 57928
rect 519905 57896 524400 57898
rect 519905 57840 519910 57896
rect 519966 57840 524400 57896
rect 519905 57838 524400 57840
rect 519905 57835 519971 57838
rect 523200 57808 524400 57838
rect 521101 56946 521167 56949
rect 518788 56944 521167 56946
rect 518788 56888 521106 56944
rect 521162 56888 521167 56944
rect 518788 56886 521167 56888
rect 521101 56883 521167 56886
rect 116853 56810 116919 56813
rect 116853 56808 119140 56810
rect 116853 56752 116858 56808
rect 116914 56752 119140 56808
rect 116853 56750 119140 56752
rect 116853 56747 116919 56750
rect 519813 56402 519879 56405
rect 523200 56402 524400 56432
rect 519813 56400 524400 56402
rect 519813 56344 519818 56400
rect 519874 56344 524400 56400
rect 519813 56342 524400 56344
rect 519813 56339 519879 56342
rect 523200 56312 524400 56342
rect 520733 55586 520799 55589
rect 518788 55584 520799 55586
rect 518788 55528 520738 55584
rect 520794 55528 520799 55584
rect 518788 55526 520799 55528
rect 520733 55523 520799 55526
rect 116945 54906 117011 54909
rect 519077 54906 519143 54909
rect 523200 54906 524400 54936
rect 116945 54904 119140 54906
rect 116945 54848 116950 54904
rect 117006 54848 119140 54904
rect 116945 54846 119140 54848
rect 519077 54904 524400 54906
rect 519077 54848 519082 54904
rect 519138 54848 524400 54904
rect 519077 54846 524400 54848
rect 116945 54843 117011 54846
rect 519077 54843 519143 54846
rect 523200 54816 524400 54846
rect 519905 54226 519971 54229
rect 518788 54224 519971 54226
rect 518788 54168 519910 54224
rect 519966 54168 519971 54224
rect 518788 54166 519971 54168
rect 519905 54163 519971 54166
rect 520181 53410 520247 53413
rect 523200 53410 524400 53440
rect 520181 53408 524400 53410
rect 520181 53352 520186 53408
rect 520242 53352 524400 53408
rect 520181 53350 524400 53352
rect 520181 53347 520247 53350
rect 523200 53320 524400 53350
rect 114185 53138 114251 53141
rect 110860 53136 114251 53138
rect 110860 53080 114190 53136
rect 114246 53080 114251 53136
rect 110860 53078 114251 53080
rect 114185 53075 114251 53078
rect 117037 53002 117103 53005
rect 117037 53000 119140 53002
rect 117037 52944 117042 53000
rect 117098 52944 119140 53000
rect 117037 52942 119140 52944
rect 117037 52939 117103 52942
rect 519813 52866 519879 52869
rect 518788 52864 519879 52866
rect 518788 52808 519818 52864
rect 519874 52808 519879 52864
rect 518788 52806 519879 52808
rect 519813 52803 519879 52806
rect 520089 51914 520155 51917
rect 523200 51914 524400 51944
rect 520089 51912 524400 51914
rect 520089 51856 520094 51912
rect 520150 51856 524400 51912
rect 520089 51854 524400 51856
rect 520089 51851 520155 51854
rect 523200 51824 524400 51854
rect 519077 51506 519143 51509
rect 518788 51504 519143 51506
rect 518788 51448 519082 51504
rect 519138 51448 519143 51504
rect 518788 51446 519143 51448
rect 519077 51443 519143 51446
rect 117129 51098 117195 51101
rect 117129 51096 119140 51098
rect 117129 51040 117134 51096
rect 117190 51040 119140 51096
rect 117129 51038 119140 51040
rect 117129 51035 117195 51038
rect 519077 50418 519143 50421
rect 523200 50418 524400 50448
rect 519077 50416 524400 50418
rect 519077 50360 519082 50416
rect 519138 50360 524400 50416
rect 519077 50358 524400 50360
rect 519077 50355 519143 50358
rect 523200 50328 524400 50358
rect 520181 50146 520247 50149
rect 518788 50144 520247 50146
rect 518788 50088 520186 50144
rect 520242 50088 520247 50144
rect 518788 50086 520247 50088
rect 520181 50083 520247 50086
rect 117221 49194 117287 49197
rect 117221 49192 119140 49194
rect 117221 49136 117226 49192
rect 117282 49136 119140 49192
rect 117221 49134 119140 49136
rect 117221 49131 117287 49134
rect 520181 48922 520247 48925
rect 523200 48922 524400 48952
rect 520181 48920 524400 48922
rect 520181 48864 520186 48920
rect 520242 48864 524400 48920
rect 520181 48862 524400 48864
rect 520181 48859 520247 48862
rect 523200 48832 524400 48862
rect 520089 48786 520155 48789
rect 518788 48784 520155 48786
rect 518788 48728 520094 48784
rect 520150 48728 520155 48784
rect 518788 48726 520155 48728
rect 520089 48723 520155 48726
rect 519077 47426 519143 47429
rect 518788 47424 519143 47426
rect 518788 47368 519082 47424
rect 519138 47368 519143 47424
rect 518788 47366 519143 47368
rect 519077 47363 519143 47366
rect 519445 47290 519511 47293
rect 523200 47290 524400 47320
rect 519445 47288 524400 47290
rect 519445 47232 519450 47288
rect 519506 47232 524400 47288
rect 519445 47230 524400 47232
rect 519445 47227 519511 47230
rect 523200 47200 524400 47230
rect 116485 47154 116551 47157
rect 116485 47152 119140 47154
rect 116485 47096 116490 47152
rect 116546 47096 119140 47152
rect 116485 47094 119140 47096
rect 116485 47091 116551 47094
rect 520181 46066 520247 46069
rect 518788 46064 520247 46066
rect 518788 46008 520186 46064
rect 520242 46008 520247 46064
rect 518788 46006 520247 46008
rect 520181 46003 520247 46006
rect 519721 45794 519787 45797
rect 523200 45794 524400 45824
rect 519721 45792 524400 45794
rect 519721 45736 519726 45792
rect 519782 45736 524400 45792
rect 519721 45734 524400 45736
rect 519721 45731 519787 45734
rect 523200 45704 524400 45734
rect 116209 45250 116275 45253
rect 116209 45248 119140 45250
rect 116209 45192 116214 45248
rect 116270 45192 119140 45248
rect 116209 45190 119140 45192
rect 116209 45187 116275 45190
rect 519445 44706 519511 44709
rect 518788 44704 519511 44706
rect 518788 44648 519450 44704
rect 519506 44648 519511 44704
rect 518788 44646 519511 44648
rect 519445 44643 519511 44646
rect 520181 44298 520247 44301
rect 523200 44298 524400 44328
rect 520181 44296 524400 44298
rect 520181 44240 520186 44296
rect 520242 44240 524400 44296
rect 520181 44238 524400 44240
rect 520181 44235 520247 44238
rect 523200 44208 524400 44238
rect 116301 43346 116367 43349
rect 519721 43346 519787 43349
rect 116301 43344 119140 43346
rect 116301 43288 116306 43344
rect 116362 43288 119140 43344
rect 116301 43286 119140 43288
rect 518788 43344 519787 43346
rect 518788 43288 519726 43344
rect 519782 43288 519787 43344
rect 518788 43286 519787 43288
rect 116301 43283 116367 43286
rect 519721 43283 519787 43286
rect 520733 42802 520799 42805
rect 523200 42802 524400 42832
rect 520733 42800 524400 42802
rect 520733 42744 520738 42800
rect 520794 42744 524400 42800
rect 520733 42742 524400 42744
rect 520733 42739 520799 42742
rect 523200 42712 524400 42742
rect 520181 41986 520247 41989
rect 518788 41984 520247 41986
rect 518788 41928 520186 41984
rect 520242 41928 520247 41984
rect 518788 41926 520247 41928
rect 520181 41923 520247 41926
rect 114093 41850 114159 41853
rect 110860 41848 114159 41850
rect 110860 41792 114098 41848
rect 114154 41792 114159 41848
rect 110860 41790 114159 41792
rect 114093 41787 114159 41790
rect 116117 41442 116183 41445
rect 116117 41440 119140 41442
rect 116117 41384 116122 41440
rect 116178 41384 119140 41440
rect 116117 41382 119140 41384
rect 116117 41379 116183 41382
rect 520733 41306 520799 41309
rect 518758 41304 520799 41306
rect 518758 41248 520738 41304
rect 520794 41248 520799 41304
rect 518758 41246 520799 41248
rect 518758 40596 518818 41246
rect 520733 41243 520799 41246
rect 520917 41306 520983 41309
rect 523200 41306 524400 41336
rect 520917 41304 524400 41306
rect 520917 41248 520922 41304
rect 520978 41248 524400 41304
rect 520917 41246 524400 41248
rect 520917 41243 520983 41246
rect 523200 41216 524400 41246
rect 520917 39946 520983 39949
rect 518758 39944 520983 39946
rect 518758 39888 520922 39944
rect 520978 39888 520983 39944
rect 518758 39886 520983 39888
rect 116393 39538 116459 39541
rect 116393 39536 119140 39538
rect 116393 39480 116398 39536
rect 116454 39480 119140 39536
rect 116393 39478 119140 39480
rect 116393 39475 116459 39478
rect 518758 39236 518818 39886
rect 520917 39883 520983 39886
rect 520917 39810 520983 39813
rect 523200 39810 524400 39840
rect 520917 39808 524400 39810
rect 520917 39752 520922 39808
rect 520978 39752 524400 39808
rect 520917 39750 524400 39752
rect 520917 39747 520983 39750
rect 523200 39720 524400 39750
rect 521101 38314 521167 38317
rect 523200 38314 524400 38344
rect 521101 38312 524400 38314
rect 521101 38256 521106 38312
rect 521162 38256 524400 38312
rect 521101 38254 524400 38256
rect 521101 38251 521167 38254
rect 523200 38224 524400 38254
rect 520917 37906 520983 37909
rect 518788 37904 520983 37906
rect 518788 37848 520922 37904
rect 520978 37848 520983 37904
rect 518788 37846 520983 37848
rect 520917 37843 520983 37846
rect 116209 37634 116275 37637
rect 116209 37632 119140 37634
rect 116209 37576 116214 37632
rect 116270 37576 119140 37632
rect 116209 37574 119140 37576
rect 116209 37571 116275 37574
rect 521101 37226 521167 37229
rect 518758 37224 521167 37226
rect 518758 37168 521106 37224
rect 521162 37168 521167 37224
rect 518758 37166 521167 37168
rect 518758 36516 518818 37166
rect 521101 37163 521167 37166
rect 521561 36818 521627 36821
rect 523200 36818 524400 36848
rect 521561 36816 524400 36818
rect 521561 36760 521566 36816
rect 521622 36760 524400 36816
rect 521561 36758 524400 36760
rect 521561 36755 521627 36758
rect 523200 36728 524400 36758
rect 521561 36002 521627 36005
rect 521561 36000 521670 36002
rect 521561 35944 521566 36000
rect 521622 35944 521670 36000
rect 521561 35939 521670 35944
rect 521610 35866 521670 35939
rect 518758 35806 521670 35866
rect 116117 35730 116183 35733
rect 116117 35728 119140 35730
rect 116117 35672 116122 35728
rect 116178 35672 119140 35728
rect 116117 35670 119140 35672
rect 116117 35667 116183 35670
rect 518758 35156 518818 35806
rect 520917 35322 520983 35325
rect 523200 35322 524400 35352
rect 520917 35320 524400 35322
rect 520917 35264 520922 35320
rect 520978 35264 524400 35320
rect 520917 35262 524400 35264
rect 520917 35259 520983 35262
rect 523200 35232 524400 35262
rect 520917 34506 520983 34509
rect 518758 34504 520983 34506
rect 518758 34448 520922 34504
rect 520978 34448 520983 34504
rect 518758 34446 520983 34448
rect 116117 33826 116183 33829
rect 116117 33824 119140 33826
rect 116117 33768 116122 33824
rect 116178 33768 119140 33824
rect 518758 33796 518818 34446
rect 520917 34443 520983 34446
rect 521101 33826 521167 33829
rect 523200 33826 524400 33856
rect 521101 33824 524400 33826
rect 116117 33766 119140 33768
rect 521101 33768 521106 33824
rect 521162 33768 524400 33824
rect 521101 33766 524400 33768
rect 116117 33763 116183 33766
rect 521101 33763 521167 33766
rect 523200 33736 524400 33766
rect 521101 33146 521167 33149
rect 518758 33144 521167 33146
rect 518758 33088 521106 33144
rect 521162 33088 521167 33144
rect 518758 33086 521167 33088
rect 518758 32436 518818 33086
rect 521101 33083 521167 33086
rect 521101 32330 521167 32333
rect 523200 32330 524400 32360
rect 521101 32328 524400 32330
rect 521101 32272 521106 32328
rect 521162 32272 524400 32328
rect 521101 32270 524400 32272
rect 521101 32267 521167 32270
rect 523200 32240 524400 32270
rect 116117 31786 116183 31789
rect 116117 31784 119140 31786
rect 116117 31728 116122 31784
rect 116178 31728 119140 31784
rect 116117 31726 119140 31728
rect 116117 31723 116183 31726
rect 521101 31650 521167 31653
rect 518758 31648 521167 31650
rect 518758 31592 521106 31648
rect 521162 31592 521167 31648
rect 518758 31590 521167 31592
rect 518758 31076 518818 31590
rect 521101 31587 521167 31590
rect 523200 30834 524400 30864
rect 518850 30774 524400 30834
rect 114001 30426 114067 30429
rect 110860 30424 114067 30426
rect 110860 30368 114006 30424
rect 114062 30368 114067 30424
rect 110860 30366 114067 30368
rect 114001 30363 114067 30366
rect 518850 30290 518910 30774
rect 523200 30744 524400 30774
rect 518758 30230 518910 30290
rect 116117 29882 116183 29885
rect 116117 29880 119140 29882
rect 116117 29824 116122 29880
rect 116178 29824 119140 29880
rect 116117 29822 119140 29824
rect 116117 29819 116183 29822
rect 518758 29716 518818 30230
rect 520917 29338 520983 29341
rect 523200 29338 524400 29368
rect 520917 29336 524400 29338
rect 520917 29280 520922 29336
rect 520978 29280 524400 29336
rect 520917 29278 524400 29280
rect 520917 29275 520983 29278
rect 523200 29248 524400 29278
rect 520917 28386 520983 28389
rect 518788 28384 520983 28386
rect 518788 28328 520922 28384
rect 520978 28328 520983 28384
rect 518788 28326 520983 28328
rect 520917 28323 520983 28326
rect 116117 27978 116183 27981
rect 116117 27976 119140 27978
rect 116117 27920 116122 27976
rect 116178 27920 119140 27976
rect 116117 27918 119140 27920
rect 116117 27915 116183 27918
rect 523200 27842 524400 27872
rect 518850 27782 524400 27842
rect 518850 27570 518910 27782
rect 523200 27752 524400 27782
rect 518758 27510 518910 27570
rect 518758 26996 518818 27510
rect 523200 26346 524400 26376
rect 521610 26286 524400 26346
rect 521610 26210 521670 26286
rect 523200 26256 524400 26286
rect 518758 26150 521670 26210
rect 116117 26074 116183 26077
rect 116117 26072 119140 26074
rect 116117 26016 116122 26072
rect 116178 26016 119140 26072
rect 116117 26014 119140 26016
rect 116117 26011 116183 26014
rect 518758 25636 518818 26150
rect 521101 24850 521167 24853
rect 523200 24850 524400 24880
rect 521101 24848 524400 24850
rect 521101 24792 521106 24848
rect 521162 24792 524400 24848
rect 521101 24790 524400 24792
rect 521101 24787 521167 24790
rect 523200 24760 524400 24790
rect 116117 24170 116183 24173
rect 116117 24168 119140 24170
rect 116117 24112 116122 24168
rect 116178 24112 119140 24168
rect 116117 24110 119140 24112
rect 116117 24107 116183 24110
rect 518758 23626 518818 24276
rect 521101 23626 521167 23629
rect 518758 23624 521167 23626
rect 518758 23568 521106 23624
rect 521162 23568 521167 23624
rect 518758 23566 521167 23568
rect 521101 23563 521167 23566
rect 520365 23218 520431 23221
rect 523200 23218 524400 23248
rect 520365 23216 524400 23218
rect 520365 23160 520370 23216
rect 520426 23160 524400 23216
rect 520365 23158 524400 23160
rect 520365 23155 520431 23158
rect 523200 23128 524400 23158
rect 116025 22266 116091 22269
rect 518758 22266 518818 22916
rect 520365 22266 520431 22269
rect 116025 22264 119140 22266
rect 116025 22208 116030 22264
rect 116086 22208 119140 22264
rect 116025 22206 119140 22208
rect 518758 22264 520431 22266
rect 518758 22208 520370 22264
rect 520426 22208 520431 22264
rect 518758 22206 520431 22208
rect 116025 22203 116091 22206
rect 520365 22203 520431 22206
rect 520917 21722 520983 21725
rect 523200 21722 524400 21752
rect 520917 21720 524400 21722
rect 520917 21664 520922 21720
rect 520978 21664 524400 21720
rect 520917 21662 524400 21664
rect 520917 21659 520983 21662
rect 523200 21632 524400 21662
rect 518758 20906 518818 21556
rect 520917 20906 520983 20909
rect 518758 20904 520983 20906
rect 518758 20848 520922 20904
rect 520978 20848 520983 20904
rect 518758 20846 520983 20848
rect 520917 20843 520983 20846
rect 116209 20362 116275 20365
rect 116209 20360 119140 20362
rect 116209 20304 116214 20360
rect 116270 20304 119140 20360
rect 116209 20302 119140 20304
rect 116209 20299 116275 20302
rect 521101 20226 521167 20229
rect 523200 20226 524400 20256
rect 521101 20224 524400 20226
rect 518758 19546 518818 20196
rect 521101 20168 521106 20224
rect 521162 20168 524400 20224
rect 521101 20166 524400 20168
rect 521101 20163 521167 20166
rect 523200 20136 524400 20166
rect 521101 19546 521167 19549
rect 518758 19544 521167 19546
rect 518758 19488 521106 19544
rect 521162 19488 521167 19544
rect 518758 19486 521167 19488
rect 521101 19483 521167 19486
rect 113909 19002 113975 19005
rect 110860 19000 113975 19002
rect 110860 18944 113914 19000
rect 113970 18944 113975 19000
rect 110860 18942 113975 18944
rect 113909 18939 113975 18942
rect 116117 18458 116183 18461
rect 116117 18456 119140 18458
rect 116117 18400 116122 18456
rect 116178 18400 119140 18456
rect 116117 18398 119140 18400
rect 116117 18395 116183 18398
rect 518758 18186 518818 18836
rect 523200 18730 524400 18760
rect 521150 18670 524400 18730
rect 521150 18186 521210 18670
rect 523200 18640 524400 18670
rect 518758 18126 521210 18186
rect 518758 16826 518818 17476
rect 523200 17234 524400 17264
rect 521150 17174 524400 17234
rect 521150 16826 521210 17174
rect 523200 17144 524400 17174
rect 518758 16766 521210 16826
rect 116209 16418 116275 16421
rect 116209 16416 119140 16418
rect 116209 16360 116214 16416
rect 116270 16360 119140 16416
rect 116209 16358 119140 16360
rect 116209 16355 116275 16358
rect 518758 15466 518818 16116
rect 523200 15738 524400 15768
rect 521150 15678 524400 15738
rect 521150 15466 521210 15678
rect 523200 15648 524400 15678
rect 518758 15406 521210 15466
rect 115933 14514 115999 14517
rect 115933 14512 119140 14514
rect 115933 14456 115938 14512
rect 115994 14456 119140 14512
rect 115933 14454 119140 14456
rect 115933 14451 115999 14454
rect 523200 14152 524400 14272
rect 523200 12656 524400 12776
rect 116526 12548 116532 12612
rect 116596 12610 116602 12612
rect 116596 12550 119140 12610
rect 116596 12548 116602 12550
rect 523200 11160 524400 11280
rect 116710 10644 116716 10708
rect 116780 10706 116786 10708
rect 116780 10646 119140 10706
rect 116780 10644 116786 10646
rect 523200 9664 524400 9784
rect 117262 8740 117268 8804
rect 117332 8802 117338 8804
rect 117332 8742 119140 8802
rect 117332 8740 117338 8742
rect 523200 8168 524400 8288
rect 113817 7714 113883 7717
rect 110860 7712 113883 7714
rect 110860 7656 113822 7712
rect 113878 7656 113883 7712
rect 110860 7654 113883 7656
rect 113817 7651 113883 7654
rect 116158 6836 116164 6900
rect 116228 6898 116234 6900
rect 116228 6838 119140 6898
rect 116228 6836 116234 6838
rect 523200 6672 524400 6792
rect 523200 5176 524400 5296
rect 116117 4994 116183 4997
rect 116117 4992 119140 4994
rect 116117 4936 116122 4992
rect 116178 4936 119140 4992
rect 116117 4934 119140 4936
rect 116117 4931 116183 4934
rect 523200 3680 524400 3800
rect 116117 3090 116183 3093
rect 116117 3088 119140 3090
rect 116117 3032 116122 3088
rect 116178 3032 119140 3088
rect 116117 3030 119140 3032
rect 116117 3027 116183 3030
rect 53649 2682 53715 2685
rect 82997 2682 83063 2685
rect 53649 2680 83063 2682
rect 53649 2624 53654 2680
rect 53710 2624 83002 2680
rect 83058 2624 83063 2680
rect 53649 2622 83063 2624
rect 53649 2619 53715 2622
rect 82997 2619 83063 2622
rect 58709 2546 58775 2549
rect 82077 2546 82143 2549
rect 58709 2544 82143 2546
rect 58709 2488 58714 2544
rect 58770 2488 82082 2544
rect 82138 2488 82143 2544
rect 58709 2486 82143 2488
rect 58709 2483 58775 2486
rect 82077 2483 82143 2486
rect 82353 2546 82419 2549
rect 83089 2546 83155 2549
rect 82353 2544 83155 2546
rect 82353 2488 82358 2544
rect 82414 2488 83094 2544
rect 83150 2488 83155 2544
rect 82353 2486 83155 2488
rect 82353 2483 82419 2486
rect 83089 2483 83155 2486
rect 56133 2410 56199 2413
rect 63493 2410 63559 2413
rect 56133 2408 63559 2410
rect 56133 2352 56138 2408
rect 56194 2352 63498 2408
rect 63554 2352 63559 2408
rect 56133 2350 63559 2352
rect 56133 2347 56199 2350
rect 63493 2347 63559 2350
rect 66345 2410 66411 2413
rect 82721 2410 82787 2413
rect 66345 2408 82787 2410
rect 66345 2352 66350 2408
rect 66406 2352 82726 2408
rect 82782 2352 82787 2408
rect 66345 2350 82787 2352
rect 66345 2347 66411 2350
rect 82721 2347 82787 2350
rect 523200 2184 524400 2304
rect 19333 1866 19399 1869
rect 116526 1866 116532 1868
rect 19333 1864 116532 1866
rect 19333 1808 19338 1864
rect 19394 1808 116532 1864
rect 19333 1806 116532 1808
rect 19333 1803 19399 1806
rect 116526 1804 116532 1806
rect 116596 1804 116602 1868
rect 15929 1730 15995 1733
rect 116710 1730 116716 1732
rect 15929 1728 116716 1730
rect 15929 1672 15934 1728
rect 15990 1672 116716 1728
rect 15929 1670 116716 1672
rect 15929 1667 15995 1670
rect 116710 1668 116716 1670
rect 116780 1668 116786 1732
rect 12617 1594 12683 1597
rect 117262 1594 117268 1596
rect 12617 1592 117268 1594
rect 12617 1536 12622 1592
rect 12678 1536 117268 1592
rect 12617 1534 117268 1536
rect 12617 1531 12683 1534
rect 117262 1532 117268 1534
rect 117332 1532 117338 1596
rect 229277 1594 229343 1597
rect 293585 1594 293651 1597
rect 229277 1592 293651 1594
rect 229277 1536 229282 1592
rect 229338 1536 293590 1592
rect 293646 1536 293651 1592
rect 229277 1534 293651 1536
rect 229277 1531 229343 1534
rect 293585 1531 293651 1534
rect 9305 1458 9371 1461
rect 116158 1458 116164 1460
rect 9305 1456 116164 1458
rect 9305 1400 9310 1456
rect 9366 1400 116164 1456
rect 9305 1398 116164 1400
rect 9305 1395 9371 1398
rect 116158 1396 116164 1398
rect 116228 1396 116234 1460
rect 163773 1458 163839 1461
rect 243629 1458 243695 1461
rect 163773 1456 243695 1458
rect 163773 1400 163778 1456
rect 163834 1400 243634 1456
rect 243690 1400 243695 1456
rect 163773 1398 243695 1400
rect 163773 1395 163839 1398
rect 243629 1395 243695 1398
rect 360285 1458 360351 1461
rect 393589 1458 393655 1461
rect 360285 1456 393655 1458
rect 360285 1400 360290 1456
rect 360346 1400 393594 1456
rect 393650 1400 393655 1456
rect 360285 1398 393655 1400
rect 360285 1395 360351 1398
rect 393589 1395 393655 1398
rect 523200 688 524400 808
<< via3 >>
rect 116532 12548 116596 12612
rect 116716 10644 116780 10708
rect 117268 8740 117332 8804
rect 116164 6836 116228 6900
rect 116532 1804 116596 1868
rect 116716 1668 116780 1732
rect 117268 1532 117332 1596
rect 116164 1396 116228 1460
<< metal4 >>
rect 1664 144454 1984 144496
rect 1664 144218 1706 144454
rect 1942 144218 1984 144454
rect 1664 144134 1984 144218
rect 1664 143898 1706 144134
rect 1942 143898 1984 144134
rect 1664 143856 1984 143898
rect 109956 144454 110276 144496
rect 109956 144218 109998 144454
rect 110234 144218 110276 144454
rect 109956 144134 110276 144218
rect 109956 143898 109998 144134
rect 110234 143898 110276 144134
rect 109956 143856 110276 143898
rect 119664 144454 119984 144496
rect 119664 144218 119706 144454
rect 119942 144218 119984 144454
rect 119664 144134 119984 144218
rect 119664 143898 119706 144134
rect 119942 143898 119984 144134
rect 119664 143856 119984 143898
rect 517940 144454 518260 144496
rect 517940 144218 517982 144454
rect 518218 144218 518260 144454
rect 517940 144134 518260 144218
rect 517940 143898 517982 144134
rect 518218 143898 518260 144134
rect 517940 143856 518260 143898
rect 1096 131454 1332 131496
rect 1096 131134 1332 131218
rect 1096 130856 1332 130898
rect 110616 131454 110936 131496
rect 110616 131218 110658 131454
rect 110894 131218 110936 131454
rect 110616 131134 110936 131218
rect 110616 130898 110658 131134
rect 110894 130898 110936 131134
rect 110616 130856 110936 130898
rect 119004 131454 119324 131496
rect 119004 131218 119046 131454
rect 119282 131218 119324 131454
rect 119004 131134 119324 131218
rect 119004 130898 119046 131134
rect 119282 130898 119324 131134
rect 119004 130856 119324 130898
rect 518600 131454 518920 131496
rect 518600 131218 518642 131454
rect 518878 131218 518920 131454
rect 518600 131134 518920 131218
rect 518600 130898 518642 131134
rect 518878 130898 518920 131134
rect 518600 130856 518920 130898
rect 1664 118454 1984 118496
rect 1664 118218 1706 118454
rect 1942 118218 1984 118454
rect 1664 118134 1984 118218
rect 1664 117898 1706 118134
rect 1942 117898 1984 118134
rect 1664 117856 1984 117898
rect 109956 118454 110276 118496
rect 109956 118218 109998 118454
rect 110234 118218 110276 118454
rect 109956 118134 110276 118218
rect 109956 117898 109998 118134
rect 110234 117898 110276 118134
rect 109956 117856 110276 117898
rect 119664 118454 119984 118496
rect 119664 118218 119706 118454
rect 119942 118218 119984 118454
rect 119664 118134 119984 118218
rect 119664 117898 119706 118134
rect 119942 117898 119984 118134
rect 119664 117856 119984 117898
rect 517940 118454 518260 118496
rect 517940 118218 517982 118454
rect 518218 118218 518260 118454
rect 517940 118134 518260 118218
rect 517940 117898 517982 118134
rect 518218 117898 518260 118134
rect 517940 117856 518260 117898
rect 1096 105454 1332 105496
rect 1096 105134 1332 105218
rect 1096 104856 1332 104898
rect 110616 105454 110936 105496
rect 110616 105218 110658 105454
rect 110894 105218 110936 105454
rect 110616 105134 110936 105218
rect 110616 104898 110658 105134
rect 110894 104898 110936 105134
rect 110616 104856 110936 104898
rect 119004 105454 119324 105496
rect 119004 105218 119046 105454
rect 119282 105218 119324 105454
rect 119004 105134 119324 105218
rect 119004 104898 119046 105134
rect 119282 104898 119324 105134
rect 119004 104856 119324 104898
rect 518600 105454 518920 105496
rect 518600 105218 518642 105454
rect 518878 105218 518920 105454
rect 518600 105134 518920 105218
rect 518600 104898 518642 105134
rect 518878 104898 518920 105134
rect 518600 104856 518920 104898
rect 1664 92454 1984 92496
rect 1664 92218 1706 92454
rect 1942 92218 1984 92454
rect 1664 92134 1984 92218
rect 1664 91898 1706 92134
rect 1942 91898 1984 92134
rect 1664 91856 1984 91898
rect 109956 92454 110276 92496
rect 109956 92218 109998 92454
rect 110234 92218 110276 92454
rect 109956 92134 110276 92218
rect 109956 91898 109998 92134
rect 110234 91898 110276 92134
rect 109956 91856 110276 91898
rect 119664 92454 119984 92496
rect 119664 92218 119706 92454
rect 119942 92218 119984 92454
rect 119664 92134 119984 92218
rect 119664 91898 119706 92134
rect 119942 91898 119984 92134
rect 119664 91856 119984 91898
rect 517940 92454 518260 92496
rect 517940 92218 517982 92454
rect 518218 92218 518260 92454
rect 517940 92134 518260 92218
rect 517940 91898 517982 92134
rect 518218 91898 518260 92134
rect 517940 91856 518260 91898
rect 1096 79454 1332 79496
rect 1096 79134 1332 79218
rect 1096 78856 1332 78898
rect 110616 79454 110936 79496
rect 110616 79218 110658 79454
rect 110894 79218 110936 79454
rect 110616 79134 110936 79218
rect 110616 78898 110658 79134
rect 110894 78898 110936 79134
rect 110616 78856 110936 78898
rect 119004 79454 119324 79496
rect 119004 79218 119046 79454
rect 119282 79218 119324 79454
rect 119004 79134 119324 79218
rect 119004 78898 119046 79134
rect 119282 78898 119324 79134
rect 119004 78856 119324 78898
rect 518600 79454 518920 79496
rect 518600 79218 518642 79454
rect 518878 79218 518920 79454
rect 518600 79134 518920 79218
rect 518600 78898 518642 79134
rect 518878 78898 518920 79134
rect 518600 78856 518920 78898
rect 1664 66454 1984 66496
rect 1664 66218 1706 66454
rect 1942 66218 1984 66454
rect 1664 66134 1984 66218
rect 1664 65898 1706 66134
rect 1942 65898 1984 66134
rect 1664 65856 1984 65898
rect 109956 66454 110276 66496
rect 109956 66218 109998 66454
rect 110234 66218 110276 66454
rect 109956 66134 110276 66218
rect 109956 65898 109998 66134
rect 110234 65898 110276 66134
rect 109956 65856 110276 65898
rect 119664 66454 119984 66496
rect 119664 66218 119706 66454
rect 119942 66218 119984 66454
rect 119664 66134 119984 66218
rect 119664 65898 119706 66134
rect 119942 65898 119984 66134
rect 119664 65856 119984 65898
rect 517940 66454 518260 66496
rect 517940 66218 517982 66454
rect 518218 66218 518260 66454
rect 517940 66134 518260 66218
rect 517940 65898 517982 66134
rect 518218 65898 518260 66134
rect 517940 65856 518260 65898
rect 1096 53454 1332 53496
rect 1096 53134 1332 53218
rect 1096 52856 1332 52898
rect 110616 53454 110936 53496
rect 110616 53218 110658 53454
rect 110894 53218 110936 53454
rect 110616 53134 110936 53218
rect 110616 52898 110658 53134
rect 110894 52898 110936 53134
rect 110616 52856 110936 52898
rect 119004 53454 119324 53496
rect 119004 53218 119046 53454
rect 119282 53218 119324 53454
rect 119004 53134 119324 53218
rect 119004 52898 119046 53134
rect 119282 52898 119324 53134
rect 119004 52856 119324 52898
rect 518600 53454 518920 53496
rect 518600 53218 518642 53454
rect 518878 53218 518920 53454
rect 518600 53134 518920 53218
rect 518600 52898 518642 53134
rect 518878 52898 518920 53134
rect 518600 52856 518920 52898
rect 1664 40454 1984 40496
rect 1664 40218 1706 40454
rect 1942 40218 1984 40454
rect 1664 40134 1984 40218
rect 1664 39898 1706 40134
rect 1942 39898 1984 40134
rect 1664 39856 1984 39898
rect 109956 40454 110276 40496
rect 109956 40218 109998 40454
rect 110234 40218 110276 40454
rect 109956 40134 110276 40218
rect 109956 39898 109998 40134
rect 110234 39898 110276 40134
rect 109956 39856 110276 39898
rect 119664 40454 119984 40496
rect 119664 40218 119706 40454
rect 119942 40218 119984 40454
rect 119664 40134 119984 40218
rect 119664 39898 119706 40134
rect 119942 39898 119984 40134
rect 119664 39856 119984 39898
rect 517940 40454 518260 40496
rect 517940 40218 517982 40454
rect 518218 40218 518260 40454
rect 517940 40134 518260 40218
rect 517940 39898 517982 40134
rect 518218 39898 518260 40134
rect 517940 39856 518260 39898
rect 1096 27454 1332 27496
rect 1096 27134 1332 27218
rect 1096 26856 1332 26898
rect 110616 27454 110936 27496
rect 110616 27218 110658 27454
rect 110894 27218 110936 27454
rect 110616 27134 110936 27218
rect 110616 26898 110658 27134
rect 110894 26898 110936 27134
rect 110616 26856 110936 26898
rect 119004 27454 119324 27496
rect 119004 27218 119046 27454
rect 119282 27218 119324 27454
rect 119004 27134 119324 27218
rect 119004 26898 119046 27134
rect 119282 26898 119324 27134
rect 119004 26856 119324 26898
rect 518600 27454 518920 27496
rect 518600 27218 518642 27454
rect 518878 27218 518920 27454
rect 518600 27134 518920 27218
rect 518600 26898 518642 27134
rect 518878 26898 518920 27134
rect 518600 26856 518920 26898
rect 1664 14454 1984 14496
rect 1664 14218 1706 14454
rect 1942 14218 1984 14454
rect 1664 14134 1984 14218
rect 1664 13898 1706 14134
rect 1942 13898 1984 14134
rect 1664 13856 1984 13898
rect 109956 14454 110276 14496
rect 109956 14218 109998 14454
rect 110234 14218 110276 14454
rect 109956 14134 110276 14218
rect 109956 13898 109998 14134
rect 110234 13898 110276 14134
rect 109956 13856 110276 13898
rect 119664 14454 119984 14496
rect 119664 14218 119706 14454
rect 119942 14218 119984 14454
rect 119664 14134 119984 14218
rect 119664 13898 119706 14134
rect 119942 13898 119984 14134
rect 119664 13856 119984 13898
rect 517940 14454 518260 14496
rect 517940 14218 517982 14454
rect 518218 14218 518260 14454
rect 517940 14134 518260 14218
rect 517940 13898 517982 14134
rect 518218 13898 518260 14134
rect 517940 13856 518260 13898
rect 116531 12612 116597 12613
rect 116531 12548 116532 12612
rect 116596 12548 116597 12612
rect 116531 12547 116597 12548
rect 116163 6900 116229 6901
rect 116163 6836 116164 6900
rect 116228 6836 116229 6900
rect 116163 6835 116229 6836
rect 116166 1461 116226 6835
rect 116534 1869 116594 12547
rect 116715 10708 116781 10709
rect 116715 10644 116716 10708
rect 116780 10644 116781 10708
rect 116715 10643 116781 10644
rect 116531 1868 116597 1869
rect 116531 1804 116532 1868
rect 116596 1804 116597 1868
rect 116531 1803 116597 1804
rect 116718 1733 116778 10643
rect 117267 8804 117333 8805
rect 117267 8740 117268 8804
rect 117332 8740 117333 8804
rect 117267 8739 117333 8740
rect 116715 1732 116781 1733
rect 116715 1668 116716 1732
rect 116780 1668 116781 1732
rect 116715 1667 116781 1668
rect 117270 1597 117330 8739
rect 117267 1596 117333 1597
rect 117267 1532 117268 1596
rect 117332 1532 117333 1596
rect 117267 1531 117333 1532
rect 116163 1460 116229 1461
rect 116163 1396 116164 1460
rect 116228 1396 116229 1460
rect 116163 1395 116229 1396
<< via4 >>
rect 1706 144218 1942 144454
rect 1706 143898 1942 144134
rect 109998 144218 110234 144454
rect 109998 143898 110234 144134
rect 119706 144218 119942 144454
rect 119706 143898 119942 144134
rect 517982 144218 518218 144454
rect 517982 143898 518218 144134
rect 1096 131218 1332 131454
rect 1096 130898 1332 131134
rect 110658 131218 110894 131454
rect 110658 130898 110894 131134
rect 119046 131218 119282 131454
rect 119046 130898 119282 131134
rect 518642 131218 518878 131454
rect 518642 130898 518878 131134
rect 1706 118218 1942 118454
rect 1706 117898 1942 118134
rect 109998 118218 110234 118454
rect 109998 117898 110234 118134
rect 119706 118218 119942 118454
rect 119706 117898 119942 118134
rect 517982 118218 518218 118454
rect 517982 117898 518218 118134
rect 1096 105218 1332 105454
rect 1096 104898 1332 105134
rect 110658 105218 110894 105454
rect 110658 104898 110894 105134
rect 119046 105218 119282 105454
rect 119046 104898 119282 105134
rect 518642 105218 518878 105454
rect 518642 104898 518878 105134
rect 1706 92218 1942 92454
rect 1706 91898 1942 92134
rect 109998 92218 110234 92454
rect 109998 91898 110234 92134
rect 119706 92218 119942 92454
rect 119706 91898 119942 92134
rect 517982 92218 518218 92454
rect 517982 91898 518218 92134
rect 1096 79218 1332 79454
rect 1096 78898 1332 79134
rect 110658 79218 110894 79454
rect 110658 78898 110894 79134
rect 119046 79218 119282 79454
rect 119046 78898 119282 79134
rect 518642 79218 518878 79454
rect 518642 78898 518878 79134
rect 1706 66218 1942 66454
rect 1706 65898 1942 66134
rect 109998 66218 110234 66454
rect 109998 65898 110234 66134
rect 119706 66218 119942 66454
rect 119706 65898 119942 66134
rect 517982 66218 518218 66454
rect 517982 65898 518218 66134
rect 1096 53218 1332 53454
rect 1096 52898 1332 53134
rect 110658 53218 110894 53454
rect 110658 52898 110894 53134
rect 119046 53218 119282 53454
rect 119046 52898 119282 53134
rect 518642 53218 518878 53454
rect 518642 52898 518878 53134
rect 1706 40218 1942 40454
rect 1706 39898 1942 40134
rect 109998 40218 110234 40454
rect 109998 39898 110234 40134
rect 119706 40218 119942 40454
rect 119706 39898 119942 40134
rect 517982 40218 518218 40454
rect 517982 39898 518218 40134
rect 1096 27218 1332 27454
rect 1096 26898 1332 27134
rect 110658 27218 110894 27454
rect 110658 26898 110894 27134
rect 119046 27218 119282 27454
rect 119046 26898 119282 27134
rect 518642 27218 518878 27454
rect 518642 26898 518878 27134
rect 1706 14218 1942 14454
rect 1706 13898 1942 14134
rect 109998 14218 110234 14454
rect 109998 13898 110234 14134
rect 119706 14218 119942 14454
rect 119706 13898 119942 14134
rect 517982 14218 518218 14454
rect 517982 13898 518218 14134
<< metal5 >>
rect 1104 156856 522836 157496
rect 1104 144454 2200 144496
rect 1104 144218 1706 144454
rect 1942 144218 2200 144454
rect 1104 144134 2200 144218
rect 1104 143898 1706 144134
rect 1942 143898 2200 144134
rect 1104 143856 2200 143898
rect 109800 144454 120200 144496
rect 109800 144218 109998 144454
rect 110234 144218 119706 144454
rect 119942 144218 120200 144454
rect 109800 144134 120200 144218
rect 109800 143898 109998 144134
rect 110234 143898 119706 144134
rect 119942 143898 120200 144134
rect 109800 143856 120200 143898
rect 517800 144454 522836 144496
rect 517800 144218 517982 144454
rect 518218 144218 522836 144454
rect 517800 144134 522836 144218
rect 517800 143898 517982 144134
rect 518218 143898 522836 144134
rect 517800 143856 522836 143898
rect 1072 131454 2200 131496
rect 1072 131218 1096 131454
rect 1332 131218 2200 131454
rect 1072 131134 2200 131218
rect 1072 130898 1096 131134
rect 1332 130898 2200 131134
rect 1072 130856 2200 130898
rect 109800 131454 120200 131496
rect 109800 131218 110658 131454
rect 110894 131218 119046 131454
rect 119282 131218 120200 131454
rect 109800 131134 120200 131218
rect 109800 130898 110658 131134
rect 110894 130898 119046 131134
rect 119282 130898 120200 131134
rect 109800 130856 120200 130898
rect 517800 131454 522836 131496
rect 517800 131218 518642 131454
rect 518878 131218 522836 131454
rect 517800 131134 522836 131218
rect 517800 130898 518642 131134
rect 518878 130898 522836 131134
rect 517800 130856 522836 130898
rect 1104 118454 2200 118496
rect 1104 118218 1706 118454
rect 1942 118218 2200 118454
rect 1104 118134 2200 118218
rect 1104 117898 1706 118134
rect 1942 117898 2200 118134
rect 1104 117856 2200 117898
rect 109800 118454 120200 118496
rect 109800 118218 109998 118454
rect 110234 118218 119706 118454
rect 119942 118218 120200 118454
rect 109800 118134 120200 118218
rect 109800 117898 109998 118134
rect 110234 117898 119706 118134
rect 119942 117898 120200 118134
rect 109800 117856 120200 117898
rect 517800 118454 522836 118496
rect 517800 118218 517982 118454
rect 518218 118218 522836 118454
rect 517800 118134 522836 118218
rect 517800 117898 517982 118134
rect 518218 117898 522836 118134
rect 517800 117856 522836 117898
rect 1072 105454 2200 105496
rect 1072 105218 1096 105454
rect 1332 105218 2200 105454
rect 1072 105134 2200 105218
rect 1072 104898 1096 105134
rect 1332 104898 2200 105134
rect 1072 104856 2200 104898
rect 109800 105454 120200 105496
rect 109800 105218 110658 105454
rect 110894 105218 119046 105454
rect 119282 105218 120200 105454
rect 109800 105134 120200 105218
rect 109800 104898 110658 105134
rect 110894 104898 119046 105134
rect 119282 104898 120200 105134
rect 109800 104856 120200 104898
rect 517800 105454 522836 105496
rect 517800 105218 518642 105454
rect 518878 105218 522836 105454
rect 517800 105134 522836 105218
rect 517800 104898 518642 105134
rect 518878 104898 522836 105134
rect 517800 104856 522836 104898
rect 1104 92454 2200 92496
rect 1104 92218 1706 92454
rect 1942 92218 2200 92454
rect 1104 92134 2200 92218
rect 1104 91898 1706 92134
rect 1942 91898 2200 92134
rect 1104 91856 2200 91898
rect 109800 92454 120200 92496
rect 109800 92218 109998 92454
rect 110234 92218 119706 92454
rect 119942 92218 120200 92454
rect 109800 92134 120200 92218
rect 109800 91898 109998 92134
rect 110234 91898 119706 92134
rect 119942 91898 120200 92134
rect 109800 91856 120200 91898
rect 517800 92454 522836 92496
rect 517800 92218 517982 92454
rect 518218 92218 522836 92454
rect 517800 92134 522836 92218
rect 517800 91898 517982 92134
rect 518218 91898 522836 92134
rect 517800 91856 522836 91898
rect 1072 79454 2200 79496
rect 1072 79218 1096 79454
rect 1332 79218 2200 79454
rect 1072 79134 2200 79218
rect 1072 78898 1096 79134
rect 1332 78898 2200 79134
rect 1072 78856 2200 78898
rect 109800 79454 120200 79496
rect 109800 79218 110658 79454
rect 110894 79218 119046 79454
rect 119282 79218 120200 79454
rect 109800 79134 120200 79218
rect 109800 78898 110658 79134
rect 110894 78898 119046 79134
rect 119282 78898 120200 79134
rect 109800 78856 120200 78898
rect 517800 79454 522836 79496
rect 517800 79218 518642 79454
rect 518878 79218 522836 79454
rect 517800 79134 522836 79218
rect 517800 78898 518642 79134
rect 518878 78898 522836 79134
rect 517800 78856 522836 78898
rect 1104 66454 2200 66496
rect 1104 66218 1706 66454
rect 1942 66218 2200 66454
rect 1104 66134 2200 66218
rect 1104 65898 1706 66134
rect 1942 65898 2200 66134
rect 1104 65856 2200 65898
rect 109800 66454 120200 66496
rect 109800 66218 109998 66454
rect 110234 66218 119706 66454
rect 119942 66218 120200 66454
rect 109800 66134 120200 66218
rect 109800 65898 109998 66134
rect 110234 65898 119706 66134
rect 119942 65898 120200 66134
rect 109800 65856 120200 65898
rect 517800 66454 522836 66496
rect 517800 66218 517982 66454
rect 518218 66218 522836 66454
rect 517800 66134 522836 66218
rect 517800 65898 517982 66134
rect 518218 65898 522836 66134
rect 517800 65856 522836 65898
rect 1072 53454 2200 53496
rect 1072 53218 1096 53454
rect 1332 53218 2200 53454
rect 1072 53134 2200 53218
rect 1072 52898 1096 53134
rect 1332 52898 2200 53134
rect 1072 52856 2200 52898
rect 109800 53454 120200 53496
rect 109800 53218 110658 53454
rect 110894 53218 119046 53454
rect 119282 53218 120200 53454
rect 109800 53134 120200 53218
rect 109800 52898 110658 53134
rect 110894 52898 119046 53134
rect 119282 52898 120200 53134
rect 109800 52856 120200 52898
rect 517800 53454 522836 53496
rect 517800 53218 518642 53454
rect 518878 53218 522836 53454
rect 517800 53134 522836 53218
rect 517800 52898 518642 53134
rect 518878 52898 522836 53134
rect 517800 52856 522836 52898
rect 1104 40454 2200 40496
rect 1104 40218 1706 40454
rect 1942 40218 2200 40454
rect 1104 40134 2200 40218
rect 1104 39898 1706 40134
rect 1942 39898 2200 40134
rect 1104 39856 2200 39898
rect 109800 40454 120200 40496
rect 109800 40218 109998 40454
rect 110234 40218 119706 40454
rect 119942 40218 120200 40454
rect 109800 40134 120200 40218
rect 109800 39898 109998 40134
rect 110234 39898 119706 40134
rect 119942 39898 120200 40134
rect 109800 39856 120200 39898
rect 517800 40454 522836 40496
rect 517800 40218 517982 40454
rect 518218 40218 522836 40454
rect 517800 40134 522836 40218
rect 517800 39898 517982 40134
rect 518218 39898 522836 40134
rect 517800 39856 522836 39898
rect 1072 27454 2200 27496
rect 1072 27218 1096 27454
rect 1332 27218 2200 27454
rect 1072 27134 2200 27218
rect 1072 26898 1096 27134
rect 1332 26898 2200 27134
rect 1072 26856 2200 26898
rect 109800 27454 120200 27496
rect 109800 27218 110658 27454
rect 110894 27218 119046 27454
rect 119282 27218 120200 27454
rect 109800 27134 120200 27218
rect 109800 26898 110658 27134
rect 110894 26898 119046 27134
rect 119282 26898 120200 27134
rect 109800 26856 120200 26898
rect 517800 27454 522836 27496
rect 517800 27218 518642 27454
rect 518878 27218 522836 27454
rect 517800 27134 522836 27218
rect 517800 26898 518642 27134
rect 518878 26898 522836 27134
rect 517800 26856 522836 26898
rect 1104 14454 2200 14496
rect 1104 14218 1706 14454
rect 1942 14218 2200 14454
rect 1104 14134 2200 14218
rect 1104 13898 1706 14134
rect 1942 13898 2200 14134
rect 1104 13856 2200 13898
rect 109800 14454 120200 14496
rect 109800 14218 109998 14454
rect 110234 14218 119706 14454
rect 119942 14218 120200 14454
rect 109800 14134 120200 14218
rect 109800 13898 109998 14134
rect 110234 13898 119706 14134
rect 119942 13898 120200 14134
rect 109800 13856 120200 13898
rect 517800 14454 522836 14496
rect 517800 14218 517982 14454
rect 518218 14218 522836 14454
rect 517800 14134 522836 14218
rect 517800 13898 517982 14134
rect 518218 13898 522836 14134
rect 517800 13856 522836 13898
use mgmt_core  core
timestamp 1648060287
transform 1 0 119000 0 1 2000
box 0 0 400000 148000
use DFFRAM  DFFRAM_0
timestamp 1648060287
transform 1 0 1000 0 1 2000
box 4 0 110000 148000
<< labels >>
rlabel metal5 s 1104 26856 2200 27496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 26856 120200 27496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 26856 522836 27496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 52856 2200 53496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 52856 120200 53496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 52856 522836 53496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 78856 2200 79496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 78856 120200 79496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 78856 522836 79496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 104856 2200 105496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 104856 120200 105496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 104856 522836 105496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 130856 2200 131496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 130856 120200 131496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 130856 522836 131496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 156856 522836 157496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 13856 2200 14496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 13856 120200 14496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 13856 522836 14496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 39856 2200 40496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 39856 120200 40496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 39856 522836 40496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 65856 2200 66496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 65856 120200 66496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 65856 522836 66496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 91856 2200 92496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 91856 120200 92496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 91856 522836 92496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 117856 2200 118496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 117856 120200 118496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 117856 522836 118496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 143856 2200 144496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 143856 120200 144496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 143856 522836 144496 6 VPWR
port 1 nsew power input
rlabel metal2 s 294786 -400 294842 800 6 core_clk
port 2 nsew signal input
rlabel metal2 s 98274 -400 98330 800 6 core_rstn
port 3 nsew signal input
rlabel metal3 s 523200 63792 524400 63912 6 debug_in
port 4 nsew signal input
rlabel metal3 s 523200 65288 524400 65408 6 debug_mode
port 5 nsew signal tristate
rlabel metal3 s 523200 66784 524400 66904 6 debug_oeb
port 6 nsew signal tristate
rlabel metal3 s 523200 68280 524400 68400 6 debug_out
port 7 nsew signal tristate
rlabel metal3 s 523200 145120 524400 145240 6 flash_clk
port 8 nsew signal tristate
rlabel metal3 s 523200 143624 524400 143744 6 flash_csb
port 9 nsew signal tristate
rlabel metal3 s 523200 146616 524400 146736 6 flash_io0_di
port 10 nsew signal input
rlabel metal3 s 523200 148112 524400 148232 6 flash_io0_do
port 11 nsew signal tristate
rlabel metal3 s 523200 149608 524400 149728 6 flash_io0_oeb
port 12 nsew signal tristate
rlabel metal3 s 523200 151104 524400 151224 6 flash_io1_di
port 13 nsew signal input
rlabel metal3 s 523200 152600 524400 152720 6 flash_io1_do
port 14 nsew signal tristate
rlabel metal3 s 523200 154096 524400 154216 6 flash_io1_oeb
port 15 nsew signal tristate
rlabel metal3 s 523200 155592 524400 155712 6 flash_io2_di
port 16 nsew signal input
rlabel metal3 s 523200 157088 524400 157208 6 flash_io2_do
port 17 nsew signal tristate
rlabel metal3 s 523200 158584 524400 158704 6 flash_io2_oeb
port 18 nsew signal tristate
rlabel metal3 s 523200 160080 524400 160200 6 flash_io3_di
port 19 nsew signal input
rlabel metal3 s 523200 161576 524400 161696 6 flash_io3_do
port 20 nsew signal tristate
rlabel metal3 s 523200 163072 524400 163192 6 flash_io3_oeb
port 21 nsew signal tristate
rlabel metal2 s 32770 -400 32826 800 6 gpio_in_pad
port 22 nsew signal input
rlabel metal2 s 163778 -400 163834 800 6 gpio_inenb_pad
port 23 nsew signal tristate
rlabel metal2 s 229282 -400 229338 800 6 gpio_mode0_pad
port 24 nsew signal tristate
rlabel metal2 s 360290 -400 360346 800 6 gpio_mode1_pad
port 25 nsew signal tristate
rlabel metal2 s 425794 -400 425850 800 6 gpio_out_pad
port 26 nsew signal tristate
rlabel metal2 s 491298 -400 491354 800 6 gpio_outenb_pad
port 27 nsew signal tristate
rlabel metal3 s 523200 90856 524400 90976 6 hk_ack_i
port 28 nsew signal input
rlabel metal3 s 523200 93848 524400 93968 6 hk_cyc_o
port 29 nsew signal tristate
rlabel metal3 s 523200 95480 524400 95600 6 hk_dat_i[0]
port 30 nsew signal input
rlabel metal3 s 523200 110440 524400 110560 6 hk_dat_i[10]
port 31 nsew signal input
rlabel metal3 s 523200 111936 524400 112056 6 hk_dat_i[11]
port 32 nsew signal input
rlabel metal3 s 523200 113432 524400 113552 6 hk_dat_i[12]
port 33 nsew signal input
rlabel metal3 s 523200 114928 524400 115048 6 hk_dat_i[13]
port 34 nsew signal input
rlabel metal3 s 523200 116424 524400 116544 6 hk_dat_i[14]
port 35 nsew signal input
rlabel metal3 s 523200 118056 524400 118176 6 hk_dat_i[15]
port 36 nsew signal input
rlabel metal3 s 523200 119552 524400 119672 6 hk_dat_i[16]
port 37 nsew signal input
rlabel metal3 s 523200 121048 524400 121168 6 hk_dat_i[17]
port 38 nsew signal input
rlabel metal3 s 523200 122544 524400 122664 6 hk_dat_i[18]
port 39 nsew signal input
rlabel metal3 s 523200 124040 524400 124160 6 hk_dat_i[19]
port 40 nsew signal input
rlabel metal3 s 523200 96976 524400 97096 6 hk_dat_i[1]
port 41 nsew signal input
rlabel metal3 s 523200 125536 524400 125656 6 hk_dat_i[20]
port 42 nsew signal input
rlabel metal3 s 523200 127032 524400 127152 6 hk_dat_i[21]
port 43 nsew signal input
rlabel metal3 s 523200 128528 524400 128648 6 hk_dat_i[22]
port 44 nsew signal input
rlabel metal3 s 523200 130024 524400 130144 6 hk_dat_i[23]
port 45 nsew signal input
rlabel metal3 s 523200 131520 524400 131640 6 hk_dat_i[24]
port 46 nsew signal input
rlabel metal3 s 523200 133016 524400 133136 6 hk_dat_i[25]
port 47 nsew signal input
rlabel metal3 s 523200 134512 524400 134632 6 hk_dat_i[26]
port 48 nsew signal input
rlabel metal3 s 523200 136008 524400 136128 6 hk_dat_i[27]
port 49 nsew signal input
rlabel metal3 s 523200 137504 524400 137624 6 hk_dat_i[28]
port 50 nsew signal input
rlabel metal3 s 523200 139000 524400 139120 6 hk_dat_i[29]
port 51 nsew signal input
rlabel metal3 s 523200 98472 524400 98592 6 hk_dat_i[2]
port 52 nsew signal input
rlabel metal3 s 523200 140496 524400 140616 6 hk_dat_i[30]
port 53 nsew signal input
rlabel metal3 s 523200 142128 524400 142248 6 hk_dat_i[31]
port 54 nsew signal input
rlabel metal3 s 523200 99968 524400 100088 6 hk_dat_i[3]
port 55 nsew signal input
rlabel metal3 s 523200 101464 524400 101584 6 hk_dat_i[4]
port 56 nsew signal input
rlabel metal3 s 523200 102960 524400 103080 6 hk_dat_i[5]
port 57 nsew signal input
rlabel metal3 s 523200 104456 524400 104576 6 hk_dat_i[6]
port 58 nsew signal input
rlabel metal3 s 523200 105952 524400 106072 6 hk_dat_i[7]
port 59 nsew signal input
rlabel metal3 s 523200 107448 524400 107568 6 hk_dat_i[8]
port 60 nsew signal input
rlabel metal3 s 523200 108944 524400 109064 6 hk_dat_i[9]
port 61 nsew signal input
rlabel metal3 s 523200 92352 524400 92472 6 hk_stb_o
port 62 nsew signal tristate
rlabel metal2 s 521842 163200 521898 164400 6 irq[0]
port 63 nsew signal input
rlabel metal2 s 522670 163200 522726 164400 6 irq[1]
port 64 nsew signal input
rlabel metal2 s 523498 163200 523554 164400 6 irq[2]
port 65 nsew signal input
rlabel metal3 s 523200 74400 524400 74520 6 irq[3]
port 66 nsew signal input
rlabel metal3 s 523200 72904 524400 73024 6 irq[4]
port 67 nsew signal input
rlabel metal3 s 523200 71408 524400 71528 6 irq[5]
port 68 nsew signal input
rlabel metal2 s 386 163200 442 164400 6 la_iena[0]
port 69 nsew signal tristate
rlabel metal2 s 336830 163200 336886 164400 6 la_iena[100]
port 70 nsew signal tristate
rlabel metal2 s 340142 163200 340198 164400 6 la_iena[101]
port 71 nsew signal tristate
rlabel metal2 s 343546 163200 343602 164400 6 la_iena[102]
port 72 nsew signal tristate
rlabel metal2 s 346858 163200 346914 164400 6 la_iena[103]
port 73 nsew signal tristate
rlabel metal2 s 350262 163200 350318 164400 6 la_iena[104]
port 74 nsew signal tristate
rlabel metal2 s 353666 163200 353722 164400 6 la_iena[105]
port 75 nsew signal tristate
rlabel metal2 s 356978 163200 357034 164400 6 la_iena[106]
port 76 nsew signal tristate
rlabel metal2 s 360382 163200 360438 164400 6 la_iena[107]
port 77 nsew signal tristate
rlabel metal2 s 363694 163200 363750 164400 6 la_iena[108]
port 78 nsew signal tristate
rlabel metal2 s 367098 163200 367154 164400 6 la_iena[109]
port 79 nsew signal tristate
rlabel metal2 s 33966 163200 34022 164400 6 la_iena[10]
port 80 nsew signal tristate
rlabel metal2 s 370410 163200 370466 164400 6 la_iena[110]
port 81 nsew signal tristate
rlabel metal2 s 373814 163200 373870 164400 6 la_iena[111]
port 82 nsew signal tristate
rlabel metal2 s 377218 163200 377274 164400 6 la_iena[112]
port 83 nsew signal tristate
rlabel metal2 s 380530 163200 380586 164400 6 la_iena[113]
port 84 nsew signal tristate
rlabel metal2 s 383934 163200 383990 164400 6 la_iena[114]
port 85 nsew signal tristate
rlabel metal2 s 387246 163200 387302 164400 6 la_iena[115]
port 86 nsew signal tristate
rlabel metal2 s 390650 163200 390706 164400 6 la_iena[116]
port 87 nsew signal tristate
rlabel metal2 s 393962 163200 394018 164400 6 la_iena[117]
port 88 nsew signal tristate
rlabel metal2 s 397366 163200 397422 164400 6 la_iena[118]
port 89 nsew signal tristate
rlabel metal2 s 400770 163200 400826 164400 6 la_iena[119]
port 90 nsew signal tristate
rlabel metal2 s 37370 163200 37426 164400 6 la_iena[11]
port 91 nsew signal tristate
rlabel metal2 s 404082 163200 404138 164400 6 la_iena[120]
port 92 nsew signal tristate
rlabel metal2 s 407486 163200 407542 164400 6 la_iena[121]
port 93 nsew signal tristate
rlabel metal2 s 410798 163200 410854 164400 6 la_iena[122]
port 94 nsew signal tristate
rlabel metal2 s 414202 163200 414258 164400 6 la_iena[123]
port 95 nsew signal tristate
rlabel metal2 s 417514 163200 417570 164400 6 la_iena[124]
port 96 nsew signal tristate
rlabel metal2 s 420918 163200 420974 164400 6 la_iena[125]
port 97 nsew signal tristate
rlabel metal2 s 424322 163200 424378 164400 6 la_iena[126]
port 98 nsew signal tristate
rlabel metal2 s 427634 163200 427690 164400 6 la_iena[127]
port 99 nsew signal tristate
rlabel metal2 s 40682 163200 40738 164400 6 la_iena[12]
port 100 nsew signal tristate
rlabel metal2 s 44086 163200 44142 164400 6 la_iena[13]
port 101 nsew signal tristate
rlabel metal2 s 47490 163200 47546 164400 6 la_iena[14]
port 102 nsew signal tristate
rlabel metal2 s 50802 163200 50858 164400 6 la_iena[15]
port 103 nsew signal tristate
rlabel metal2 s 54206 163200 54262 164400 6 la_iena[16]
port 104 nsew signal tristate
rlabel metal2 s 57518 163200 57574 164400 6 la_iena[17]
port 105 nsew signal tristate
rlabel metal2 s 60922 163200 60978 164400 6 la_iena[18]
port 106 nsew signal tristate
rlabel metal2 s 64234 163200 64290 164400 6 la_iena[19]
port 107 nsew signal tristate
rlabel metal2 s 3698 163200 3754 164400 6 la_iena[1]
port 108 nsew signal tristate
rlabel metal2 s 67638 163200 67694 164400 6 la_iena[20]
port 109 nsew signal tristate
rlabel metal2 s 71042 163200 71098 164400 6 la_iena[21]
port 110 nsew signal tristate
rlabel metal2 s 74354 163200 74410 164400 6 la_iena[22]
port 111 nsew signal tristate
rlabel metal2 s 77758 163200 77814 164400 6 la_iena[23]
port 112 nsew signal tristate
rlabel metal2 s 81070 163200 81126 164400 6 la_iena[24]
port 113 nsew signal tristate
rlabel metal2 s 84474 163200 84530 164400 6 la_iena[25]
port 114 nsew signal tristate
rlabel metal2 s 87786 163200 87842 164400 6 la_iena[26]
port 115 nsew signal tristate
rlabel metal2 s 91190 163200 91246 164400 6 la_iena[27]
port 116 nsew signal tristate
rlabel metal2 s 94594 163200 94650 164400 6 la_iena[28]
port 117 nsew signal tristate
rlabel metal2 s 97906 163200 97962 164400 6 la_iena[29]
port 118 nsew signal tristate
rlabel metal2 s 7102 163200 7158 164400 6 la_iena[2]
port 119 nsew signal tristate
rlabel metal2 s 101310 163200 101366 164400 6 la_iena[30]
port 120 nsew signal tristate
rlabel metal2 s 104622 163200 104678 164400 6 la_iena[31]
port 121 nsew signal tristate
rlabel metal2 s 108026 163200 108082 164400 6 la_iena[32]
port 122 nsew signal tristate
rlabel metal2 s 111338 163200 111394 164400 6 la_iena[33]
port 123 nsew signal tristate
rlabel metal2 s 114742 163200 114798 164400 6 la_iena[34]
port 124 nsew signal tristate
rlabel metal2 s 118146 163200 118202 164400 6 la_iena[35]
port 125 nsew signal tristate
rlabel metal2 s 121458 163200 121514 164400 6 la_iena[36]
port 126 nsew signal tristate
rlabel metal2 s 124862 163200 124918 164400 6 la_iena[37]
port 127 nsew signal tristate
rlabel metal2 s 128174 163200 128230 164400 6 la_iena[38]
port 128 nsew signal tristate
rlabel metal2 s 131578 163200 131634 164400 6 la_iena[39]
port 129 nsew signal tristate
rlabel metal2 s 10414 163200 10470 164400 6 la_iena[3]
port 130 nsew signal tristate
rlabel metal2 s 134890 163200 134946 164400 6 la_iena[40]
port 131 nsew signal tristate
rlabel metal2 s 138294 163200 138350 164400 6 la_iena[41]
port 132 nsew signal tristate
rlabel metal2 s 141698 163200 141754 164400 6 la_iena[42]
port 133 nsew signal tristate
rlabel metal2 s 145010 163200 145066 164400 6 la_iena[43]
port 134 nsew signal tristate
rlabel metal2 s 148414 163200 148470 164400 6 la_iena[44]
port 135 nsew signal tristate
rlabel metal2 s 151726 163200 151782 164400 6 la_iena[45]
port 136 nsew signal tristate
rlabel metal2 s 155130 163200 155186 164400 6 la_iena[46]
port 137 nsew signal tristate
rlabel metal2 s 158442 163200 158498 164400 6 la_iena[47]
port 138 nsew signal tristate
rlabel metal2 s 161846 163200 161902 164400 6 la_iena[48]
port 139 nsew signal tristate
rlabel metal2 s 165250 163200 165306 164400 6 la_iena[49]
port 140 nsew signal tristate
rlabel metal2 s 13818 163200 13874 164400 6 la_iena[4]
port 141 nsew signal tristate
rlabel metal2 s 168562 163200 168618 164400 6 la_iena[50]
port 142 nsew signal tristate
rlabel metal2 s 171966 163200 172022 164400 6 la_iena[51]
port 143 nsew signal tristate
rlabel metal2 s 175278 163200 175334 164400 6 la_iena[52]
port 144 nsew signal tristate
rlabel metal2 s 178682 163200 178738 164400 6 la_iena[53]
port 145 nsew signal tristate
rlabel metal2 s 181994 163200 182050 164400 6 la_iena[54]
port 146 nsew signal tristate
rlabel metal2 s 185398 163200 185454 164400 6 la_iena[55]
port 147 nsew signal tristate
rlabel metal2 s 188802 163200 188858 164400 6 la_iena[56]
port 148 nsew signal tristate
rlabel metal2 s 192114 163200 192170 164400 6 la_iena[57]
port 149 nsew signal tristate
rlabel metal2 s 195518 163200 195574 164400 6 la_iena[58]
port 150 nsew signal tristate
rlabel metal2 s 198830 163200 198886 164400 6 la_iena[59]
port 151 nsew signal tristate
rlabel metal2 s 17130 163200 17186 164400 6 la_iena[5]
port 152 nsew signal tristate
rlabel metal2 s 202234 163200 202290 164400 6 la_iena[60]
port 153 nsew signal tristate
rlabel metal2 s 205546 163200 205602 164400 6 la_iena[61]
port 154 nsew signal tristate
rlabel metal2 s 208950 163200 209006 164400 6 la_iena[62]
port 155 nsew signal tristate
rlabel metal2 s 212354 163200 212410 164400 6 la_iena[63]
port 156 nsew signal tristate
rlabel metal2 s 215666 163200 215722 164400 6 la_iena[64]
port 157 nsew signal tristate
rlabel metal2 s 219070 163200 219126 164400 6 la_iena[65]
port 158 nsew signal tristate
rlabel metal2 s 222382 163200 222438 164400 6 la_iena[66]
port 159 nsew signal tristate
rlabel metal2 s 225786 163200 225842 164400 6 la_iena[67]
port 160 nsew signal tristate
rlabel metal2 s 229098 163200 229154 164400 6 la_iena[68]
port 161 nsew signal tristate
rlabel metal2 s 232502 163200 232558 164400 6 la_iena[69]
port 162 nsew signal tristate
rlabel metal2 s 20534 163200 20590 164400 6 la_iena[6]
port 163 nsew signal tristate
rlabel metal2 s 235906 163200 235962 164400 6 la_iena[70]
port 164 nsew signal tristate
rlabel metal2 s 239218 163200 239274 164400 6 la_iena[71]
port 165 nsew signal tristate
rlabel metal2 s 242622 163200 242678 164400 6 la_iena[72]
port 166 nsew signal tristate
rlabel metal2 s 245934 163200 245990 164400 6 la_iena[73]
port 167 nsew signal tristate
rlabel metal2 s 249338 163200 249394 164400 6 la_iena[74]
port 168 nsew signal tristate
rlabel metal2 s 252650 163200 252706 164400 6 la_iena[75]
port 169 nsew signal tristate
rlabel metal2 s 256054 163200 256110 164400 6 la_iena[76]
port 170 nsew signal tristate
rlabel metal2 s 259458 163200 259514 164400 6 la_iena[77]
port 171 nsew signal tristate
rlabel metal2 s 262770 163200 262826 164400 6 la_iena[78]
port 172 nsew signal tristate
rlabel metal2 s 266174 163200 266230 164400 6 la_iena[79]
port 173 nsew signal tristate
rlabel metal2 s 23938 163200 23994 164400 6 la_iena[7]
port 174 nsew signal tristate
rlabel metal2 s 269486 163200 269542 164400 6 la_iena[80]
port 175 nsew signal tristate
rlabel metal2 s 272890 163200 272946 164400 6 la_iena[81]
port 176 nsew signal tristate
rlabel metal2 s 276202 163200 276258 164400 6 la_iena[82]
port 177 nsew signal tristate
rlabel metal2 s 279606 163200 279662 164400 6 la_iena[83]
port 178 nsew signal tristate
rlabel metal2 s 283010 163200 283066 164400 6 la_iena[84]
port 179 nsew signal tristate
rlabel metal2 s 286322 163200 286378 164400 6 la_iena[85]
port 180 nsew signal tristate
rlabel metal2 s 289726 163200 289782 164400 6 la_iena[86]
port 181 nsew signal tristate
rlabel metal2 s 293038 163200 293094 164400 6 la_iena[87]
port 182 nsew signal tristate
rlabel metal2 s 296442 163200 296498 164400 6 la_iena[88]
port 183 nsew signal tristate
rlabel metal2 s 299754 163200 299810 164400 6 la_iena[89]
port 184 nsew signal tristate
rlabel metal2 s 27250 163200 27306 164400 6 la_iena[8]
port 185 nsew signal tristate
rlabel metal2 s 303158 163200 303214 164400 6 la_iena[90]
port 186 nsew signal tristate
rlabel metal2 s 306562 163200 306618 164400 6 la_iena[91]
port 187 nsew signal tristate
rlabel metal2 s 309874 163200 309930 164400 6 la_iena[92]
port 188 nsew signal tristate
rlabel metal2 s 313278 163200 313334 164400 6 la_iena[93]
port 189 nsew signal tristate
rlabel metal2 s 316590 163200 316646 164400 6 la_iena[94]
port 190 nsew signal tristate
rlabel metal2 s 319994 163200 320050 164400 6 la_iena[95]
port 191 nsew signal tristate
rlabel metal2 s 323306 163200 323362 164400 6 la_iena[96]
port 192 nsew signal tristate
rlabel metal2 s 326710 163200 326766 164400 6 la_iena[97]
port 193 nsew signal tristate
rlabel metal2 s 330114 163200 330170 164400 6 la_iena[98]
port 194 nsew signal tristate
rlabel metal2 s 333426 163200 333482 164400 6 la_iena[99]
port 195 nsew signal tristate
rlabel metal2 s 30654 163200 30710 164400 6 la_iena[9]
port 196 nsew signal tristate
rlabel metal2 s 1214 163200 1270 164400 6 la_input[0]
port 197 nsew signal input
rlabel metal2 s 337658 163200 337714 164400 6 la_input[100]
port 198 nsew signal input
rlabel metal2 s 340970 163200 341026 164400 6 la_input[101]
port 199 nsew signal input
rlabel metal2 s 344374 163200 344430 164400 6 la_input[102]
port 200 nsew signal input
rlabel metal2 s 347778 163200 347834 164400 6 la_input[103]
port 201 nsew signal input
rlabel metal2 s 351090 163200 351146 164400 6 la_input[104]
port 202 nsew signal input
rlabel metal2 s 354494 163200 354550 164400 6 la_input[105]
port 203 nsew signal input
rlabel metal2 s 357806 163200 357862 164400 6 la_input[106]
port 204 nsew signal input
rlabel metal2 s 361210 163200 361266 164400 6 la_input[107]
port 205 nsew signal input
rlabel metal2 s 364522 163200 364578 164400 6 la_input[108]
port 206 nsew signal input
rlabel metal2 s 367926 163200 367982 164400 6 la_input[109]
port 207 nsew signal input
rlabel metal2 s 34794 163200 34850 164400 6 la_input[10]
port 208 nsew signal input
rlabel metal2 s 371330 163200 371386 164400 6 la_input[110]
port 209 nsew signal input
rlabel metal2 s 374642 163200 374698 164400 6 la_input[111]
port 210 nsew signal input
rlabel metal2 s 378046 163200 378102 164400 6 la_input[112]
port 211 nsew signal input
rlabel metal2 s 381358 163200 381414 164400 6 la_input[113]
port 212 nsew signal input
rlabel metal2 s 384762 163200 384818 164400 6 la_input[114]
port 213 nsew signal input
rlabel metal2 s 388074 163200 388130 164400 6 la_input[115]
port 214 nsew signal input
rlabel metal2 s 391478 163200 391534 164400 6 la_input[116]
port 215 nsew signal input
rlabel metal2 s 394882 163200 394938 164400 6 la_input[117]
port 216 nsew signal input
rlabel metal2 s 398194 163200 398250 164400 6 la_input[118]
port 217 nsew signal input
rlabel metal2 s 401598 163200 401654 164400 6 la_input[119]
port 218 nsew signal input
rlabel metal2 s 38198 163200 38254 164400 6 la_input[11]
port 219 nsew signal input
rlabel metal2 s 404910 163200 404966 164400 6 la_input[120]
port 220 nsew signal input
rlabel metal2 s 408314 163200 408370 164400 6 la_input[121]
port 221 nsew signal input
rlabel metal2 s 411626 163200 411682 164400 6 la_input[122]
port 222 nsew signal input
rlabel metal2 s 415030 163200 415086 164400 6 la_input[123]
port 223 nsew signal input
rlabel metal2 s 418434 163200 418490 164400 6 la_input[124]
port 224 nsew signal input
rlabel metal2 s 421746 163200 421802 164400 6 la_input[125]
port 225 nsew signal input
rlabel metal2 s 425150 163200 425206 164400 6 la_input[126]
port 226 nsew signal input
rlabel metal2 s 428462 163200 428518 164400 6 la_input[127]
port 227 nsew signal input
rlabel metal2 s 41602 163200 41658 164400 6 la_input[12]
port 228 nsew signal input
rlabel metal2 s 44914 163200 44970 164400 6 la_input[13]
port 229 nsew signal input
rlabel metal2 s 48318 163200 48374 164400 6 la_input[14]
port 230 nsew signal input
rlabel metal2 s 51630 163200 51686 164400 6 la_input[15]
port 231 nsew signal input
rlabel metal2 s 55034 163200 55090 164400 6 la_input[16]
port 232 nsew signal input
rlabel metal2 s 58346 163200 58402 164400 6 la_input[17]
port 233 nsew signal input
rlabel metal2 s 61750 163200 61806 164400 6 la_input[18]
port 234 nsew signal input
rlabel metal2 s 65154 163200 65210 164400 6 la_input[19]
port 235 nsew signal input
rlabel metal2 s 4526 163200 4582 164400 6 la_input[1]
port 236 nsew signal input
rlabel metal2 s 68466 163200 68522 164400 6 la_input[20]
port 237 nsew signal input
rlabel metal2 s 71870 163200 71926 164400 6 la_input[21]
port 238 nsew signal input
rlabel metal2 s 75182 163200 75238 164400 6 la_input[22]
port 239 nsew signal input
rlabel metal2 s 78586 163200 78642 164400 6 la_input[23]
port 240 nsew signal input
rlabel metal2 s 81898 163200 81954 164400 6 la_input[24]
port 241 nsew signal input
rlabel metal2 s 85302 163200 85358 164400 6 la_input[25]
port 242 nsew signal input
rlabel metal2 s 88706 163200 88762 164400 6 la_input[26]
port 243 nsew signal input
rlabel metal2 s 92018 163200 92074 164400 6 la_input[27]
port 244 nsew signal input
rlabel metal2 s 95422 163200 95478 164400 6 la_input[28]
port 245 nsew signal input
rlabel metal2 s 98734 163200 98790 164400 6 la_input[29]
port 246 nsew signal input
rlabel metal2 s 7930 163200 7986 164400 6 la_input[2]
port 247 nsew signal input
rlabel metal2 s 102138 163200 102194 164400 6 la_input[30]
port 248 nsew signal input
rlabel metal2 s 105450 163200 105506 164400 6 la_input[31]
port 249 nsew signal input
rlabel metal2 s 108854 163200 108910 164400 6 la_input[32]
port 250 nsew signal input
rlabel metal2 s 112258 163200 112314 164400 6 la_input[33]
port 251 nsew signal input
rlabel metal2 s 115570 163200 115626 164400 6 la_input[34]
port 252 nsew signal input
rlabel metal2 s 118974 163200 119030 164400 6 la_input[35]
port 253 nsew signal input
rlabel metal2 s 122286 163200 122342 164400 6 la_input[36]
port 254 nsew signal input
rlabel metal2 s 125690 163200 125746 164400 6 la_input[37]
port 255 nsew signal input
rlabel metal2 s 129002 163200 129058 164400 6 la_input[38]
port 256 nsew signal input
rlabel metal2 s 132406 163200 132462 164400 6 la_input[39]
port 257 nsew signal input
rlabel metal2 s 11242 163200 11298 164400 6 la_input[3]
port 258 nsew signal input
rlabel metal2 s 135810 163200 135866 164400 6 la_input[40]
port 259 nsew signal input
rlabel metal2 s 139122 163200 139178 164400 6 la_input[41]
port 260 nsew signal input
rlabel metal2 s 142526 163200 142582 164400 6 la_input[42]
port 261 nsew signal input
rlabel metal2 s 145838 163200 145894 164400 6 la_input[43]
port 262 nsew signal input
rlabel metal2 s 149242 163200 149298 164400 6 la_input[44]
port 263 nsew signal input
rlabel metal2 s 152554 163200 152610 164400 6 la_input[45]
port 264 nsew signal input
rlabel metal2 s 155958 163200 156014 164400 6 la_input[46]
port 265 nsew signal input
rlabel metal2 s 159362 163200 159418 164400 6 la_input[47]
port 266 nsew signal input
rlabel metal2 s 162674 163200 162730 164400 6 la_input[48]
port 267 nsew signal input
rlabel metal2 s 166078 163200 166134 164400 6 la_input[49]
port 268 nsew signal input
rlabel metal2 s 14646 163200 14702 164400 6 la_input[4]
port 269 nsew signal input
rlabel metal2 s 169390 163200 169446 164400 6 la_input[50]
port 270 nsew signal input
rlabel metal2 s 172794 163200 172850 164400 6 la_input[51]
port 271 nsew signal input
rlabel metal2 s 176106 163200 176162 164400 6 la_input[52]
port 272 nsew signal input
rlabel metal2 s 179510 163200 179566 164400 6 la_input[53]
port 273 nsew signal input
rlabel metal2 s 182914 163200 182970 164400 6 la_input[54]
port 274 nsew signal input
rlabel metal2 s 186226 163200 186282 164400 6 la_input[55]
port 275 nsew signal input
rlabel metal2 s 189630 163200 189686 164400 6 la_input[56]
port 276 nsew signal input
rlabel metal2 s 192942 163200 192998 164400 6 la_input[57]
port 277 nsew signal input
rlabel metal2 s 196346 163200 196402 164400 6 la_input[58]
port 278 nsew signal input
rlabel metal2 s 199658 163200 199714 164400 6 la_input[59]
port 279 nsew signal input
rlabel metal2 s 18050 163200 18106 164400 6 la_input[5]
port 280 nsew signal input
rlabel metal2 s 203062 163200 203118 164400 6 la_input[60]
port 281 nsew signal input
rlabel metal2 s 206466 163200 206522 164400 6 la_input[61]
port 282 nsew signal input
rlabel metal2 s 209778 163200 209834 164400 6 la_input[62]
port 283 nsew signal input
rlabel metal2 s 213182 163200 213238 164400 6 la_input[63]
port 284 nsew signal input
rlabel metal2 s 216494 163200 216550 164400 6 la_input[64]
port 285 nsew signal input
rlabel metal2 s 219898 163200 219954 164400 6 la_input[65]
port 286 nsew signal input
rlabel metal2 s 223210 163200 223266 164400 6 la_input[66]
port 287 nsew signal input
rlabel metal2 s 226614 163200 226670 164400 6 la_input[67]
port 288 nsew signal input
rlabel metal2 s 230018 163200 230074 164400 6 la_input[68]
port 289 nsew signal input
rlabel metal2 s 233330 163200 233386 164400 6 la_input[69]
port 290 nsew signal input
rlabel metal2 s 21362 163200 21418 164400 6 la_input[6]
port 291 nsew signal input
rlabel metal2 s 236734 163200 236790 164400 6 la_input[70]
port 292 nsew signal input
rlabel metal2 s 240046 163200 240102 164400 6 la_input[71]
port 293 nsew signal input
rlabel metal2 s 243450 163200 243506 164400 6 la_input[72]
port 294 nsew signal input
rlabel metal2 s 246762 163200 246818 164400 6 la_input[73]
port 295 nsew signal input
rlabel metal2 s 250166 163200 250222 164400 6 la_input[74]
port 296 nsew signal input
rlabel metal2 s 253570 163200 253626 164400 6 la_input[75]
port 297 nsew signal input
rlabel metal2 s 256882 163200 256938 164400 6 la_input[76]
port 298 nsew signal input
rlabel metal2 s 260286 163200 260342 164400 6 la_input[77]
port 299 nsew signal input
rlabel metal2 s 263598 163200 263654 164400 6 la_input[78]
port 300 nsew signal input
rlabel metal2 s 267002 163200 267058 164400 6 la_input[79]
port 301 nsew signal input
rlabel metal2 s 24766 163200 24822 164400 6 la_input[7]
port 302 nsew signal input
rlabel metal2 s 270314 163200 270370 164400 6 la_input[80]
port 303 nsew signal input
rlabel metal2 s 273718 163200 273774 164400 6 la_input[81]
port 304 nsew signal input
rlabel metal2 s 277122 163200 277178 164400 6 la_input[82]
port 305 nsew signal input
rlabel metal2 s 280434 163200 280490 164400 6 la_input[83]
port 306 nsew signal input
rlabel metal2 s 283838 163200 283894 164400 6 la_input[84]
port 307 nsew signal input
rlabel metal2 s 287150 163200 287206 164400 6 la_input[85]
port 308 nsew signal input
rlabel metal2 s 290554 163200 290610 164400 6 la_input[86]
port 309 nsew signal input
rlabel metal2 s 293866 163200 293922 164400 6 la_input[87]
port 310 nsew signal input
rlabel metal2 s 297270 163200 297326 164400 6 la_input[88]
port 311 nsew signal input
rlabel metal2 s 300674 163200 300730 164400 6 la_input[89]
port 312 nsew signal input
rlabel metal2 s 28078 163200 28134 164400 6 la_input[8]
port 313 nsew signal input
rlabel metal2 s 303986 163200 304042 164400 6 la_input[90]
port 314 nsew signal input
rlabel metal2 s 307390 163200 307446 164400 6 la_input[91]
port 315 nsew signal input
rlabel metal2 s 310702 163200 310758 164400 6 la_input[92]
port 316 nsew signal input
rlabel metal2 s 314106 163200 314162 164400 6 la_input[93]
port 317 nsew signal input
rlabel metal2 s 317418 163200 317474 164400 6 la_input[94]
port 318 nsew signal input
rlabel metal2 s 320822 163200 320878 164400 6 la_input[95]
port 319 nsew signal input
rlabel metal2 s 324226 163200 324282 164400 6 la_input[96]
port 320 nsew signal input
rlabel metal2 s 327538 163200 327594 164400 6 la_input[97]
port 321 nsew signal input
rlabel metal2 s 330942 163200 330998 164400 6 la_input[98]
port 322 nsew signal input
rlabel metal2 s 334254 163200 334310 164400 6 la_input[99]
port 323 nsew signal input
rlabel metal2 s 31482 163200 31538 164400 6 la_input[9]
port 324 nsew signal input
rlabel metal2 s 2042 163200 2098 164400 6 la_oenb[0]
port 325 nsew signal tristate
rlabel metal2 s 338486 163200 338542 164400 6 la_oenb[100]
port 326 nsew signal tristate
rlabel metal2 s 341890 163200 341946 164400 6 la_oenb[101]
port 327 nsew signal tristate
rlabel metal2 s 345202 163200 345258 164400 6 la_oenb[102]
port 328 nsew signal tristate
rlabel metal2 s 348606 163200 348662 164400 6 la_oenb[103]
port 329 nsew signal tristate
rlabel metal2 s 351918 163200 351974 164400 6 la_oenb[104]
port 330 nsew signal tristate
rlabel metal2 s 355322 163200 355378 164400 6 la_oenb[105]
port 331 nsew signal tristate
rlabel metal2 s 358634 163200 358690 164400 6 la_oenb[106]
port 332 nsew signal tristate
rlabel metal2 s 362038 163200 362094 164400 6 la_oenb[107]
port 333 nsew signal tristate
rlabel metal2 s 365442 163200 365498 164400 6 la_oenb[108]
port 334 nsew signal tristate
rlabel metal2 s 368754 163200 368810 164400 6 la_oenb[109]
port 335 nsew signal tristate
rlabel metal2 s 35714 163200 35770 164400 6 la_oenb[10]
port 336 nsew signal tristate
rlabel metal2 s 372158 163200 372214 164400 6 la_oenb[110]
port 337 nsew signal tristate
rlabel metal2 s 375470 163200 375526 164400 6 la_oenb[111]
port 338 nsew signal tristate
rlabel metal2 s 378874 163200 378930 164400 6 la_oenb[112]
port 339 nsew signal tristate
rlabel metal2 s 382186 163200 382242 164400 6 la_oenb[113]
port 340 nsew signal tristate
rlabel metal2 s 385590 163200 385646 164400 6 la_oenb[114]
port 341 nsew signal tristate
rlabel metal2 s 388994 163200 389050 164400 6 la_oenb[115]
port 342 nsew signal tristate
rlabel metal2 s 392306 163200 392362 164400 6 la_oenb[116]
port 343 nsew signal tristate
rlabel metal2 s 395710 163200 395766 164400 6 la_oenb[117]
port 344 nsew signal tristate
rlabel metal2 s 399022 163200 399078 164400 6 la_oenb[118]
port 345 nsew signal tristate
rlabel metal2 s 402426 163200 402482 164400 6 la_oenb[119]
port 346 nsew signal tristate
rlabel metal2 s 39026 163200 39082 164400 6 la_oenb[11]
port 347 nsew signal tristate
rlabel metal2 s 405738 163200 405794 164400 6 la_oenb[120]
port 348 nsew signal tristate
rlabel metal2 s 409142 163200 409198 164400 6 la_oenb[121]
port 349 nsew signal tristate
rlabel metal2 s 412546 163200 412602 164400 6 la_oenb[122]
port 350 nsew signal tristate
rlabel metal2 s 415858 163200 415914 164400 6 la_oenb[123]
port 351 nsew signal tristate
rlabel metal2 s 419262 163200 419318 164400 6 la_oenb[124]
port 352 nsew signal tristate
rlabel metal2 s 422574 163200 422630 164400 6 la_oenb[125]
port 353 nsew signal tristate
rlabel metal2 s 425978 163200 426034 164400 6 la_oenb[126]
port 354 nsew signal tristate
rlabel metal2 s 429290 163200 429346 164400 6 la_oenb[127]
port 355 nsew signal tristate
rlabel metal2 s 42430 163200 42486 164400 6 la_oenb[12]
port 356 nsew signal tristate
rlabel metal2 s 45742 163200 45798 164400 6 la_oenb[13]
port 357 nsew signal tristate
rlabel metal2 s 49146 163200 49202 164400 6 la_oenb[14]
port 358 nsew signal tristate
rlabel metal2 s 52458 163200 52514 164400 6 la_oenb[15]
port 359 nsew signal tristate
rlabel metal2 s 55862 163200 55918 164400 6 la_oenb[16]
port 360 nsew signal tristate
rlabel metal2 s 59266 163200 59322 164400 6 la_oenb[17]
port 361 nsew signal tristate
rlabel metal2 s 62578 163200 62634 164400 6 la_oenb[18]
port 362 nsew signal tristate
rlabel metal2 s 65982 163200 66038 164400 6 la_oenb[19]
port 363 nsew signal tristate
rlabel metal2 s 5354 163200 5410 164400 6 la_oenb[1]
port 364 nsew signal tristate
rlabel metal2 s 69294 163200 69350 164400 6 la_oenb[20]
port 365 nsew signal tristate
rlabel metal2 s 72698 163200 72754 164400 6 la_oenb[21]
port 366 nsew signal tristate
rlabel metal2 s 76010 163200 76066 164400 6 la_oenb[22]
port 367 nsew signal tristate
rlabel metal2 s 79414 163200 79470 164400 6 la_oenb[23]
port 368 nsew signal tristate
rlabel metal2 s 82818 163200 82874 164400 6 la_oenb[24]
port 369 nsew signal tristate
rlabel metal2 s 86130 163200 86186 164400 6 la_oenb[25]
port 370 nsew signal tristate
rlabel metal2 s 89534 163200 89590 164400 6 la_oenb[26]
port 371 nsew signal tristate
rlabel metal2 s 92846 163200 92902 164400 6 la_oenb[27]
port 372 nsew signal tristate
rlabel metal2 s 96250 163200 96306 164400 6 la_oenb[28]
port 373 nsew signal tristate
rlabel metal2 s 99562 163200 99618 164400 6 la_oenb[29]
port 374 nsew signal tristate
rlabel metal2 s 8758 163200 8814 164400 6 la_oenb[2]
port 375 nsew signal tristate
rlabel metal2 s 102966 163200 103022 164400 6 la_oenb[30]
port 376 nsew signal tristate
rlabel metal2 s 106370 163200 106426 164400 6 la_oenb[31]
port 377 nsew signal tristate
rlabel metal2 s 109682 163200 109738 164400 6 la_oenb[32]
port 378 nsew signal tristate
rlabel metal2 s 113086 163200 113142 164400 6 la_oenb[33]
port 379 nsew signal tristate
rlabel metal2 s 116398 163200 116454 164400 6 la_oenb[34]
port 380 nsew signal tristate
rlabel metal2 s 119802 163200 119858 164400 6 la_oenb[35]
port 381 nsew signal tristate
rlabel metal2 s 123114 163200 123170 164400 6 la_oenb[36]
port 382 nsew signal tristate
rlabel metal2 s 126518 163200 126574 164400 6 la_oenb[37]
port 383 nsew signal tristate
rlabel metal2 s 129922 163200 129978 164400 6 la_oenb[38]
port 384 nsew signal tristate
rlabel metal2 s 133234 163200 133290 164400 6 la_oenb[39]
port 385 nsew signal tristate
rlabel metal2 s 12162 163200 12218 164400 6 la_oenb[3]
port 386 nsew signal tristate
rlabel metal2 s 136638 163200 136694 164400 6 la_oenb[40]
port 387 nsew signal tristate
rlabel metal2 s 139950 163200 140006 164400 6 la_oenb[41]
port 388 nsew signal tristate
rlabel metal2 s 143354 163200 143410 164400 6 la_oenb[42]
port 389 nsew signal tristate
rlabel metal2 s 146666 163200 146722 164400 6 la_oenb[43]
port 390 nsew signal tristate
rlabel metal2 s 150070 163200 150126 164400 6 la_oenb[44]
port 391 nsew signal tristate
rlabel metal2 s 153474 163200 153530 164400 6 la_oenb[45]
port 392 nsew signal tristate
rlabel metal2 s 156786 163200 156842 164400 6 la_oenb[46]
port 393 nsew signal tristate
rlabel metal2 s 160190 163200 160246 164400 6 la_oenb[47]
port 394 nsew signal tristate
rlabel metal2 s 163502 163200 163558 164400 6 la_oenb[48]
port 395 nsew signal tristate
rlabel metal2 s 166906 163200 166962 164400 6 la_oenb[49]
port 396 nsew signal tristate
rlabel metal2 s 15474 163200 15530 164400 6 la_oenb[4]
port 397 nsew signal tristate
rlabel metal2 s 170218 163200 170274 164400 6 la_oenb[50]
port 398 nsew signal tristate
rlabel metal2 s 173622 163200 173678 164400 6 la_oenb[51]
port 399 nsew signal tristate
rlabel metal2 s 177026 163200 177082 164400 6 la_oenb[52]
port 400 nsew signal tristate
rlabel metal2 s 180338 163200 180394 164400 6 la_oenb[53]
port 401 nsew signal tristate
rlabel metal2 s 183742 163200 183798 164400 6 la_oenb[54]
port 402 nsew signal tristate
rlabel metal2 s 187054 163200 187110 164400 6 la_oenb[55]
port 403 nsew signal tristate
rlabel metal2 s 190458 163200 190514 164400 6 la_oenb[56]
port 404 nsew signal tristate
rlabel metal2 s 193770 163200 193826 164400 6 la_oenb[57]
port 405 nsew signal tristate
rlabel metal2 s 197174 163200 197230 164400 6 la_oenb[58]
port 406 nsew signal tristate
rlabel metal2 s 200578 163200 200634 164400 6 la_oenb[59]
port 407 nsew signal tristate
rlabel metal2 s 18878 163200 18934 164400 6 la_oenb[5]
port 408 nsew signal tristate
rlabel metal2 s 203890 163200 203946 164400 6 la_oenb[60]
port 409 nsew signal tristate
rlabel metal2 s 207294 163200 207350 164400 6 la_oenb[61]
port 410 nsew signal tristate
rlabel metal2 s 210606 163200 210662 164400 6 la_oenb[62]
port 411 nsew signal tristate
rlabel metal2 s 214010 163200 214066 164400 6 la_oenb[63]
port 412 nsew signal tristate
rlabel metal2 s 217322 163200 217378 164400 6 la_oenb[64]
port 413 nsew signal tristate
rlabel metal2 s 220726 163200 220782 164400 6 la_oenb[65]
port 414 nsew signal tristate
rlabel metal2 s 224130 163200 224186 164400 6 la_oenb[66]
port 415 nsew signal tristate
rlabel metal2 s 227442 163200 227498 164400 6 la_oenb[67]
port 416 nsew signal tristate
rlabel metal2 s 230846 163200 230902 164400 6 la_oenb[68]
port 417 nsew signal tristate
rlabel metal2 s 234158 163200 234214 164400 6 la_oenb[69]
port 418 nsew signal tristate
rlabel metal2 s 22190 163200 22246 164400 6 la_oenb[6]
port 419 nsew signal tristate
rlabel metal2 s 237562 163200 237618 164400 6 la_oenb[70]
port 420 nsew signal tristate
rlabel metal2 s 240874 163200 240930 164400 6 la_oenb[71]
port 421 nsew signal tristate
rlabel metal2 s 244278 163200 244334 164400 6 la_oenb[72]
port 422 nsew signal tristate
rlabel metal2 s 247682 163200 247738 164400 6 la_oenb[73]
port 423 nsew signal tristate
rlabel metal2 s 250994 163200 251050 164400 6 la_oenb[74]
port 424 nsew signal tristate
rlabel metal2 s 254398 163200 254454 164400 6 la_oenb[75]
port 425 nsew signal tristate
rlabel metal2 s 257710 163200 257766 164400 6 la_oenb[76]
port 426 nsew signal tristate
rlabel metal2 s 261114 163200 261170 164400 6 la_oenb[77]
port 427 nsew signal tristate
rlabel metal2 s 264426 163200 264482 164400 6 la_oenb[78]
port 428 nsew signal tristate
rlabel metal2 s 267830 163200 267886 164400 6 la_oenb[79]
port 429 nsew signal tristate
rlabel metal2 s 25594 163200 25650 164400 6 la_oenb[7]
port 430 nsew signal tristate
rlabel metal2 s 271234 163200 271290 164400 6 la_oenb[80]
port 431 nsew signal tristate
rlabel metal2 s 274546 163200 274602 164400 6 la_oenb[81]
port 432 nsew signal tristate
rlabel metal2 s 277950 163200 278006 164400 6 la_oenb[82]
port 433 nsew signal tristate
rlabel metal2 s 281262 163200 281318 164400 6 la_oenb[83]
port 434 nsew signal tristate
rlabel metal2 s 284666 163200 284722 164400 6 la_oenb[84]
port 435 nsew signal tristate
rlabel metal2 s 287978 163200 288034 164400 6 la_oenb[85]
port 436 nsew signal tristate
rlabel metal2 s 291382 163200 291438 164400 6 la_oenb[86]
port 437 nsew signal tristate
rlabel metal2 s 294786 163200 294842 164400 6 la_oenb[87]
port 438 nsew signal tristate
rlabel metal2 s 298098 163200 298154 164400 6 la_oenb[88]
port 439 nsew signal tristate
rlabel metal2 s 301502 163200 301558 164400 6 la_oenb[89]
port 440 nsew signal tristate
rlabel metal2 s 28906 163200 28962 164400 6 la_oenb[8]
port 441 nsew signal tristate
rlabel metal2 s 304814 163200 304870 164400 6 la_oenb[90]
port 442 nsew signal tristate
rlabel metal2 s 308218 163200 308274 164400 6 la_oenb[91]
port 443 nsew signal tristate
rlabel metal2 s 311530 163200 311586 164400 6 la_oenb[92]
port 444 nsew signal tristate
rlabel metal2 s 314934 163200 314990 164400 6 la_oenb[93]
port 445 nsew signal tristate
rlabel metal2 s 318338 163200 318394 164400 6 la_oenb[94]
port 446 nsew signal tristate
rlabel metal2 s 321650 163200 321706 164400 6 la_oenb[95]
port 447 nsew signal tristate
rlabel metal2 s 325054 163200 325110 164400 6 la_oenb[96]
port 448 nsew signal tristate
rlabel metal2 s 328366 163200 328422 164400 6 la_oenb[97]
port 449 nsew signal tristate
rlabel metal2 s 331770 163200 331826 164400 6 la_oenb[98]
port 450 nsew signal tristate
rlabel metal2 s 335082 163200 335138 164400 6 la_oenb[99]
port 451 nsew signal tristate
rlabel metal2 s 32310 163200 32366 164400 6 la_oenb[9]
port 452 nsew signal tristate
rlabel metal2 s 2870 163200 2926 164400 6 la_output[0]
port 453 nsew signal tristate
rlabel metal2 s 339314 163200 339370 164400 6 la_output[100]
port 454 nsew signal tristate
rlabel metal2 s 342718 163200 342774 164400 6 la_output[101]
port 455 nsew signal tristate
rlabel metal2 s 346030 163200 346086 164400 6 la_output[102]
port 456 nsew signal tristate
rlabel metal2 s 349434 163200 349490 164400 6 la_output[103]
port 457 nsew signal tristate
rlabel metal2 s 352746 163200 352802 164400 6 la_output[104]
port 458 nsew signal tristate
rlabel metal2 s 356150 163200 356206 164400 6 la_output[105]
port 459 nsew signal tristate
rlabel metal2 s 359554 163200 359610 164400 6 la_output[106]
port 460 nsew signal tristate
rlabel metal2 s 362866 163200 362922 164400 6 la_output[107]
port 461 nsew signal tristate
rlabel metal2 s 366270 163200 366326 164400 6 la_output[108]
port 462 nsew signal tristate
rlabel metal2 s 369582 163200 369638 164400 6 la_output[109]
port 463 nsew signal tristate
rlabel metal2 s 36542 163200 36598 164400 6 la_output[10]
port 464 nsew signal tristate
rlabel metal2 s 372986 163200 373042 164400 6 la_output[110]
port 465 nsew signal tristate
rlabel metal2 s 376298 163200 376354 164400 6 la_output[111]
port 466 nsew signal tristate
rlabel metal2 s 379702 163200 379758 164400 6 la_output[112]
port 467 nsew signal tristate
rlabel metal2 s 383106 163200 383162 164400 6 la_output[113]
port 468 nsew signal tristate
rlabel metal2 s 386418 163200 386474 164400 6 la_output[114]
port 469 nsew signal tristate
rlabel metal2 s 389822 163200 389878 164400 6 la_output[115]
port 470 nsew signal tristate
rlabel metal2 s 393134 163200 393190 164400 6 la_output[116]
port 471 nsew signal tristate
rlabel metal2 s 396538 163200 396594 164400 6 la_output[117]
port 472 nsew signal tristate
rlabel metal2 s 399850 163200 399906 164400 6 la_output[118]
port 473 nsew signal tristate
rlabel metal2 s 403254 163200 403310 164400 6 la_output[119]
port 474 nsew signal tristate
rlabel metal2 s 39854 163200 39910 164400 6 la_output[11]
port 475 nsew signal tristate
rlabel metal2 s 406658 163200 406714 164400 6 la_output[120]
port 476 nsew signal tristate
rlabel metal2 s 409970 163200 410026 164400 6 la_output[121]
port 477 nsew signal tristate
rlabel metal2 s 413374 163200 413430 164400 6 la_output[122]
port 478 nsew signal tristate
rlabel metal2 s 416686 163200 416742 164400 6 la_output[123]
port 479 nsew signal tristate
rlabel metal2 s 420090 163200 420146 164400 6 la_output[124]
port 480 nsew signal tristate
rlabel metal2 s 423402 163200 423458 164400 6 la_output[125]
port 481 nsew signal tristate
rlabel metal2 s 426806 163200 426862 164400 6 la_output[126]
port 482 nsew signal tristate
rlabel metal2 s 430210 163200 430266 164400 6 la_output[127]
port 483 nsew signal tristate
rlabel metal2 s 43258 163200 43314 164400 6 la_output[12]
port 484 nsew signal tristate
rlabel metal2 s 46570 163200 46626 164400 6 la_output[13]
port 485 nsew signal tristate
rlabel metal2 s 49974 163200 50030 164400 6 la_output[14]
port 486 nsew signal tristate
rlabel metal2 s 53378 163200 53434 164400 6 la_output[15]
port 487 nsew signal tristate
rlabel metal2 s 56690 163200 56746 164400 6 la_output[16]
port 488 nsew signal tristate
rlabel metal2 s 60094 163200 60150 164400 6 la_output[17]
port 489 nsew signal tristate
rlabel metal2 s 63406 163200 63462 164400 6 la_output[18]
port 490 nsew signal tristate
rlabel metal2 s 66810 163200 66866 164400 6 la_output[19]
port 491 nsew signal tristate
rlabel metal2 s 6274 163200 6330 164400 6 la_output[1]
port 492 nsew signal tristate
rlabel metal2 s 70122 163200 70178 164400 6 la_output[20]
port 493 nsew signal tristate
rlabel metal2 s 73526 163200 73582 164400 6 la_output[21]
port 494 nsew signal tristate
rlabel metal2 s 76930 163200 76986 164400 6 la_output[22]
port 495 nsew signal tristate
rlabel metal2 s 80242 163200 80298 164400 6 la_output[23]
port 496 nsew signal tristate
rlabel metal2 s 83646 163200 83702 164400 6 la_output[24]
port 497 nsew signal tristate
rlabel metal2 s 86958 163200 87014 164400 6 la_output[25]
port 498 nsew signal tristate
rlabel metal2 s 90362 163200 90418 164400 6 la_output[26]
port 499 nsew signal tristate
rlabel metal2 s 93674 163200 93730 164400 6 la_output[27]
port 500 nsew signal tristate
rlabel metal2 s 97078 163200 97134 164400 6 la_output[28]
port 501 nsew signal tristate
rlabel metal2 s 100482 163200 100538 164400 6 la_output[29]
port 502 nsew signal tristate
rlabel metal2 s 9586 163200 9642 164400 6 la_output[2]
port 503 nsew signal tristate
rlabel metal2 s 103794 163200 103850 164400 6 la_output[30]
port 504 nsew signal tristate
rlabel metal2 s 107198 163200 107254 164400 6 la_output[31]
port 505 nsew signal tristate
rlabel metal2 s 110510 163200 110566 164400 6 la_output[32]
port 506 nsew signal tristate
rlabel metal2 s 113914 163200 113970 164400 6 la_output[33]
port 507 nsew signal tristate
rlabel metal2 s 117226 163200 117282 164400 6 la_output[34]
port 508 nsew signal tristate
rlabel metal2 s 120630 163200 120686 164400 6 la_output[35]
port 509 nsew signal tristate
rlabel metal2 s 124034 163200 124090 164400 6 la_output[36]
port 510 nsew signal tristate
rlabel metal2 s 127346 163200 127402 164400 6 la_output[37]
port 511 nsew signal tristate
rlabel metal2 s 130750 163200 130806 164400 6 la_output[38]
port 512 nsew signal tristate
rlabel metal2 s 134062 163200 134118 164400 6 la_output[39]
port 513 nsew signal tristate
rlabel metal2 s 12990 163200 13046 164400 6 la_output[3]
port 514 nsew signal tristate
rlabel metal2 s 137466 163200 137522 164400 6 la_output[40]
port 515 nsew signal tristate
rlabel metal2 s 140778 163200 140834 164400 6 la_output[41]
port 516 nsew signal tristate
rlabel metal2 s 144182 163200 144238 164400 6 la_output[42]
port 517 nsew signal tristate
rlabel metal2 s 147586 163200 147642 164400 6 la_output[43]
port 518 nsew signal tristate
rlabel metal2 s 150898 163200 150954 164400 6 la_output[44]
port 519 nsew signal tristate
rlabel metal2 s 154302 163200 154358 164400 6 la_output[45]
port 520 nsew signal tristate
rlabel metal2 s 157614 163200 157670 164400 6 la_output[46]
port 521 nsew signal tristate
rlabel metal2 s 161018 163200 161074 164400 6 la_output[47]
port 522 nsew signal tristate
rlabel metal2 s 164330 163200 164386 164400 6 la_output[48]
port 523 nsew signal tristate
rlabel metal2 s 167734 163200 167790 164400 6 la_output[49]
port 524 nsew signal tristate
rlabel metal2 s 16302 163200 16358 164400 6 la_output[4]
port 525 nsew signal tristate
rlabel metal2 s 171138 163200 171194 164400 6 la_output[50]
port 526 nsew signal tristate
rlabel metal2 s 174450 163200 174506 164400 6 la_output[51]
port 527 nsew signal tristate
rlabel metal2 s 177854 163200 177910 164400 6 la_output[52]
port 528 nsew signal tristate
rlabel metal2 s 181166 163200 181222 164400 6 la_output[53]
port 529 nsew signal tristate
rlabel metal2 s 184570 163200 184626 164400 6 la_output[54]
port 530 nsew signal tristate
rlabel metal2 s 187882 163200 187938 164400 6 la_output[55]
port 531 nsew signal tristate
rlabel metal2 s 191286 163200 191342 164400 6 la_output[56]
port 532 nsew signal tristate
rlabel metal2 s 194690 163200 194746 164400 6 la_output[57]
port 533 nsew signal tristate
rlabel metal2 s 198002 163200 198058 164400 6 la_output[58]
port 534 nsew signal tristate
rlabel metal2 s 201406 163200 201462 164400 6 la_output[59]
port 535 nsew signal tristate
rlabel metal2 s 19706 163200 19762 164400 6 la_output[5]
port 536 nsew signal tristate
rlabel metal2 s 204718 163200 204774 164400 6 la_output[60]
port 537 nsew signal tristate
rlabel metal2 s 208122 163200 208178 164400 6 la_output[61]
port 538 nsew signal tristate
rlabel metal2 s 211434 163200 211490 164400 6 la_output[62]
port 539 nsew signal tristate
rlabel metal2 s 214838 163200 214894 164400 6 la_output[63]
port 540 nsew signal tristate
rlabel metal2 s 218242 163200 218298 164400 6 la_output[64]
port 541 nsew signal tristate
rlabel metal2 s 221554 163200 221610 164400 6 la_output[65]
port 542 nsew signal tristate
rlabel metal2 s 224958 163200 225014 164400 6 la_output[66]
port 543 nsew signal tristate
rlabel metal2 s 228270 163200 228326 164400 6 la_output[67]
port 544 nsew signal tristate
rlabel metal2 s 231674 163200 231730 164400 6 la_output[68]
port 545 nsew signal tristate
rlabel metal2 s 234986 163200 235042 164400 6 la_output[69]
port 546 nsew signal tristate
rlabel metal2 s 23018 163200 23074 164400 6 la_output[6]
port 547 nsew signal tristate
rlabel metal2 s 238390 163200 238446 164400 6 la_output[70]
port 548 nsew signal tristate
rlabel metal2 s 241794 163200 241850 164400 6 la_output[71]
port 549 nsew signal tristate
rlabel metal2 s 245106 163200 245162 164400 6 la_output[72]
port 550 nsew signal tristate
rlabel metal2 s 248510 163200 248566 164400 6 la_output[73]
port 551 nsew signal tristate
rlabel metal2 s 251822 163200 251878 164400 6 la_output[74]
port 552 nsew signal tristate
rlabel metal2 s 255226 163200 255282 164400 6 la_output[75]
port 553 nsew signal tristate
rlabel metal2 s 258538 163200 258594 164400 6 la_output[76]
port 554 nsew signal tristate
rlabel metal2 s 261942 163200 261998 164400 6 la_output[77]
port 555 nsew signal tristate
rlabel metal2 s 265346 163200 265402 164400 6 la_output[78]
port 556 nsew signal tristate
rlabel metal2 s 268658 163200 268714 164400 6 la_output[79]
port 557 nsew signal tristate
rlabel metal2 s 26422 163200 26478 164400 6 la_output[7]
port 558 nsew signal tristate
rlabel metal2 s 272062 163200 272118 164400 6 la_output[80]
port 559 nsew signal tristate
rlabel metal2 s 275374 163200 275430 164400 6 la_output[81]
port 560 nsew signal tristate
rlabel metal2 s 278778 163200 278834 164400 6 la_output[82]
port 561 nsew signal tristate
rlabel metal2 s 282090 163200 282146 164400 6 la_output[83]
port 562 nsew signal tristate
rlabel metal2 s 285494 163200 285550 164400 6 la_output[84]
port 563 nsew signal tristate
rlabel metal2 s 288898 163200 288954 164400 6 la_output[85]
port 564 nsew signal tristate
rlabel metal2 s 292210 163200 292266 164400 6 la_output[86]
port 565 nsew signal tristate
rlabel metal2 s 295614 163200 295670 164400 6 la_output[87]
port 566 nsew signal tristate
rlabel metal2 s 298926 163200 298982 164400 6 la_output[88]
port 567 nsew signal tristate
rlabel metal2 s 302330 163200 302386 164400 6 la_output[89]
port 568 nsew signal tristate
rlabel metal2 s 29826 163200 29882 164400 6 la_output[8]
port 569 nsew signal tristate
rlabel metal2 s 305642 163200 305698 164400 6 la_output[90]
port 570 nsew signal tristate
rlabel metal2 s 309046 163200 309102 164400 6 la_output[91]
port 571 nsew signal tristate
rlabel metal2 s 312450 163200 312506 164400 6 la_output[92]
port 572 nsew signal tristate
rlabel metal2 s 315762 163200 315818 164400 6 la_output[93]
port 573 nsew signal tristate
rlabel metal2 s 319166 163200 319222 164400 6 la_output[94]
port 574 nsew signal tristate
rlabel metal2 s 322478 163200 322534 164400 6 la_output[95]
port 575 nsew signal tristate
rlabel metal2 s 325882 163200 325938 164400 6 la_output[96]
port 576 nsew signal tristate
rlabel metal2 s 329194 163200 329250 164400 6 la_output[97]
port 577 nsew signal tristate
rlabel metal2 s 332598 163200 332654 164400 6 la_output[98]
port 578 nsew signal tristate
rlabel metal2 s 336002 163200 336058 164400 6 la_output[99]
port 579 nsew signal tristate
rlabel metal2 s 33138 163200 33194 164400 6 la_output[9]
port 580 nsew signal tristate
rlabel metal2 s 431038 163200 431094 164400 6 mprj_ack_i
port 581 nsew signal input
rlabel metal2 s 435178 163200 435234 164400 6 mprj_adr_o[0]
port 582 nsew signal tristate
rlabel metal2 s 463790 163200 463846 164400 6 mprj_adr_o[10]
port 583 nsew signal tristate
rlabel metal2 s 466366 163200 466422 164400 6 mprj_adr_o[11]
port 584 nsew signal tristate
rlabel metal2 s 468850 163200 468906 164400 6 mprj_adr_o[12]
port 585 nsew signal tristate
rlabel metal2 s 471426 163200 471482 164400 6 mprj_adr_o[13]
port 586 nsew signal tristate
rlabel metal2 s 473910 163200 473966 164400 6 mprj_adr_o[14]
port 587 nsew signal tristate
rlabel metal2 s 476394 163200 476450 164400 6 mprj_adr_o[15]
port 588 nsew signal tristate
rlabel metal2 s 478970 163200 479026 164400 6 mprj_adr_o[16]
port 589 nsew signal tristate
rlabel metal2 s 481454 163200 481510 164400 6 mprj_adr_o[17]
port 590 nsew signal tristate
rlabel metal2 s 484030 163200 484086 164400 6 mprj_adr_o[18]
port 591 nsew signal tristate
rlabel metal2 s 486514 163200 486570 164400 6 mprj_adr_o[19]
port 592 nsew signal tristate
rlabel metal2 s 438582 163200 438638 164400 6 mprj_adr_o[1]
port 593 nsew signal tristate
rlabel metal2 s 489090 163200 489146 164400 6 mprj_adr_o[20]
port 594 nsew signal tristate
rlabel metal2 s 491574 163200 491630 164400 6 mprj_adr_o[21]
port 595 nsew signal tristate
rlabel metal2 s 494058 163200 494114 164400 6 mprj_adr_o[22]
port 596 nsew signal tristate
rlabel metal2 s 496634 163200 496690 164400 6 mprj_adr_o[23]
port 597 nsew signal tristate
rlabel metal2 s 499118 163200 499174 164400 6 mprj_adr_o[24]
port 598 nsew signal tristate
rlabel metal2 s 501694 163200 501750 164400 6 mprj_adr_o[25]
port 599 nsew signal tristate
rlabel metal2 s 504178 163200 504234 164400 6 mprj_adr_o[26]
port 600 nsew signal tristate
rlabel metal2 s 506754 163200 506810 164400 6 mprj_adr_o[27]
port 601 nsew signal tristate
rlabel metal2 s 509238 163200 509294 164400 6 mprj_adr_o[28]
port 602 nsew signal tristate
rlabel metal2 s 511722 163200 511778 164400 6 mprj_adr_o[29]
port 603 nsew signal tristate
rlabel metal2 s 441986 163200 442042 164400 6 mprj_adr_o[2]
port 604 nsew signal tristate
rlabel metal2 s 514298 163200 514354 164400 6 mprj_adr_o[30]
port 605 nsew signal tristate
rlabel metal2 s 516782 163200 516838 164400 6 mprj_adr_o[31]
port 606 nsew signal tristate
rlabel metal2 s 445298 163200 445354 164400 6 mprj_adr_o[3]
port 607 nsew signal tristate
rlabel metal2 s 448702 163200 448758 164400 6 mprj_adr_o[4]
port 608 nsew signal tristate
rlabel metal2 s 451186 163200 451242 164400 6 mprj_adr_o[5]
port 609 nsew signal tristate
rlabel metal2 s 453762 163200 453818 164400 6 mprj_adr_o[6]
port 610 nsew signal tristate
rlabel metal2 s 456246 163200 456302 164400 6 mprj_adr_o[7]
port 611 nsew signal tristate
rlabel metal2 s 458730 163200 458786 164400 6 mprj_adr_o[8]
port 612 nsew signal tristate
rlabel metal2 s 461306 163200 461362 164400 6 mprj_adr_o[9]
port 613 nsew signal tristate
rlabel metal2 s 431866 163200 431922 164400 6 mprj_cyc_o
port 614 nsew signal tristate
rlabel metal2 s 436098 163200 436154 164400 6 mprj_dat_i[0]
port 615 nsew signal input
rlabel metal2 s 464618 163200 464674 164400 6 mprj_dat_i[10]
port 616 nsew signal input
rlabel metal2 s 467194 163200 467250 164400 6 mprj_dat_i[11]
port 617 nsew signal input
rlabel metal2 s 469678 163200 469734 164400 6 mprj_dat_i[12]
port 618 nsew signal input
rlabel metal2 s 472254 163200 472310 164400 6 mprj_dat_i[13]
port 619 nsew signal input
rlabel metal2 s 474738 163200 474794 164400 6 mprj_dat_i[14]
port 620 nsew signal input
rlabel metal2 s 477314 163200 477370 164400 6 mprj_dat_i[15]
port 621 nsew signal input
rlabel metal2 s 479798 163200 479854 164400 6 mprj_dat_i[16]
port 622 nsew signal input
rlabel metal2 s 482282 163200 482338 164400 6 mprj_dat_i[17]
port 623 nsew signal input
rlabel metal2 s 484858 163200 484914 164400 6 mprj_dat_i[18]
port 624 nsew signal input
rlabel metal2 s 487342 163200 487398 164400 6 mprj_dat_i[19]
port 625 nsew signal input
rlabel metal2 s 439410 163200 439466 164400 6 mprj_dat_i[1]
port 626 nsew signal input
rlabel metal2 s 489918 163200 489974 164400 6 mprj_dat_i[20]
port 627 nsew signal input
rlabel metal2 s 492402 163200 492458 164400 6 mprj_dat_i[21]
port 628 nsew signal input
rlabel metal2 s 494978 163200 495034 164400 6 mprj_dat_i[22]
port 629 nsew signal input
rlabel metal2 s 497462 163200 497518 164400 6 mprj_dat_i[23]
port 630 nsew signal input
rlabel metal2 s 499946 163200 500002 164400 6 mprj_dat_i[24]
port 631 nsew signal input
rlabel metal2 s 502522 163200 502578 164400 6 mprj_dat_i[25]
port 632 nsew signal input
rlabel metal2 s 505006 163200 505062 164400 6 mprj_dat_i[26]
port 633 nsew signal input
rlabel metal2 s 507582 163200 507638 164400 6 mprj_dat_i[27]
port 634 nsew signal input
rlabel metal2 s 510066 163200 510122 164400 6 mprj_dat_i[28]
port 635 nsew signal input
rlabel metal2 s 512642 163200 512698 164400 6 mprj_dat_i[29]
port 636 nsew signal input
rlabel metal2 s 442814 163200 442870 164400 6 mprj_dat_i[2]
port 637 nsew signal input
rlabel metal2 s 515126 163200 515182 164400 6 mprj_dat_i[30]
port 638 nsew signal input
rlabel metal2 s 517610 163200 517666 164400 6 mprj_dat_i[31]
port 639 nsew signal input
rlabel metal2 s 446126 163200 446182 164400 6 mprj_dat_i[3]
port 640 nsew signal input
rlabel metal2 s 449530 163200 449586 164400 6 mprj_dat_i[4]
port 641 nsew signal input
rlabel metal2 s 452014 163200 452070 164400 6 mprj_dat_i[5]
port 642 nsew signal input
rlabel metal2 s 454590 163200 454646 164400 6 mprj_dat_i[6]
port 643 nsew signal input
rlabel metal2 s 457074 163200 457130 164400 6 mprj_dat_i[7]
port 644 nsew signal input
rlabel metal2 s 459650 163200 459706 164400 6 mprj_dat_i[8]
port 645 nsew signal input
rlabel metal2 s 462134 163200 462190 164400 6 mprj_dat_i[9]
port 646 nsew signal input
rlabel metal2 s 436926 163200 436982 164400 6 mprj_dat_o[0]
port 647 nsew signal tristate
rlabel metal2 s 465538 163200 465594 164400 6 mprj_dat_o[10]
port 648 nsew signal tristate
rlabel metal2 s 468022 163200 468078 164400 6 mprj_dat_o[11]
port 649 nsew signal tristate
rlabel metal2 s 470506 163200 470562 164400 6 mprj_dat_o[12]
port 650 nsew signal tristate
rlabel metal2 s 473082 163200 473138 164400 6 mprj_dat_o[13]
port 651 nsew signal tristate
rlabel metal2 s 475566 163200 475622 164400 6 mprj_dat_o[14]
port 652 nsew signal tristate
rlabel metal2 s 478142 163200 478198 164400 6 mprj_dat_o[15]
port 653 nsew signal tristate
rlabel metal2 s 480626 163200 480682 164400 6 mprj_dat_o[16]
port 654 nsew signal tristate
rlabel metal2 s 483202 163200 483258 164400 6 mprj_dat_o[17]
port 655 nsew signal tristate
rlabel metal2 s 485686 163200 485742 164400 6 mprj_dat_o[18]
port 656 nsew signal tristate
rlabel metal2 s 488170 163200 488226 164400 6 mprj_dat_o[19]
port 657 nsew signal tristate
rlabel metal2 s 440238 163200 440294 164400 6 mprj_dat_o[1]
port 658 nsew signal tristate
rlabel metal2 s 490746 163200 490802 164400 6 mprj_dat_o[20]
port 659 nsew signal tristate
rlabel metal2 s 493230 163200 493286 164400 6 mprj_dat_o[21]
port 660 nsew signal tristate
rlabel metal2 s 495806 163200 495862 164400 6 mprj_dat_o[22]
port 661 nsew signal tristate
rlabel metal2 s 498290 163200 498346 164400 6 mprj_dat_o[23]
port 662 nsew signal tristate
rlabel metal2 s 500866 163200 500922 164400 6 mprj_dat_o[24]
port 663 nsew signal tristate
rlabel metal2 s 503350 163200 503406 164400 6 mprj_dat_o[25]
port 664 nsew signal tristate
rlabel metal2 s 505834 163200 505890 164400 6 mprj_dat_o[26]
port 665 nsew signal tristate
rlabel metal2 s 508410 163200 508466 164400 6 mprj_dat_o[27]
port 666 nsew signal tristate
rlabel metal2 s 510894 163200 510950 164400 6 mprj_dat_o[28]
port 667 nsew signal tristate
rlabel metal2 s 513470 163200 513526 164400 6 mprj_dat_o[29]
port 668 nsew signal tristate
rlabel metal2 s 443642 163200 443698 164400 6 mprj_dat_o[2]
port 669 nsew signal tristate
rlabel metal2 s 515954 163200 516010 164400 6 mprj_dat_o[30]
port 670 nsew signal tristate
rlabel metal2 s 518530 163200 518586 164400 6 mprj_dat_o[31]
port 671 nsew signal tristate
rlabel metal2 s 446954 163200 447010 164400 6 mprj_dat_o[3]
port 672 nsew signal tristate
rlabel metal2 s 450358 163200 450414 164400 6 mprj_dat_o[4]
port 673 nsew signal tristate
rlabel metal2 s 452842 163200 452898 164400 6 mprj_dat_o[5]
port 674 nsew signal tristate
rlabel metal2 s 455418 163200 455474 164400 6 mprj_dat_o[6]
port 675 nsew signal tristate
rlabel metal2 s 457902 163200 457958 164400 6 mprj_dat_o[7]
port 676 nsew signal tristate
rlabel metal2 s 460478 163200 460534 164400 6 mprj_dat_o[8]
port 677 nsew signal tristate
rlabel metal2 s 462962 163200 463018 164400 6 mprj_dat_o[9]
port 678 nsew signal tristate
rlabel metal2 s 437754 163200 437810 164400 6 mprj_sel_o[0]
port 679 nsew signal tristate
rlabel metal2 s 441066 163200 441122 164400 6 mprj_sel_o[1]
port 680 nsew signal tristate
rlabel metal2 s 444470 163200 444526 164400 6 mprj_sel_o[2]
port 681 nsew signal tristate
rlabel metal2 s 447874 163200 447930 164400 6 mprj_sel_o[3]
port 682 nsew signal tristate
rlabel metal2 s 432694 163200 432750 164400 6 mprj_stb_o
port 683 nsew signal tristate
rlabel metal2 s 433522 163200 433578 164400 6 mprj_wb_iena
port 684 nsew signal tristate
rlabel metal2 s 434350 163200 434406 164400 6 mprj_we_o
port 685 nsew signal tristate
rlabel metal3 s 523200 89360 524400 89480 6 qspi_enabled
port 686 nsew signal tristate
rlabel metal3 s 523200 83376 524400 83496 6 ser_rx
port 687 nsew signal input
rlabel metal3 s 523200 84872 524400 84992 6 ser_tx
port 688 nsew signal tristate
rlabel metal3 s 523200 80384 524400 80504 6 spi_csb
port 689 nsew signal tristate
rlabel metal3 s 523200 86368 524400 86488 6 spi_enabled
port 690 nsew signal tristate
rlabel metal3 s 523200 78888 524400 79008 6 spi_sck
port 691 nsew signal tristate
rlabel metal3 s 523200 81880 524400 82000 6 spi_sdi
port 692 nsew signal input
rlabel metal3 s 523200 77392 524400 77512 6 spi_sdo
port 693 nsew signal tristate
rlabel metal3 s 523200 75896 524400 76016 6 spi_sdoenb
port 694 nsew signal tristate
rlabel metal3 s 523200 2184 524400 2304 6 sram_ro_addr[0]
port 695 nsew signal input
rlabel metal3 s 523200 3680 524400 3800 6 sram_ro_addr[1]
port 696 nsew signal input
rlabel metal3 s 523200 5176 524400 5296 6 sram_ro_addr[2]
port 697 nsew signal input
rlabel metal3 s 523200 6672 524400 6792 6 sram_ro_addr[3]
port 698 nsew signal input
rlabel metal3 s 523200 8168 524400 8288 6 sram_ro_addr[4]
port 699 nsew signal input
rlabel metal3 s 523200 9664 524400 9784 6 sram_ro_addr[5]
port 700 nsew signal input
rlabel metal3 s 523200 11160 524400 11280 6 sram_ro_addr[6]
port 701 nsew signal input
rlabel metal3 s 523200 12656 524400 12776 6 sram_ro_addr[7]
port 702 nsew signal input
rlabel metal3 s 523200 14152 524400 14272 6 sram_ro_clk
port 703 nsew signal input
rlabel metal3 s 523200 688 524400 808 6 sram_ro_csb
port 704 nsew signal input
rlabel metal3 s 523200 15648 524400 15768 6 sram_ro_data[0]
port 705 nsew signal tristate
rlabel metal3 s 523200 30744 524400 30864 6 sram_ro_data[10]
port 706 nsew signal tristate
rlabel metal3 s 523200 32240 524400 32360 6 sram_ro_data[11]
port 707 nsew signal tristate
rlabel metal3 s 523200 33736 524400 33856 6 sram_ro_data[12]
port 708 nsew signal tristate
rlabel metal3 s 523200 35232 524400 35352 6 sram_ro_data[13]
port 709 nsew signal tristate
rlabel metal3 s 523200 36728 524400 36848 6 sram_ro_data[14]
port 710 nsew signal tristate
rlabel metal3 s 523200 38224 524400 38344 6 sram_ro_data[15]
port 711 nsew signal tristate
rlabel metal3 s 523200 39720 524400 39840 6 sram_ro_data[16]
port 712 nsew signal tristate
rlabel metal3 s 523200 41216 524400 41336 6 sram_ro_data[17]
port 713 nsew signal tristate
rlabel metal3 s 523200 42712 524400 42832 6 sram_ro_data[18]
port 714 nsew signal tristate
rlabel metal3 s 523200 44208 524400 44328 6 sram_ro_data[19]
port 715 nsew signal tristate
rlabel metal3 s 523200 17144 524400 17264 6 sram_ro_data[1]
port 716 nsew signal tristate
rlabel metal3 s 523200 45704 524400 45824 6 sram_ro_data[20]
port 717 nsew signal tristate
rlabel metal3 s 523200 47200 524400 47320 6 sram_ro_data[21]
port 718 nsew signal tristate
rlabel metal3 s 523200 48832 524400 48952 6 sram_ro_data[22]
port 719 nsew signal tristate
rlabel metal3 s 523200 50328 524400 50448 6 sram_ro_data[23]
port 720 nsew signal tristate
rlabel metal3 s 523200 51824 524400 51944 6 sram_ro_data[24]
port 721 nsew signal tristate
rlabel metal3 s 523200 53320 524400 53440 6 sram_ro_data[25]
port 722 nsew signal tristate
rlabel metal3 s 523200 54816 524400 54936 6 sram_ro_data[26]
port 723 nsew signal tristate
rlabel metal3 s 523200 56312 524400 56432 6 sram_ro_data[27]
port 724 nsew signal tristate
rlabel metal3 s 523200 57808 524400 57928 6 sram_ro_data[28]
port 725 nsew signal tristate
rlabel metal3 s 523200 59304 524400 59424 6 sram_ro_data[29]
port 726 nsew signal tristate
rlabel metal3 s 523200 18640 524400 18760 6 sram_ro_data[2]
port 727 nsew signal tristate
rlabel metal3 s 523200 60800 524400 60920 6 sram_ro_data[30]
port 728 nsew signal tristate
rlabel metal3 s 523200 62296 524400 62416 6 sram_ro_data[31]
port 729 nsew signal tristate
rlabel metal3 s 523200 20136 524400 20256 6 sram_ro_data[3]
port 730 nsew signal tristate
rlabel metal3 s 523200 21632 524400 21752 6 sram_ro_data[4]
port 731 nsew signal tristate
rlabel metal3 s 523200 23128 524400 23248 6 sram_ro_data[5]
port 732 nsew signal tristate
rlabel metal3 s 523200 24760 524400 24880 6 sram_ro_data[6]
port 733 nsew signal tristate
rlabel metal3 s 523200 26256 524400 26376 6 sram_ro_data[7]
port 734 nsew signal tristate
rlabel metal3 s 523200 27752 524400 27872 6 sram_ro_data[8]
port 735 nsew signal tristate
rlabel metal3 s 523200 29248 524400 29368 6 sram_ro_data[9]
port 736 nsew signal tristate
rlabel metal3 s 523200 69776 524400 69896 6 trap
port 737 nsew signal tristate
rlabel metal3 s 523200 87864 524400 87984 6 uart_enabled
port 738 nsew signal tristate
rlabel metal2 s 519358 163200 519414 164400 6 user_irq_ena[0]
port 739 nsew signal tristate
rlabel metal2 s 520186 163200 520242 164400 6 user_irq_ena[1]
port 740 nsew signal tristate
rlabel metal2 s 521014 163200 521070 164400 6 user_irq_ena[2]
port 741 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 524000 164000
<< end >>
