magic
tech sky130A
magscale 1 2
timestamp 1665506905
<< obsli1 >>
rect 920 2159 98992 137649
<< obsm1 >>
rect 920 1708 99990 138032
<< metal2 >>
rect 2870 139200 2926 140000
rect 5906 139200 5962 140000
rect 8942 139200 8998 140000
rect 11978 139200 12034 140000
rect 15014 139200 15070 140000
rect 18050 139200 18106 140000
rect 21086 139200 21142 140000
rect 24122 139200 24178 140000
rect 27158 139200 27214 140000
rect 30194 139200 30250 140000
rect 33230 139200 33286 140000
rect 36266 139200 36322 140000
rect 39302 139200 39358 140000
rect 42338 139200 42394 140000
rect 45374 139200 45430 140000
rect 48410 139200 48466 140000
rect 51446 139200 51502 140000
rect 54482 139200 54538 140000
rect 57518 139200 57574 140000
rect 60554 139200 60610 140000
rect 63590 139200 63646 140000
rect 66626 139200 66682 140000
rect 69662 139200 69718 140000
rect 72698 139200 72754 140000
rect 75734 139200 75790 140000
rect 78770 139200 78826 140000
rect 81806 139200 81862 140000
rect 84842 139200 84898 140000
rect 87878 139200 87934 140000
rect 90914 139200 90970 140000
rect 93950 139200 94006 140000
rect 96986 139200 97042 140000
<< obsm2 >>
rect 1030 139144 2814 139346
rect 2982 139144 5850 139346
rect 6018 139144 8886 139346
rect 9054 139144 11922 139346
rect 12090 139144 14958 139346
rect 15126 139144 17994 139346
rect 18162 139144 21030 139346
rect 21198 139144 24066 139346
rect 24234 139144 27102 139346
rect 27270 139144 30138 139346
rect 30306 139144 33174 139346
rect 33342 139144 36210 139346
rect 36378 139144 39246 139346
rect 39414 139144 42282 139346
rect 42450 139144 45318 139346
rect 45486 139144 48354 139346
rect 48522 139144 51390 139346
rect 51558 139144 54426 139346
rect 54594 139144 57462 139346
rect 57630 139144 60498 139346
rect 60666 139144 63534 139346
rect 63702 139144 66570 139346
rect 66738 139144 69606 139346
rect 69774 139144 72642 139346
rect 72810 139144 75678 139346
rect 75846 139144 78714 139346
rect 78882 139144 81750 139346
rect 81918 139144 84786 139346
rect 84954 139144 87822 139346
rect 87990 139144 90858 139346
rect 91026 139144 93894 139346
rect 94062 139144 96930 139346
rect 97098 139144 99984 139346
rect 1030 1702 99984 139144
<< metal3 >>
rect 99200 137232 100000 137352
rect 99200 134240 100000 134360
rect 99200 131248 100000 131368
rect 99200 128256 100000 128376
rect 99200 125264 100000 125384
rect 99200 122272 100000 122392
rect 99200 119280 100000 119400
rect 99200 116288 100000 116408
rect 99200 113296 100000 113416
rect 99200 110304 100000 110424
rect 99200 107312 100000 107432
rect 99200 104320 100000 104440
rect 99200 101328 100000 101448
rect 99200 98336 100000 98456
rect 99200 95344 100000 95464
rect 99200 92352 100000 92472
rect 99200 89360 100000 89480
rect 99200 86368 100000 86488
rect 99200 83376 100000 83496
rect 99200 80384 100000 80504
rect 99200 77392 100000 77512
rect 99200 74400 100000 74520
rect 99200 71408 100000 71528
rect 99200 68416 100000 68536
rect 99200 65424 100000 65544
rect 99200 62432 100000 62552
rect 99200 59440 100000 59560
rect 99200 56448 100000 56568
rect 99200 53456 100000 53576
rect 99200 50464 100000 50584
rect 99200 47472 100000 47592
rect 99200 44480 100000 44600
rect 99200 41488 100000 41608
rect 99200 38496 100000 38616
rect 99200 35504 100000 35624
rect 99200 32512 100000 32632
rect 99200 29520 100000 29640
rect 99200 26528 100000 26648
rect 99200 23536 100000 23656
rect 99200 20544 100000 20664
rect 99200 17552 100000 17672
rect 99200 14560 100000 14680
rect 99200 11568 100000 11688
rect 99200 8576 100000 8696
rect 99200 5584 100000 5704
rect 99200 2592 100000 2712
<< obsm3 >>
rect 1025 137432 99807 137665
rect 1025 137152 99120 137432
rect 1025 134440 99807 137152
rect 1025 134160 99120 134440
rect 1025 131448 99807 134160
rect 1025 131168 99120 131448
rect 1025 128456 99807 131168
rect 1025 128176 99120 128456
rect 1025 125464 99807 128176
rect 1025 125184 99120 125464
rect 1025 122472 99807 125184
rect 1025 122192 99120 122472
rect 1025 119480 99807 122192
rect 1025 119200 99120 119480
rect 1025 116488 99807 119200
rect 1025 116208 99120 116488
rect 1025 113496 99807 116208
rect 1025 113216 99120 113496
rect 1025 110504 99807 113216
rect 1025 110224 99120 110504
rect 1025 107512 99807 110224
rect 1025 107232 99120 107512
rect 1025 104520 99807 107232
rect 1025 104240 99120 104520
rect 1025 101528 99807 104240
rect 1025 101248 99120 101528
rect 1025 98536 99807 101248
rect 1025 98256 99120 98536
rect 1025 95544 99807 98256
rect 1025 95264 99120 95544
rect 1025 92552 99807 95264
rect 1025 92272 99120 92552
rect 1025 89560 99807 92272
rect 1025 89280 99120 89560
rect 1025 86568 99807 89280
rect 1025 86288 99120 86568
rect 1025 83576 99807 86288
rect 1025 83296 99120 83576
rect 1025 80584 99807 83296
rect 1025 80304 99120 80584
rect 1025 77592 99807 80304
rect 1025 77312 99120 77592
rect 1025 74600 99807 77312
rect 1025 74320 99120 74600
rect 1025 71608 99807 74320
rect 1025 71328 99120 71608
rect 1025 68616 99807 71328
rect 1025 68336 99120 68616
rect 1025 65624 99807 68336
rect 1025 65344 99120 65624
rect 1025 62632 99807 65344
rect 1025 62352 99120 62632
rect 1025 59640 99807 62352
rect 1025 59360 99120 59640
rect 1025 56648 99807 59360
rect 1025 56368 99120 56648
rect 1025 53656 99807 56368
rect 1025 53376 99120 53656
rect 1025 50664 99807 53376
rect 1025 50384 99120 50664
rect 1025 47672 99807 50384
rect 1025 47392 99120 47672
rect 1025 44680 99807 47392
rect 1025 44400 99120 44680
rect 1025 41688 99807 44400
rect 1025 41408 99120 41688
rect 1025 38696 99807 41408
rect 1025 38416 99120 38696
rect 1025 35704 99807 38416
rect 1025 35424 99120 35704
rect 1025 32712 99807 35424
rect 1025 32432 99120 32712
rect 1025 29720 99807 32432
rect 1025 29440 99120 29720
rect 1025 26728 99807 29440
rect 1025 26448 99120 26728
rect 1025 23736 99807 26448
rect 1025 23456 99120 23736
rect 1025 20744 99807 23456
rect 1025 20464 99120 20744
rect 1025 17752 99807 20464
rect 1025 17472 99120 17752
rect 1025 14760 99807 17472
rect 1025 14480 99120 14760
rect 1025 11768 99807 14480
rect 1025 11488 99120 11768
rect 1025 8776 99807 11488
rect 1025 8496 99120 8776
rect 1025 5784 99807 8496
rect 1025 5504 99120 5784
rect 1025 2792 99807 5504
rect 1025 2512 99120 2792
rect 1025 1396 99807 2512
<< metal4 >>
rect -1260 -4 -940 139812
rect -600 656 -280 139152
rect 4024 -4 4344 139812
rect 19384 -4 19704 139812
rect 34744 -4 35064 139812
rect 50104 -4 50424 139812
rect 65464 -4 65784 139812
rect 80824 -4 81144 139812
rect 96184 -4 96504 139812
rect 100192 656 100512 139152
rect 100852 -4 101172 139812
<< obsm4 >>
rect 1347 1395 3944 136373
rect 4424 1395 19304 136373
rect 19784 1395 34664 136373
rect 35144 1395 50024 136373
rect 50504 1395 65384 136373
rect 65864 1395 80744 136373
rect 81224 1395 96104 136373
rect 96584 1395 97829 136373
<< metal5 >>
rect -1260 139492 101172 139812
rect -600 138832 100512 139152
rect -1260 135346 101172 135666
rect -1260 122346 101172 122666
rect -1260 109346 101172 109666
rect -1260 96346 101172 96666
rect -1260 83346 101172 83666
rect -1260 70346 101172 70666
rect -1260 57346 101172 57666
rect -1260 44346 101172 44666
rect -1260 31346 101172 31666
rect -1260 18346 101172 18666
rect -1260 5346 101172 5666
rect -600 656 100512 976
rect -1260 -4 101172 316
<< labels >>
rlabel metal3 s 99200 2592 100000 2712 6 A0[0]
port 1 nsew signal input
rlabel metal3 s 99200 5584 100000 5704 6 A0[1]
port 2 nsew signal input
rlabel metal3 s 99200 8576 100000 8696 6 A0[2]
port 3 nsew signal input
rlabel metal3 s 99200 11568 100000 11688 6 A0[3]
port 4 nsew signal input
rlabel metal3 s 99200 14560 100000 14680 6 A0[4]
port 5 nsew signal input
rlabel metal3 s 99200 17552 100000 17672 6 A0[5]
port 6 nsew signal input
rlabel metal3 s 99200 20544 100000 20664 6 A0[6]
port 7 nsew signal input
rlabel metal3 s 99200 23536 100000 23656 6 A0[7]
port 8 nsew signal input
rlabel metal3 s 99200 89360 100000 89480 6 CLK
port 9 nsew signal input
rlabel metal3 s 99200 41488 100000 41608 6 Di0[0]
port 10 nsew signal input
rlabel metal3 s 99200 71408 100000 71528 6 Di0[10]
port 11 nsew signal input
rlabel metal3 s 99200 74400 100000 74520 6 Di0[11]
port 12 nsew signal input
rlabel metal3 s 99200 77392 100000 77512 6 Di0[12]
port 13 nsew signal input
rlabel metal3 s 99200 80384 100000 80504 6 Di0[13]
port 14 nsew signal input
rlabel metal3 s 99200 83376 100000 83496 6 Di0[14]
port 15 nsew signal input
rlabel metal3 s 99200 86368 100000 86488 6 Di0[15]
port 16 nsew signal input
rlabel metal3 s 99200 92352 100000 92472 6 Di0[16]
port 17 nsew signal input
rlabel metal3 s 99200 95344 100000 95464 6 Di0[17]
port 18 nsew signal input
rlabel metal3 s 99200 98336 100000 98456 6 Di0[18]
port 19 nsew signal input
rlabel metal3 s 99200 101328 100000 101448 6 Di0[19]
port 20 nsew signal input
rlabel metal3 s 99200 44480 100000 44600 6 Di0[1]
port 21 nsew signal input
rlabel metal3 s 99200 104320 100000 104440 6 Di0[20]
port 22 nsew signal input
rlabel metal3 s 99200 107312 100000 107432 6 Di0[21]
port 23 nsew signal input
rlabel metal3 s 99200 110304 100000 110424 6 Di0[22]
port 24 nsew signal input
rlabel metal3 s 99200 113296 100000 113416 6 Di0[23]
port 25 nsew signal input
rlabel metal3 s 99200 116288 100000 116408 6 Di0[24]
port 26 nsew signal input
rlabel metal3 s 99200 119280 100000 119400 6 Di0[25]
port 27 nsew signal input
rlabel metal3 s 99200 122272 100000 122392 6 Di0[26]
port 28 nsew signal input
rlabel metal3 s 99200 125264 100000 125384 6 Di0[27]
port 29 nsew signal input
rlabel metal3 s 99200 128256 100000 128376 6 Di0[28]
port 30 nsew signal input
rlabel metal3 s 99200 131248 100000 131368 6 Di0[29]
port 31 nsew signal input
rlabel metal3 s 99200 47472 100000 47592 6 Di0[2]
port 32 nsew signal input
rlabel metal3 s 99200 134240 100000 134360 6 Di0[30]
port 33 nsew signal input
rlabel metal3 s 99200 137232 100000 137352 6 Di0[31]
port 34 nsew signal input
rlabel metal3 s 99200 50464 100000 50584 6 Di0[3]
port 35 nsew signal input
rlabel metal3 s 99200 53456 100000 53576 6 Di0[4]
port 36 nsew signal input
rlabel metal3 s 99200 56448 100000 56568 6 Di0[5]
port 37 nsew signal input
rlabel metal3 s 99200 59440 100000 59560 6 Di0[6]
port 38 nsew signal input
rlabel metal3 s 99200 62432 100000 62552 6 Di0[7]
port 39 nsew signal input
rlabel metal3 s 99200 65424 100000 65544 6 Di0[8]
port 40 nsew signal input
rlabel metal3 s 99200 68416 100000 68536 6 Di0[9]
port 41 nsew signal input
rlabel metal2 s 2870 139200 2926 140000 6 Do0[0]
port 42 nsew signal output
rlabel metal2 s 33230 139200 33286 140000 6 Do0[10]
port 43 nsew signal output
rlabel metal2 s 36266 139200 36322 140000 6 Do0[11]
port 44 nsew signal output
rlabel metal2 s 39302 139200 39358 140000 6 Do0[12]
port 45 nsew signal output
rlabel metal2 s 42338 139200 42394 140000 6 Do0[13]
port 46 nsew signal output
rlabel metal2 s 45374 139200 45430 140000 6 Do0[14]
port 47 nsew signal output
rlabel metal2 s 48410 139200 48466 140000 6 Do0[15]
port 48 nsew signal output
rlabel metal2 s 51446 139200 51502 140000 6 Do0[16]
port 49 nsew signal output
rlabel metal2 s 54482 139200 54538 140000 6 Do0[17]
port 50 nsew signal output
rlabel metal2 s 57518 139200 57574 140000 6 Do0[18]
port 51 nsew signal output
rlabel metal2 s 60554 139200 60610 140000 6 Do0[19]
port 52 nsew signal output
rlabel metal2 s 5906 139200 5962 140000 6 Do0[1]
port 53 nsew signal output
rlabel metal2 s 63590 139200 63646 140000 6 Do0[20]
port 54 nsew signal output
rlabel metal2 s 66626 139200 66682 140000 6 Do0[21]
port 55 nsew signal output
rlabel metal2 s 69662 139200 69718 140000 6 Do0[22]
port 56 nsew signal output
rlabel metal2 s 72698 139200 72754 140000 6 Do0[23]
port 57 nsew signal output
rlabel metal2 s 75734 139200 75790 140000 6 Do0[24]
port 58 nsew signal output
rlabel metal2 s 78770 139200 78826 140000 6 Do0[25]
port 59 nsew signal output
rlabel metal2 s 81806 139200 81862 140000 6 Do0[26]
port 60 nsew signal output
rlabel metal2 s 84842 139200 84898 140000 6 Do0[27]
port 61 nsew signal output
rlabel metal2 s 87878 139200 87934 140000 6 Do0[28]
port 62 nsew signal output
rlabel metal2 s 90914 139200 90970 140000 6 Do0[29]
port 63 nsew signal output
rlabel metal2 s 8942 139200 8998 140000 6 Do0[2]
port 64 nsew signal output
rlabel metal2 s 93950 139200 94006 140000 6 Do0[30]
port 65 nsew signal output
rlabel metal2 s 96986 139200 97042 140000 6 Do0[31]
port 66 nsew signal output
rlabel metal2 s 11978 139200 12034 140000 6 Do0[3]
port 67 nsew signal output
rlabel metal2 s 15014 139200 15070 140000 6 Do0[4]
port 68 nsew signal output
rlabel metal2 s 18050 139200 18106 140000 6 Do0[5]
port 69 nsew signal output
rlabel metal2 s 21086 139200 21142 140000 6 Do0[6]
port 70 nsew signal output
rlabel metal2 s 24122 139200 24178 140000 6 Do0[7]
port 71 nsew signal output
rlabel metal2 s 27158 139200 27214 140000 6 Do0[8]
port 72 nsew signal output
rlabel metal2 s 30194 139200 30250 140000 6 Do0[9]
port 73 nsew signal output
rlabel metal3 s 99200 38496 100000 38616 6 EN0
port 74 nsew signal input
rlabel metal4 s -1260 -4 -940 139812 4 VGND
port 75 nsew ground bidirectional
rlabel metal5 s -1260 -4 101172 316 6 VGND
port 75 nsew ground bidirectional
rlabel metal5 s -1260 139492 101172 139812 6 VGND
port 75 nsew ground bidirectional
rlabel metal4 s 100852 -4 101172 139812 6 VGND
port 75 nsew ground bidirectional
rlabel metal4 s 19384 -4 19704 139812 6 VGND
port 75 nsew ground bidirectional
rlabel metal4 s 50104 -4 50424 139812 6 VGND
port 75 nsew ground bidirectional
rlabel metal4 s 80824 -4 81144 139812 6 VGND
port 75 nsew ground bidirectional
rlabel metal5 s -1260 18346 101172 18666 6 VGND
port 75 nsew ground bidirectional
rlabel metal5 s -1260 44346 101172 44666 6 VGND
port 75 nsew ground bidirectional
rlabel metal5 s -1260 70346 101172 70666 6 VGND
port 75 nsew ground bidirectional
rlabel metal5 s -1260 96346 101172 96666 6 VGND
port 75 nsew ground bidirectional
rlabel metal5 s -1260 122346 101172 122666 6 VGND
port 75 nsew ground bidirectional
rlabel metal4 s -600 656 -280 139152 4 VPWR
port 76 nsew power bidirectional
rlabel metal5 s -600 656 100512 976 6 VPWR
port 76 nsew power bidirectional
rlabel metal5 s -600 138832 100512 139152 6 VPWR
port 76 nsew power bidirectional
rlabel metal4 s 100192 656 100512 139152 6 VPWR
port 76 nsew power bidirectional
rlabel metal4 s 4024 -4 4344 139812 6 VPWR
port 76 nsew power bidirectional
rlabel metal4 s 34744 -4 35064 139812 6 VPWR
port 76 nsew power bidirectional
rlabel metal4 s 65464 -4 65784 139812 6 VPWR
port 76 nsew power bidirectional
rlabel metal4 s 96184 -4 96504 139812 6 VPWR
port 76 nsew power bidirectional
rlabel metal5 s -1260 5346 101172 5666 6 VPWR
port 76 nsew power bidirectional
rlabel metal5 s -1260 31346 101172 31666 6 VPWR
port 76 nsew power bidirectional
rlabel metal5 s -1260 57346 101172 57666 6 VPWR
port 76 nsew power bidirectional
rlabel metal5 s -1260 83346 101172 83666 6 VPWR
port 76 nsew power bidirectional
rlabel metal5 s -1260 109346 101172 109666 6 VPWR
port 76 nsew power bidirectional
rlabel metal5 s -1260 135346 101172 135666 6 VPWR
port 76 nsew power bidirectional
rlabel metal3 s 99200 26528 100000 26648 6 WE0[0]
port 77 nsew signal input
rlabel metal3 s 99200 29520 100000 29640 6 WE0[1]
port 78 nsew signal input
rlabel metal3 s 99200 32512 100000 32632 6 WE0[2]
port 79 nsew signal input
rlabel metal3 s 99200 35504 100000 35624 6 WE0[3]
port 80 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 100000 140000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 56297974
string GDS_FILE /home/kareem_farid/caravel_mgmt_soc_litex/openlane/RAM256/runs/22_10_11_09_17/results/signoff/RAM256.magic.gds
string GDS_START 184572
<< end >>

