magic
tech sky130A
magscale 1 2
timestamp 1638311292
<< metal1 >>
rect 31386 158516 31392 158568
rect 31444 158556 31450 158568
rect 142706 158556 142712 158568
rect 31444 158528 142712 158556
rect 31444 158516 31450 158528
rect 142706 158516 142712 158528
rect 142764 158516 142770 158568
rect 96062 158448 96068 158500
rect 96120 158488 96126 158500
rect 192386 158488 192392 158500
rect 96120 158460 192392 158488
rect 96120 158448 96126 158460
rect 192386 158448 192392 158460
rect 192444 158448 192450 158500
rect 89346 158380 89352 158432
rect 89404 158420 89410 158432
rect 186682 158420 186688 158432
rect 89404 158392 186688 158420
rect 89404 158380 89410 158392
rect 186682 158380 186688 158392
rect 186740 158380 186746 158432
rect 82630 158312 82636 158364
rect 82688 158352 82694 158364
rect 182082 158352 182088 158364
rect 82688 158324 182088 158352
rect 82688 158312 82694 158324
rect 182082 158312 182088 158324
rect 182140 158312 182146 158364
rect 75914 158244 75920 158296
rect 75972 158284 75978 158296
rect 177022 158284 177028 158296
rect 75972 158256 177028 158284
rect 75972 158244 75978 158256
rect 177022 158244 177028 158256
rect 177080 158244 177086 158296
rect 69198 158176 69204 158228
rect 69256 158216 69262 158228
rect 171870 158216 171876 158228
rect 69256 158188 171876 158216
rect 69256 158176 69262 158188
rect 171870 158176 171876 158188
rect 171928 158176 171934 158228
rect 72602 158108 72608 158160
rect 72660 158148 72666 158160
rect 174446 158148 174452 158160
rect 72660 158120 174452 158148
rect 72660 158108 72666 158120
rect 174446 158108 174452 158120
rect 174504 158108 174510 158160
rect 65886 158040 65892 158092
rect 65944 158080 65950 158092
rect 169294 158080 169300 158092
rect 65944 158052 169300 158080
rect 65944 158040 65950 158052
rect 169294 158040 169300 158052
rect 169352 158040 169358 158092
rect 62482 157972 62488 158024
rect 62540 158012 62546 158024
rect 165982 158012 165988 158024
rect 62540 157984 165988 158012
rect 62540 157972 62546 157984
rect 165982 157972 165988 157984
rect 166040 157972 166046 158024
rect 59078 157904 59084 157956
rect 59136 157944 59142 157956
rect 163866 157944 163872 157956
rect 59136 157916 163872 157944
rect 59136 157904 59142 157916
rect 163866 157904 163872 157916
rect 163924 157904 163930 157956
rect 55766 157836 55772 157888
rect 55824 157876 55830 157888
rect 161658 157876 161664 157888
rect 55824 157848 161664 157876
rect 55824 157836 55830 157848
rect 161658 157836 161664 157848
rect 161716 157836 161722 157888
rect 52362 157768 52368 157820
rect 52420 157808 52426 157820
rect 158990 157808 158996 157820
rect 52420 157780 158996 157808
rect 52420 157768 52426 157780
rect 158990 157768 158996 157780
rect 159048 157768 159054 157820
rect 45646 157700 45652 157752
rect 45704 157740 45710 157752
rect 153746 157740 153752 157752
rect 45704 157712 153752 157740
rect 45704 157700 45710 157712
rect 153746 157700 153752 157712
rect 153804 157700 153810 157752
rect 49050 157632 49056 157684
rect 49108 157672 49114 157684
rect 156322 157672 156328 157684
rect 49108 157644 156328 157672
rect 49108 157632 49114 157644
rect 156322 157632 156328 157644
rect 156380 157632 156386 157684
rect 42334 157564 42340 157616
rect 42392 157604 42398 157616
rect 151262 157604 151268 157616
rect 42392 157576 151268 157604
rect 42392 157564 42398 157576
rect 151262 157564 151268 157576
rect 151320 157564 151326 157616
rect 38930 157496 38936 157548
rect 38988 157536 38994 157548
rect 147674 157536 147680 157548
rect 38988 157508 147680 157536
rect 38988 157496 38994 157508
rect 147674 157496 147680 157508
rect 147732 157496 147738 157548
rect 35618 157428 35624 157480
rect 35676 157468 35682 157480
rect 146202 157468 146208 157480
rect 35676 157440 146208 157468
rect 35676 157428 35682 157440
rect 146202 157428 146208 157440
rect 146260 157428 146266 157480
rect 102778 157360 102784 157412
rect 102836 157400 102842 157412
rect 197538 157400 197544 157412
rect 102836 157372 197544 157400
rect 102836 157360 102842 157372
rect 197538 157360 197544 157372
rect 197596 157360 197602 157412
rect 47394 157292 47400 157344
rect 47452 157332 47458 157344
rect 155126 157332 155132 157344
rect 47452 157304 155132 157332
rect 47452 157292 47458 157304
rect 155126 157292 155132 157304
rect 155184 157292 155190 157344
rect 156046 157292 156052 157344
rect 156104 157332 156110 157344
rect 160278 157332 160284 157344
rect 156104 157304 160284 157332
rect 156104 157292 156110 157304
rect 160278 157292 160284 157304
rect 160336 157292 160342 157344
rect 161934 157292 161940 157344
rect 161992 157332 161998 157344
rect 165430 157332 165436 157344
rect 161992 157304 165436 157332
rect 161992 157292 161998 157304
rect 165430 157292 165436 157304
rect 165488 157292 165494 157344
rect 172514 157292 172520 157344
rect 172572 157332 172578 157344
rect 250806 157332 250812 157344
rect 172572 157304 250812 157332
rect 172572 157292 172578 157304
rect 250806 157292 250812 157304
rect 250864 157292 250870 157344
rect 43990 157224 43996 157276
rect 44048 157264 44054 157276
rect 152550 157264 152556 157276
rect 44048 157236 152556 157264
rect 44048 157224 44054 157236
rect 152550 157224 152556 157236
rect 152608 157224 152614 157276
rect 155862 157224 155868 157276
rect 155920 157264 155926 157276
rect 162578 157264 162584 157276
rect 155920 157236 162584 157264
rect 155920 157224 155926 157236
rect 162578 157224 162584 157236
rect 162636 157224 162642 157276
rect 171686 157224 171692 157276
rect 171744 157264 171750 157276
rect 250162 157264 250168 157276
rect 171744 157236 250168 157264
rect 171744 157224 171750 157236
rect 250162 157224 250168 157236
rect 250220 157224 250226 157276
rect 37274 157156 37280 157208
rect 37332 157196 37338 157208
rect 146846 157196 146852 157208
rect 37332 157168 146852 157196
rect 37332 157156 37338 157168
rect 146846 157156 146852 157168
rect 146904 157156 146910 157208
rect 149974 157196 149980 157208
rect 146956 157168 149980 157196
rect 40678 157088 40684 157140
rect 40736 157128 40742 157140
rect 146956 157128 146984 157168
rect 149974 157156 149980 157168
rect 150032 157156 150038 157208
rect 152918 157156 152924 157208
rect 152976 157196 152982 157208
rect 157702 157196 157708 157208
rect 152976 157168 157708 157196
rect 152976 157156 152982 157168
rect 157702 157156 157708 157168
rect 157760 157156 157766 157208
rect 161566 157156 161572 157208
rect 161624 157196 161630 157208
rect 242434 157196 242440 157208
rect 161624 157168 242440 157196
rect 161624 157156 161630 157168
rect 242434 157156 242440 157168
rect 242492 157156 242498 157208
rect 40736 157100 146984 157128
rect 40736 157088 40742 157100
rect 148134 157088 148140 157140
rect 148192 157128 148198 157140
rect 148192 157100 156644 157128
rect 148192 157088 148198 157100
rect 28074 157020 28080 157072
rect 28132 157060 28138 157072
rect 140406 157060 140412 157072
rect 28132 157032 140412 157060
rect 28132 157020 28138 157032
rect 140406 157020 140412 157032
rect 140464 157020 140470 157072
rect 144822 157020 144828 157072
rect 144880 157060 144886 157072
rect 144880 157032 148272 157060
rect 144880 157020 144886 157032
rect 23842 156952 23848 157004
rect 23900 156992 23906 157004
rect 137094 156992 137100 157004
rect 23900 156964 137100 156992
rect 23900 156952 23906 156964
rect 137094 156952 137100 156964
rect 137152 156952 137158 157004
rect 143442 156952 143448 157004
rect 143500 156992 143506 157004
rect 148134 156992 148140 157004
rect 143500 156964 148140 156992
rect 143500 156952 143506 156964
rect 148134 156952 148140 156964
rect 148192 156952 148198 157004
rect 21358 156884 21364 156936
rect 21416 156924 21422 156936
rect 135346 156924 135352 156936
rect 21416 156896 135352 156924
rect 21416 156884 21422 156896
rect 135346 156884 135352 156896
rect 135404 156884 135410 156936
rect 138106 156884 138112 156936
rect 138164 156924 138170 156936
rect 148244 156924 148272 157032
rect 148318 157020 148324 157072
rect 148376 157060 148382 157072
rect 148376 157032 148456 157060
rect 148376 157020 148382 157032
rect 148428 156992 148456 157032
rect 151538 157020 151544 157072
rect 151596 157060 151602 157072
rect 156616 157060 156644 157100
rect 158254 157088 158260 157140
rect 158312 157128 158318 157140
rect 239950 157128 239956 157140
rect 158312 157100 239956 157128
rect 158312 157088 158318 157100
rect 239950 157088 239956 157100
rect 240008 157088 240014 157140
rect 232222 157060 232228 157072
rect 151596 157032 156552 157060
rect 156616 157032 232228 157060
rect 151596 157020 151602 157032
rect 156414 156992 156420 157004
rect 148428 156964 156420 156992
rect 156414 156952 156420 156964
rect 156472 156952 156478 157004
rect 156524 156992 156552 157032
rect 232222 157020 232228 157032
rect 232280 157020 232286 157072
rect 249794 157020 249800 157072
rect 249852 157060 249858 157072
rect 309870 157060 309876 157072
rect 249852 157032 309876 157060
rect 249852 157020 249858 157032
rect 309870 157020 309876 157032
rect 309928 157020 309934 157072
rect 234798 156992 234804 157004
rect 156524 156964 234804 156992
rect 234798 156952 234804 156964
rect 234856 156952 234862 157004
rect 243078 156952 243084 157004
rect 243136 156992 243142 157004
rect 304718 156992 304724 157004
rect 243136 156964 304724 156992
rect 243136 156952 243142 156964
rect 304718 156952 304724 156964
rect 304776 156952 304782 157004
rect 229554 156924 229560 156936
rect 138164 156896 146984 156924
rect 148244 156896 229560 156924
rect 138164 156884 138170 156896
rect 14642 156816 14648 156868
rect 14700 156856 14706 156868
rect 130102 156856 130108 156868
rect 14700 156828 130108 156856
rect 14700 156816 14706 156828
rect 130102 156816 130108 156828
rect 130160 156816 130166 156868
rect 141418 156816 141424 156868
rect 141476 156856 141482 156868
rect 146956 156856 146984 156896
rect 229554 156884 229560 156896
rect 229612 156884 229618 156936
rect 239674 156884 239680 156936
rect 239732 156924 239738 156936
rect 302234 156924 302240 156936
rect 239732 156896 302240 156924
rect 239732 156884 239738 156896
rect 302234 156884 302240 156896
rect 302292 156884 302298 156936
rect 224126 156856 224132 156868
rect 141476 156828 143580 156856
rect 146956 156828 224132 156856
rect 141476 156816 141482 156828
rect 7098 156748 7104 156800
rect 7156 156788 7162 156800
rect 7156 156760 122696 156788
rect 7156 156748 7162 156760
rect 3694 156680 3700 156732
rect 3752 156720 3758 156732
rect 121730 156720 121736 156732
rect 3752 156692 121736 156720
rect 3752 156680 3758 156692
rect 121730 156680 121736 156692
rect 121788 156680 121794 156732
rect 122668 156720 122696 156760
rect 122742 156748 122748 156800
rect 122800 156788 122806 156800
rect 143442 156788 143448 156800
rect 122800 156760 143448 156788
rect 122800 156748 122806 156760
rect 143442 156748 143448 156760
rect 143500 156748 143506 156800
rect 143552 156788 143580 156828
rect 224126 156816 224132 156828
rect 224184 156816 224190 156868
rect 226242 156816 226248 156868
rect 226300 156856 226306 156868
rect 291930 156856 291936 156868
rect 226300 156828 291936 156856
rect 226300 156816 226306 156828
rect 291930 156816 291936 156828
rect 291988 156816 291994 156868
rect 226886 156788 226892 156800
rect 143552 156760 226892 156788
rect 226886 156748 226892 156760
rect 226944 156748 226950 156800
rect 232958 156748 232964 156800
rect 233016 156788 233022 156800
rect 297082 156788 297088 156800
rect 233016 156760 297088 156788
rect 233016 156748 233022 156760
rect 297082 156748 297088 156760
rect 297140 156748 297146 156800
rect 124306 156720 124312 156732
rect 122668 156692 124312 156720
rect 124306 156680 124312 156692
rect 124364 156680 124370 156732
rect 131390 156680 131396 156732
rect 131448 156720 131454 156732
rect 218238 156720 218244 156732
rect 131448 156692 218244 156720
rect 131448 156680 131454 156692
rect 218238 156680 218244 156692
rect 218296 156680 218302 156732
rect 219526 156680 219532 156732
rect 219584 156720 219590 156732
rect 286778 156720 286784 156732
rect 219584 156692 286784 156720
rect 219584 156680 219590 156692
rect 286778 156680 286784 156692
rect 286836 156680 286842 156732
rect 382 156612 388 156664
rect 440 156652 446 156664
rect 118970 156652 118976 156664
rect 440 156624 118976 156652
rect 440 156612 446 156624
rect 118970 156612 118976 156624
rect 119028 156612 119034 156664
rect 124582 156612 124588 156664
rect 124640 156652 124646 156664
rect 214190 156652 214196 156664
rect 124640 156624 214196 156652
rect 124640 156612 124646 156624
rect 214190 156612 214196 156624
rect 214248 156612 214254 156664
rect 216122 156612 216128 156664
rect 216180 156652 216186 156664
rect 284110 156652 284116 156664
rect 216180 156624 284116 156652
rect 216180 156612 216186 156624
rect 284110 156612 284116 156624
rect 284168 156612 284174 156664
rect 50706 156544 50712 156596
rect 50764 156584 50770 156596
rect 152918 156584 152924 156596
rect 50764 156556 152924 156584
rect 50764 156544 50770 156556
rect 152918 156544 152924 156556
rect 152976 156544 152982 156596
rect 153010 156544 153016 156596
rect 153068 156584 153074 156596
rect 207842 156584 207848 156596
rect 153068 156556 207848 156584
rect 153068 156544 153074 156556
rect 207842 156544 207848 156556
rect 207900 156544 207906 156596
rect 54110 156476 54116 156528
rect 54168 156516 54174 156528
rect 156046 156516 156052 156528
rect 54168 156488 156052 156516
rect 54168 156476 54174 156488
rect 156046 156476 156052 156488
rect 156104 156476 156110 156528
rect 156414 156476 156420 156528
rect 156472 156516 156478 156528
rect 162118 156516 162124 156528
rect 156472 156488 162124 156516
rect 156472 156476 156478 156488
rect 162118 156476 162124 156488
rect 162176 156476 162182 156528
rect 173066 156516 173072 156528
rect 162320 156488 173072 156516
rect 60826 156408 60832 156460
rect 60884 156448 60890 156460
rect 161934 156448 161940 156460
rect 60884 156420 161940 156448
rect 60884 156408 60890 156420
rect 161934 156408 161940 156420
rect 161992 156408 161998 156460
rect 70854 156340 70860 156392
rect 70912 156380 70918 156392
rect 162320 156380 162348 156488
rect 173066 156476 173072 156488
rect 173124 156476 173130 156528
rect 174538 156476 174544 156528
rect 174596 156516 174602 156528
rect 178034 156516 178040 156528
rect 174596 156488 178040 156516
rect 174596 156476 174602 156488
rect 178034 156476 178040 156488
rect 178092 156476 178098 156528
rect 179230 156476 179236 156528
rect 179288 156516 179294 156528
rect 255958 156516 255964 156528
rect 179288 156488 255964 156516
rect 179288 156476 179294 156488
rect 255958 156476 255964 156488
rect 256016 156476 256022 156528
rect 162578 156408 162584 156460
rect 162636 156448 162642 156460
rect 176194 156448 176200 156460
rect 162636 156420 176200 156448
rect 162636 156408 162642 156420
rect 176194 156408 176200 156420
rect 176252 156408 176258 156460
rect 176286 156408 176292 156460
rect 176344 156448 176350 156460
rect 178954 156448 178960 156460
rect 176344 156420 178960 156448
rect 176344 156408 176350 156420
rect 178954 156408 178960 156420
rect 179012 156408 179018 156460
rect 183370 156408 183376 156460
rect 183428 156448 183434 156460
rect 259178 156448 259184 156460
rect 183428 156420 259184 156448
rect 183428 156408 183434 156420
rect 259178 156408 259184 156420
rect 259236 156408 259242 156460
rect 321094 156408 321100 156460
rect 321152 156448 321158 156460
rect 327258 156448 327264 156460
rect 321152 156420 327264 156448
rect 321152 156408 321158 156420
rect 327258 156408 327264 156420
rect 327316 156408 327322 156460
rect 70912 156352 162348 156380
rect 70912 156340 70918 156352
rect 162486 156340 162492 156392
rect 162544 156380 162550 156392
rect 175826 156380 175832 156392
rect 162544 156352 175832 156380
rect 162544 156340 162550 156352
rect 175826 156340 175832 156352
rect 175884 156340 175890 156392
rect 181162 156380 181168 156392
rect 176212 156352 181168 156380
rect 78398 156272 78404 156324
rect 78456 156312 78462 156324
rect 175918 156312 175924 156324
rect 78456 156284 175924 156312
rect 78456 156272 78462 156284
rect 175918 156272 175924 156284
rect 175976 156272 175982 156324
rect 176212 156312 176240 156352
rect 181162 156340 181168 156352
rect 181220 156340 181226 156392
rect 185118 156340 185124 156392
rect 185176 156380 185182 156392
rect 260006 156380 260012 156392
rect 185176 156352 260012 156380
rect 185176 156340 185182 156352
rect 260006 156340 260012 156352
rect 260064 156340 260070 156392
rect 176120 156284 176240 156312
rect 80974 156204 80980 156256
rect 81032 156244 81038 156256
rect 176120 156244 176148 156284
rect 178402 156272 178408 156324
rect 178460 156312 178466 156324
rect 178460 156284 185624 156312
rect 178460 156272 178466 156284
rect 81032 156216 176148 156244
rect 81032 156204 81038 156216
rect 176194 156204 176200 156256
rect 176252 156244 176258 156256
rect 176252 156216 185532 156244
rect 176252 156204 176258 156216
rect 121270 156136 121276 156188
rect 121328 156176 121334 156188
rect 185302 156176 185308 156188
rect 121328 156148 185308 156176
rect 121328 156136 121334 156148
rect 185302 156136 185308 156148
rect 185360 156136 185366 156188
rect 87690 156068 87696 156120
rect 87748 156108 87754 156120
rect 185394 156108 185400 156120
rect 87748 156080 185400 156108
rect 87748 156068 87754 156080
rect 185394 156068 185400 156080
rect 185452 156068 185458 156120
rect 185504 156108 185532 156216
rect 185596 156176 185624 156284
rect 185762 156272 185768 156324
rect 185820 156312 185826 156324
rect 189810 156312 189816 156324
rect 185820 156284 189816 156312
rect 185820 156272 185826 156284
rect 189810 156272 189816 156284
rect 189868 156272 189874 156324
rect 195146 156272 195152 156324
rect 195204 156312 195210 156324
rect 268102 156312 268108 156324
rect 195204 156284 268108 156312
rect 195204 156272 195210 156284
rect 268102 156272 268108 156284
rect 268160 156272 268166 156324
rect 185670 156204 185676 156256
rect 185728 156244 185734 156256
rect 191282 156244 191288 156256
rect 185728 156216 191288 156244
rect 185728 156204 185734 156216
rect 191282 156204 191288 156216
rect 191340 156204 191346 156256
rect 192662 156204 192668 156256
rect 192720 156244 192726 156256
rect 265158 156244 265164 156256
rect 192720 156216 265164 156244
rect 192720 156204 192726 156216
rect 265158 156204 265164 156216
rect 265216 156204 265222 156256
rect 255406 156176 255412 156188
rect 185596 156148 255412 156176
rect 255406 156136 255412 156148
rect 255464 156136 255470 156188
rect 223206 156108 223212 156120
rect 185504 156080 223212 156108
rect 223206 156068 223212 156080
rect 223264 156068 223270 156120
rect 94406 156000 94412 156052
rect 94464 156040 94470 156052
rect 185670 156040 185676 156052
rect 94464 156012 185676 156040
rect 94464 156000 94470 156012
rect 185670 156000 185676 156012
rect 185728 156000 185734 156052
rect 333606 156040 333612 156052
rect 328426 156012 333612 156040
rect 77570 155932 77576 155984
rect 77628 155972 77634 155984
rect 174538 155972 174544 155984
rect 77628 155944 174544 155972
rect 77628 155932 77634 155944
rect 174538 155932 174544 155944
rect 174596 155932 174602 155984
rect 175826 155932 175832 155984
rect 175884 155972 175890 155984
rect 205174 155972 205180 155984
rect 175884 155944 205180 155972
rect 175884 155932 175890 155944
rect 205174 155932 205180 155944
rect 205232 155932 205238 155984
rect 209774 155972 209780 155984
rect 209424 155944 209780 155972
rect 15470 155864 15476 155916
rect 15528 155904 15534 155916
rect 84194 155904 84200 155916
rect 15528 155876 84200 155904
rect 15528 155864 15534 155876
rect 84194 155864 84200 155876
rect 84252 155864 84258 155916
rect 84286 155864 84292 155916
rect 84344 155904 84350 155916
rect 85390 155904 85396 155916
rect 84344 155876 85396 155904
rect 84344 155864 84350 155876
rect 85390 155864 85396 155876
rect 85448 155864 85454 155916
rect 95234 155864 95240 155916
rect 95292 155904 95298 155916
rect 96522 155904 96528 155916
rect 95292 155876 96528 155904
rect 95292 155864 95298 155876
rect 96522 155864 96528 155876
rect 96580 155864 96586 155916
rect 101122 155864 101128 155916
rect 101180 155904 101186 155916
rect 102042 155904 102048 155916
rect 101180 155876 102048 155904
rect 101180 155864 101186 155876
rect 102042 155864 102048 155876
rect 102100 155864 102106 155916
rect 106182 155864 106188 155916
rect 106240 155904 106246 155916
rect 109402 155904 109408 155916
rect 106240 155876 109408 155904
rect 106240 155864 106246 155876
rect 109402 155864 109408 155876
rect 109460 155864 109466 155916
rect 109494 155864 109500 155916
rect 109552 155904 109558 155916
rect 111610 155904 111616 155916
rect 109552 155876 111616 155904
rect 109552 155864 109558 155876
rect 111610 155864 111616 155876
rect 111668 155864 111674 155916
rect 111794 155864 111800 155916
rect 111852 155904 111858 155916
rect 195698 155904 195704 155916
rect 111852 155876 195704 155904
rect 111852 155864 111858 155876
rect 195698 155864 195704 155876
rect 195756 155864 195762 155916
rect 200666 155904 200672 155916
rect 195808 155876 200672 155904
rect 26206 155808 64874 155836
rect 12066 155660 12072 155712
rect 12124 155700 12130 155712
rect 26206 155700 26234 155808
rect 12124 155672 26234 155700
rect 64846 155700 64874 155808
rect 76742 155796 76748 155848
rect 76800 155836 76806 155848
rect 76800 155808 82952 155836
rect 76800 155796 76806 155808
rect 66714 155728 66720 155780
rect 66772 155768 66778 155780
rect 82814 155768 82820 155780
rect 66772 155740 82820 155768
rect 66772 155728 66778 155740
rect 82814 155728 82820 155740
rect 82872 155728 82878 155780
rect 77110 155700 77116 155712
rect 64846 155672 77116 155700
rect 12124 155660 12130 155672
rect 77110 155660 77116 155672
rect 77168 155660 77174 155712
rect 81802 155660 81808 155712
rect 81860 155700 81866 155712
rect 82722 155700 82728 155712
rect 81860 155672 82728 155700
rect 81860 155660 81866 155672
rect 82722 155660 82728 155672
rect 82780 155660 82786 155712
rect 82924 155700 82952 155808
rect 83458 155796 83464 155848
rect 83516 155836 83522 155848
rect 173434 155836 173440 155848
rect 83516 155808 173440 155836
rect 83516 155796 83522 155808
rect 173434 155796 173440 155808
rect 173492 155796 173498 155848
rect 175642 155836 175648 155848
rect 173544 155808 175648 155836
rect 82998 155728 83004 155780
rect 83056 155768 83062 155780
rect 152918 155768 152924 155780
rect 83056 155740 152924 155768
rect 83056 155728 83062 155740
rect 152918 155728 152924 155740
rect 152976 155728 152982 155780
rect 153654 155728 153660 155780
rect 153712 155768 153718 155780
rect 156690 155768 156696 155780
rect 153712 155740 156696 155768
rect 153712 155728 153718 155740
rect 156690 155728 156696 155740
rect 156748 155728 156754 155780
rect 158806 155728 158812 155780
rect 158864 155768 158870 155780
rect 173544 155768 173572 155808
rect 175642 155796 175648 155808
rect 175700 155796 175706 155848
rect 175826 155796 175832 155848
rect 175884 155836 175890 155848
rect 177758 155836 177764 155848
rect 175884 155808 177764 155836
rect 175884 155796 175890 155808
rect 177758 155796 177764 155808
rect 177816 155796 177822 155848
rect 180058 155796 180064 155848
rect 180116 155836 180122 155848
rect 185486 155836 185492 155848
rect 180116 155808 185492 155836
rect 180116 155796 180122 155808
rect 185486 155796 185492 155808
rect 185544 155796 185550 155848
rect 187510 155836 187516 155848
rect 185596 155808 187516 155836
rect 158864 155740 173572 155768
rect 158864 155728 158870 155740
rect 174170 155728 174176 155780
rect 174228 155768 174234 155780
rect 174228 155740 177528 155768
rect 174228 155728 174234 155740
rect 164234 155700 164240 155712
rect 82924 155672 152964 155700
rect 49878 155592 49884 155644
rect 49936 155632 49942 155644
rect 134610 155632 134616 155644
rect 49936 155604 134616 155632
rect 49936 155592 49942 155604
rect 134610 155592 134616 155604
rect 134668 155592 134674 155644
rect 134702 155592 134708 155644
rect 134760 155632 134766 155644
rect 135162 155632 135168 155644
rect 134760 155604 135168 155632
rect 134760 155592 134766 155604
rect 135162 155592 135168 155604
rect 135220 155592 135226 155644
rect 136358 155592 136364 155644
rect 136416 155632 136422 155644
rect 146938 155632 146944 155644
rect 136416 155604 146944 155632
rect 136416 155592 136422 155604
rect 146938 155592 146944 155604
rect 146996 155592 147002 155644
rect 152936 155632 152964 155672
rect 153212 155672 164240 155700
rect 153212 155632 153240 155672
rect 164234 155660 164240 155672
rect 164292 155660 164298 155712
rect 164344 155672 166994 155700
rect 152936 155604 153240 155632
rect 153286 155592 153292 155644
rect 153344 155632 153350 155644
rect 164344 155632 164372 155672
rect 153344 155604 164372 155632
rect 166966 155632 166994 155672
rect 167454 155660 167460 155712
rect 167512 155700 167518 155712
rect 171042 155700 171048 155712
rect 167512 155672 171048 155700
rect 167512 155660 167518 155672
rect 171042 155660 171048 155672
rect 171100 155660 171106 155712
rect 171134 155660 171140 155712
rect 171192 155700 171198 155712
rect 176010 155700 176016 155712
rect 171192 155672 176016 155700
rect 171192 155660 171198 155672
rect 176010 155660 176016 155672
rect 176068 155660 176074 155712
rect 177500 155700 177528 155740
rect 177574 155728 177580 155780
rect 177632 155768 177638 155780
rect 185596 155768 185624 155808
rect 187510 155796 187516 155808
rect 187568 155796 187574 155848
rect 187602 155796 187608 155848
rect 187660 155836 187666 155848
rect 187660 155808 191236 155836
rect 187660 155796 187666 155808
rect 177632 155740 185624 155768
rect 177632 155728 177638 155740
rect 185670 155728 185676 155780
rect 185728 155768 185734 155780
rect 191098 155768 191104 155780
rect 185728 155740 191104 155768
rect 185728 155728 185734 155740
rect 191098 155728 191104 155740
rect 191156 155728 191162 155780
rect 191208 155768 191236 155808
rect 194318 155796 194324 155848
rect 194376 155836 194382 155848
rect 195808 155836 195836 155876
rect 200666 155864 200672 155876
rect 200724 155864 200730 155916
rect 200758 155864 200764 155916
rect 200816 155904 200822 155916
rect 205910 155904 205916 155916
rect 200816 155876 205916 155904
rect 200816 155864 200822 155876
rect 205910 155864 205916 155876
rect 205968 155864 205974 155916
rect 206922 155864 206928 155916
rect 206980 155904 206986 155916
rect 209424 155904 209452 155944
rect 209774 155932 209780 155944
rect 209832 155932 209838 155984
rect 244550 155932 244556 155984
rect 244608 155972 244614 155984
rect 246298 155972 246304 155984
rect 244608 155944 246304 155972
rect 244608 155932 244614 155944
rect 246298 155932 246304 155944
rect 246356 155932 246362 155984
rect 283006 155972 283012 155984
rect 281552 155944 283012 155972
rect 270218 155904 270224 155916
rect 206980 155876 209452 155904
rect 209608 155876 270224 155904
rect 206980 155864 206986 155876
rect 200298 155836 200304 155848
rect 194376 155808 195836 155836
rect 196728 155808 200304 155836
rect 194376 155796 194382 155808
rect 196728 155768 196756 155808
rect 200298 155796 200304 155808
rect 200356 155796 200362 155848
rect 201034 155796 201040 155848
rect 201092 155836 201098 155848
rect 209608 155836 209636 155876
rect 270218 155864 270224 155876
rect 270276 155864 270282 155916
rect 270770 155864 270776 155916
rect 270828 155904 270834 155916
rect 277210 155904 277216 155916
rect 270828 155876 277216 155904
rect 270828 155864 270834 155876
rect 277210 155864 277216 155876
rect 277268 155864 277274 155916
rect 281552 155904 281580 155944
rect 283006 155932 283012 155944
rect 283064 155932 283070 155984
rect 292206 155932 292212 155984
rect 292264 155972 292270 155984
rect 295794 155972 295800 155984
rect 292264 155944 295800 155972
rect 292264 155932 292270 155944
rect 295794 155932 295800 155944
rect 295852 155932 295858 155984
rect 321370 155932 321376 155984
rect 321428 155972 321434 155984
rect 321554 155972 321560 155984
rect 321428 155944 321560 155972
rect 321428 155932 321434 155944
rect 321554 155932 321560 155944
rect 321612 155932 321618 155984
rect 324498 155932 324504 155984
rect 324556 155972 324562 155984
rect 326614 155972 326620 155984
rect 324556 155944 326620 155972
rect 324556 155932 324562 155944
rect 326614 155932 326620 155944
rect 326672 155932 326678 155984
rect 277366 155876 281580 155904
rect 201092 155808 209636 155836
rect 201092 155796 201098 155808
rect 209682 155796 209688 155848
rect 209740 155836 209746 155848
rect 209740 155808 258074 155836
rect 209740 155796 209746 155808
rect 200390 155768 200396 155780
rect 191208 155740 196756 155768
rect 196820 155740 200396 155768
rect 196820 155700 196848 155740
rect 200390 155728 200396 155740
rect 200448 155728 200454 155780
rect 200574 155728 200580 155780
rect 200632 155768 200638 155780
rect 240410 155768 240416 155780
rect 200632 155740 240416 155768
rect 200632 155728 200638 155740
rect 240410 155728 240416 155740
rect 240468 155728 240474 155780
rect 240502 155728 240508 155780
rect 240560 155768 240566 155780
rect 240560 155740 244688 155768
rect 240560 155728 240566 155740
rect 177500 155672 196848 155700
rect 196894 155660 196900 155712
rect 196952 155700 196958 155712
rect 200206 155700 200212 155712
rect 196952 155672 200212 155700
rect 196952 155660 196958 155672
rect 200206 155660 200212 155672
rect 200264 155660 200270 155712
rect 200298 155660 200304 155712
rect 200356 155700 200362 155712
rect 244550 155700 244556 155712
rect 200356 155672 244556 155700
rect 200356 155660 200362 155672
rect 244550 155660 244556 155672
rect 244608 155660 244614 155712
rect 222746 155632 222752 155644
rect 166966 155604 222752 155632
rect 153344 155592 153350 155604
rect 222746 155592 222752 155604
rect 222804 155592 222810 155644
rect 222838 155592 222844 155644
rect 222896 155632 222902 155644
rect 223482 155632 223488 155644
rect 222896 155604 223488 155632
rect 222896 155592 222902 155604
rect 223482 155592 223488 155604
rect 223540 155592 223546 155644
rect 223574 155592 223580 155644
rect 223632 155632 223638 155644
rect 228450 155632 228456 155644
rect 223632 155604 228456 155632
rect 223632 155592 223638 155604
rect 228450 155592 228456 155604
rect 228508 155592 228514 155644
rect 230382 155592 230388 155644
rect 230440 155632 230446 155644
rect 233970 155632 233976 155644
rect 230440 155604 233976 155632
rect 230440 155592 230446 155604
rect 233970 155592 233976 155604
rect 234028 155592 234034 155644
rect 234614 155592 234620 155644
rect 234672 155632 234678 155644
rect 243538 155632 243544 155644
rect 234672 155604 243544 155632
rect 234672 155592 234678 155604
rect 243538 155592 243544 155604
rect 243596 155592 243602 155644
rect 244660 155632 244688 155740
rect 244826 155728 244832 155780
rect 244884 155768 244890 155780
rect 248138 155768 248144 155780
rect 244884 155740 248144 155768
rect 244884 155728 244890 155740
rect 248138 155728 248144 155740
rect 248196 155728 248202 155780
rect 249058 155728 249064 155780
rect 249116 155768 249122 155780
rect 257246 155768 257252 155780
rect 249116 155740 257252 155768
rect 249116 155728 249122 155740
rect 257246 155728 257252 155740
rect 257304 155728 257310 155780
rect 258046 155768 258074 155808
rect 259822 155796 259828 155848
rect 259880 155836 259886 155848
rect 277366 155836 277394 155876
rect 281626 155864 281632 155916
rect 281684 155904 281690 155916
rect 299428 155904 299434 155916
rect 281684 155876 299434 155904
rect 281684 155864 281690 155876
rect 299428 155864 299434 155876
rect 299486 155864 299492 155916
rect 299566 155864 299572 155916
rect 299624 155904 299630 155916
rect 326154 155904 326160 155916
rect 299624 155876 326160 155904
rect 299624 155864 299630 155876
rect 326154 155864 326160 155876
rect 326212 155864 326218 155916
rect 328426 155904 328454 156012
rect 333606 156000 333612 156012
rect 333664 156000 333670 156052
rect 335998 156000 336004 156052
rect 336056 156040 336062 156052
rect 336056 156012 336412 156040
rect 336056 156000 336062 156012
rect 326264 155876 328454 155904
rect 331784 155944 335400 155972
rect 259880 155808 277394 155836
rect 259880 155796 259886 155808
rect 277486 155796 277492 155848
rect 277544 155836 277550 155848
rect 282454 155836 282460 155848
rect 277544 155808 282460 155836
rect 277544 155796 277550 155808
rect 282454 155796 282460 155808
rect 282512 155796 282518 155848
rect 283282 155796 283288 155848
rect 283340 155836 283346 155848
rect 287330 155836 287336 155848
rect 283340 155808 287336 155836
rect 283340 155796 283346 155808
rect 287330 155796 287336 155808
rect 287388 155796 287394 155848
rect 287514 155796 287520 155848
rect 287572 155836 287578 155848
rect 295702 155836 295708 155848
rect 287572 155808 295708 155836
rect 287572 155796 287578 155808
rect 295702 155796 295708 155808
rect 295760 155796 295766 155848
rect 295794 155796 295800 155848
rect 295852 155836 295858 155848
rect 326264 155836 326292 155876
rect 295852 155808 326292 155836
rect 295852 155796 295858 155808
rect 326430 155796 326436 155848
rect 326488 155836 326494 155848
rect 331784 155836 331812 155944
rect 335262 155904 335268 155916
rect 333716 155876 335268 155904
rect 333716 155836 333744 155876
rect 335262 155864 335268 155876
rect 335320 155864 335326 155916
rect 335372 155904 335400 155944
rect 336384 155904 336412 156012
rect 348878 155932 348884 155984
rect 348936 155972 348942 155984
rect 356514 155972 356520 155984
rect 348936 155944 356520 155972
rect 348936 155932 348942 155944
rect 356514 155932 356520 155944
rect 356572 155932 356578 155984
rect 343910 155904 343916 155916
rect 335372 155876 336320 155904
rect 336384 155876 343916 155904
rect 326488 155808 331812 155836
rect 331876 155808 333744 155836
rect 326488 155796 326494 155808
rect 261386 155768 261392 155780
rect 258046 155740 261392 155768
rect 261386 155728 261392 155740
rect 261444 155728 261450 155780
rect 261478 155728 261484 155780
rect 261536 155768 261542 155780
rect 299474 155768 299480 155780
rect 261536 155740 299480 155768
rect 261536 155728 261542 155740
rect 299474 155728 299480 155740
rect 299532 155728 299538 155780
rect 299566 155728 299572 155780
rect 299624 155768 299630 155780
rect 311618 155768 311624 155780
rect 299624 155740 311624 155768
rect 299624 155728 299630 155740
rect 311618 155728 311624 155740
rect 311676 155728 311682 155780
rect 321370 155768 321376 155780
rect 311866 155740 321376 155768
rect 246298 155660 246304 155712
rect 246356 155700 246362 155712
rect 262122 155700 262128 155712
rect 246356 155672 262128 155700
rect 246356 155660 246362 155672
rect 262122 155660 262128 155672
rect 262180 155660 262186 155712
rect 264054 155660 264060 155712
rect 264112 155700 264118 155712
rect 266722 155700 266728 155712
rect 264112 155672 266728 155700
rect 264112 155660 264118 155672
rect 266722 155660 266728 155672
rect 266780 155660 266786 155712
rect 268194 155660 268200 155712
rect 268252 155700 268258 155712
rect 311866 155700 311894 155740
rect 321370 155728 321376 155740
rect 321428 155728 321434 155780
rect 321462 155728 321468 155780
rect 321520 155768 321526 155780
rect 331766 155768 331772 155780
rect 321520 155740 331772 155768
rect 321520 155728 321526 155740
rect 331766 155728 331772 155740
rect 331824 155728 331830 155780
rect 268252 155672 311894 155700
rect 268252 155660 268258 155672
rect 312078 155660 312084 155712
rect 312136 155700 312142 155712
rect 315942 155700 315948 155712
rect 312136 155672 315948 155700
rect 312136 155660 312142 155672
rect 315942 155660 315948 155672
rect 316000 155660 316006 155712
rect 316586 155660 316592 155712
rect 316644 155700 316650 155712
rect 320174 155700 320180 155712
rect 316644 155672 320180 155700
rect 316644 155660 316650 155672
rect 320174 155660 320180 155672
rect 320232 155660 320238 155712
rect 320266 155660 320272 155712
rect 320324 155700 320330 155712
rect 326338 155700 326344 155712
rect 320324 155672 326344 155700
rect 320324 155660 320330 155672
rect 326338 155660 326344 155672
rect 326396 155660 326402 155712
rect 326522 155660 326528 155712
rect 326580 155700 326586 155712
rect 331876 155700 331904 155808
rect 333790 155796 333796 155848
rect 333848 155836 333854 155848
rect 336182 155836 336188 155848
rect 333848 155808 336188 155836
rect 333848 155796 333854 155808
rect 336182 155796 336188 155808
rect 336240 155796 336246 155848
rect 336292 155836 336320 155876
rect 343910 155864 343916 155876
rect 343968 155864 343974 155916
rect 344646 155864 344652 155916
rect 344704 155904 344710 155916
rect 382366 155904 382372 155916
rect 344704 155876 382372 155904
rect 344704 155864 344710 155876
rect 382366 155864 382372 155876
rect 382424 155864 382430 155916
rect 402238 155904 402244 155916
rect 398944 155876 402244 155904
rect 337838 155836 337844 155848
rect 336292 155808 337844 155836
rect 337838 155796 337844 155808
rect 337896 155796 337902 155848
rect 337930 155796 337936 155848
rect 337988 155836 337994 155848
rect 340782 155836 340788 155848
rect 337988 155808 340788 155836
rect 337988 155796 337994 155808
rect 340782 155796 340788 155808
rect 340840 155796 340846 155848
rect 342162 155796 342168 155848
rect 342220 155836 342226 155848
rect 380526 155836 380532 155848
rect 342220 155808 380532 155836
rect 342220 155796 342226 155808
rect 380526 155796 380532 155808
rect 380584 155796 380590 155848
rect 381630 155796 381636 155848
rect 381688 155836 381694 155848
rect 398834 155836 398840 155848
rect 381688 155808 398840 155836
rect 381688 155796 381694 155808
rect 398834 155796 398840 155808
rect 398892 155796 398898 155848
rect 331950 155728 331956 155780
rect 332008 155768 332014 155780
rect 351270 155768 351276 155780
rect 332008 155740 351276 155768
rect 332008 155728 332014 155740
rect 351270 155728 351276 155740
rect 351328 155728 351334 155780
rect 355226 155728 355232 155780
rect 355284 155768 355290 155780
rect 357986 155768 357992 155780
rect 355284 155740 357992 155768
rect 355284 155728 355290 155740
rect 357986 155728 357992 155740
rect 358044 155728 358050 155780
rect 358078 155728 358084 155780
rect 358136 155768 358142 155780
rect 364702 155768 364708 155780
rect 358136 155740 364708 155768
rect 358136 155728 358142 155740
rect 364702 155728 364708 155740
rect 364760 155728 364766 155780
rect 364794 155728 364800 155780
rect 364852 155768 364858 155780
rect 384574 155768 384580 155780
rect 364852 155740 384580 155768
rect 364852 155728 364858 155740
rect 384574 155728 384580 155740
rect 384632 155728 384638 155780
rect 388346 155728 388352 155780
rect 388404 155768 388410 155780
rect 398944 155768 398972 155876
rect 402238 155864 402244 155876
rect 402296 155864 402302 155916
rect 411806 155864 411812 155916
rect 411864 155904 411870 155916
rect 413922 155904 413928 155916
rect 411864 155876 413928 155904
rect 411864 155864 411870 155876
rect 413922 155864 413928 155876
rect 413980 155864 413986 155916
rect 443730 155864 443736 155916
rect 443788 155904 443794 155916
rect 458266 155904 458272 155916
rect 443788 155876 458272 155904
rect 443788 155864 443794 155876
rect 458266 155864 458272 155876
rect 458324 155864 458330 155916
rect 460566 155864 460572 155916
rect 460624 155904 460630 155916
rect 470502 155904 470508 155916
rect 460624 155876 470508 155904
rect 460624 155864 460630 155876
rect 470502 155864 470508 155876
rect 470560 155864 470566 155916
rect 471422 155864 471428 155916
rect 471480 155904 471486 155916
rect 476114 155904 476120 155916
rect 471480 155876 476120 155904
rect 471480 155864 471486 155876
rect 476114 155864 476120 155876
rect 476172 155864 476178 155916
rect 476482 155864 476488 155916
rect 476540 155904 476546 155916
rect 482922 155904 482928 155916
rect 476540 155876 482928 155904
rect 476540 155864 476546 155876
rect 482922 155864 482928 155876
rect 482980 155864 482986 155916
rect 488258 155864 488264 155916
rect 488316 155904 488322 155916
rect 490374 155904 490380 155916
rect 488316 155876 490380 155904
rect 488316 155864 488322 155876
rect 490374 155864 490380 155876
rect 490432 155864 490438 155916
rect 499206 155864 499212 155916
rect 499264 155904 499270 155916
rect 500586 155904 500592 155916
rect 499264 155876 500592 155904
rect 499264 155864 499270 155876
rect 500586 155864 500592 155876
rect 500644 155864 500650 155916
rect 509050 155864 509056 155916
rect 509108 155904 509114 155916
rect 510062 155904 510068 155916
rect 509108 155876 510068 155904
rect 509108 155864 509114 155876
rect 510062 155864 510068 155876
rect 510120 155864 510126 155916
rect 516042 155864 516048 155916
rect 516100 155904 516106 155916
rect 519354 155904 519360 155916
rect 516100 155876 519360 155904
rect 516100 155864 516106 155876
rect 519354 155864 519360 155876
rect 519412 155864 519418 155916
rect 401778 155796 401784 155848
rect 401836 155836 401842 155848
rect 407298 155836 407304 155848
rect 401836 155808 407304 155836
rect 401836 155796 401842 155808
rect 407298 155796 407304 155808
rect 407356 155796 407362 155848
rect 419350 155796 419356 155848
rect 419408 155836 419414 155848
rect 423214 155836 423220 155848
rect 419408 155808 423220 155836
rect 419408 155796 419414 155808
rect 423214 155796 423220 155808
rect 423272 155796 423278 155848
rect 442074 155796 442080 155848
rect 442132 155836 442138 155848
rect 456978 155836 456984 155848
rect 442132 155808 456984 155836
rect 442132 155796 442138 155808
rect 456978 155796 456984 155808
rect 457036 155796 457042 155848
rect 458910 155796 458916 155848
rect 458968 155836 458974 155848
rect 458968 155808 465672 155836
rect 458968 155796 458974 155808
rect 388404 155740 398972 155768
rect 388404 155728 388410 155740
rect 399202 155728 399208 155780
rect 399260 155768 399266 155780
rect 416682 155768 416688 155780
rect 399260 155740 416688 155768
rect 399260 155728 399266 155740
rect 416682 155728 416688 155740
rect 416740 155728 416746 155780
rect 424410 155728 424416 155780
rect 424468 155768 424474 155780
rect 437474 155768 437480 155780
rect 424468 155740 437480 155768
rect 424468 155728 424474 155740
rect 437474 155728 437480 155740
rect 437532 155728 437538 155780
rect 439590 155728 439596 155780
rect 439648 155768 439654 155780
rect 455046 155768 455052 155780
rect 439648 155740 455052 155768
rect 439648 155728 439654 155740
rect 455046 155728 455052 155740
rect 455104 155728 455110 155780
rect 456334 155728 456340 155780
rect 456392 155768 456398 155780
rect 464338 155768 464344 155780
rect 456392 155740 464344 155768
rect 456392 155728 456398 155740
rect 464338 155728 464344 155740
rect 464396 155728 464402 155780
rect 326580 155672 331904 155700
rect 326580 155660 326586 155672
rect 332042 155660 332048 155712
rect 332100 155700 332106 155712
rect 333974 155700 333980 155712
rect 332100 155672 333980 155700
rect 332100 155660 332106 155672
rect 333974 155660 333980 155672
rect 334032 155660 334038 155712
rect 335446 155660 335452 155712
rect 335504 155700 335510 155712
rect 365346 155700 365352 155712
rect 335504 155672 351316 155700
rect 335504 155660 335510 155672
rect 292574 155632 292580 155644
rect 244660 155604 292580 155632
rect 292574 155592 292580 155604
rect 292632 155592 292638 155644
rect 295886 155592 295892 155644
rect 295944 155632 295950 155644
rect 299658 155632 299664 155644
rect 295944 155604 299664 155632
rect 295944 155592 295950 155604
rect 299658 155592 299664 155604
rect 299716 155592 299722 155644
rect 300118 155592 300124 155644
rect 300176 155632 300182 155644
rect 302786 155632 302792 155644
rect 300176 155604 302792 155632
rect 300176 155592 300182 155604
rect 302786 155592 302792 155604
rect 302844 155592 302850 155644
rect 302878 155592 302884 155644
rect 302936 155632 302942 155644
rect 340966 155632 340972 155644
rect 302936 155604 340972 155632
rect 302936 155592 302942 155604
rect 340966 155592 340972 155604
rect 341024 155592 341030 155644
rect 341058 155592 341064 155644
rect 341116 155632 341122 155644
rect 349890 155632 349896 155644
rect 341116 155604 349896 155632
rect 341116 155592 341122 155604
rect 349890 155592 349896 155604
rect 349948 155592 349954 155644
rect 351288 155632 351316 155672
rect 351472 155672 365352 155700
rect 351472 155632 351500 155672
rect 365346 155660 365352 155672
rect 365404 155660 365410 155712
rect 382458 155660 382464 155712
rect 382516 155700 382522 155712
rect 382516 155672 405044 155700
rect 382516 155660 382522 155672
rect 351288 155604 351500 155632
rect 356514 155592 356520 155644
rect 356572 155632 356578 155644
rect 365070 155632 365076 155644
rect 356572 155604 365076 155632
rect 356572 155592 356578 155604
rect 365070 155592 365076 155604
rect 365128 155592 365134 155644
rect 365254 155592 365260 155644
rect 365312 155632 365318 155644
rect 385586 155632 385592 155644
rect 365312 155604 385592 155632
rect 365312 155592 365318 155604
rect 385586 155592 385592 155604
rect 385644 155592 385650 155644
rect 398374 155592 398380 155644
rect 398432 155632 398438 155644
rect 404906 155632 404912 155644
rect 398432 155604 404912 155632
rect 398432 155592 398438 155604
rect 404906 155592 404912 155604
rect 404964 155592 404970 155644
rect 405016 155632 405044 155672
rect 405090 155660 405096 155712
rect 405148 155700 405154 155712
rect 408862 155700 408868 155712
rect 405148 155672 408868 155700
rect 405148 155660 405154 155672
rect 408862 155660 408868 155672
rect 408920 155660 408926 155712
rect 433702 155660 433708 155712
rect 433760 155700 433766 155712
rect 448606 155700 448612 155712
rect 433760 155672 448612 155700
rect 433760 155660 433766 155672
rect 448606 155660 448612 155672
rect 448664 155660 448670 155712
rect 452838 155700 452844 155712
rect 451246 155672 452844 155700
rect 411346 155632 411352 155644
rect 405016 155604 411352 155632
rect 411346 155592 411352 155604
rect 411404 155592 411410 155644
rect 412634 155592 412640 155644
rect 412692 155632 412698 155644
rect 420178 155632 420184 155644
rect 412692 155604 420184 155632
rect 412692 155592 412698 155604
rect 420178 155592 420184 155604
rect 420236 155592 420242 155644
rect 435358 155592 435364 155644
rect 435416 155632 435422 155644
rect 435416 155604 445340 155632
rect 435416 155592 435422 155604
rect 59998 155524 60004 155576
rect 60056 155564 60062 155576
rect 153654 155564 153660 155576
rect 60056 155536 153660 155564
rect 60056 155524 60062 155536
rect 153654 155524 153660 155536
rect 153712 155524 153718 155576
rect 154850 155524 154856 155576
rect 154908 155564 154914 155576
rect 155678 155564 155684 155576
rect 154908 155536 155684 155564
rect 154908 155524 154914 155536
rect 155678 155524 155684 155536
rect 155736 155524 155742 155576
rect 156506 155524 156512 155576
rect 156564 155564 156570 155576
rect 158806 155564 158812 155576
rect 156564 155536 158812 155564
rect 156564 155524 156570 155536
rect 158806 155524 158812 155536
rect 158864 155524 158870 155576
rect 159910 155524 159916 155576
rect 159968 155564 159974 155576
rect 164326 155564 164332 155576
rect 159968 155536 164332 155564
rect 159968 155524 159974 155536
rect 164326 155524 164332 155536
rect 164384 155524 164390 155576
rect 164418 155524 164424 155576
rect 164476 155564 164482 155576
rect 169754 155564 169760 155576
rect 164476 155536 169760 155564
rect 164476 155524 164482 155536
rect 169754 155524 169760 155536
rect 169812 155524 169818 155576
rect 170858 155524 170864 155576
rect 170916 155564 170922 155576
rect 173250 155564 173256 155576
rect 170916 155536 173256 155564
rect 170916 155524 170922 155536
rect 173250 155524 173256 155536
rect 173308 155524 173314 155576
rect 173342 155524 173348 155576
rect 173400 155564 173406 155576
rect 180058 155564 180064 155576
rect 173400 155536 180064 155564
rect 173400 155524 173406 155536
rect 180058 155524 180064 155536
rect 180116 155524 180122 155576
rect 180886 155524 180892 155576
rect 180944 155564 180950 155576
rect 185670 155564 185676 155576
rect 180944 155536 185676 155564
rect 180944 155524 180950 155536
rect 185670 155524 185676 155536
rect 185728 155524 185734 155576
rect 232314 155564 232320 155576
rect 186286 155536 232320 155564
rect 70026 155456 70032 155508
rect 70084 155496 70090 155508
rect 162118 155496 162124 155508
rect 70084 155468 162124 155496
rect 70084 155456 70090 155468
rect 162118 155456 162124 155468
rect 162176 155456 162182 155508
rect 164142 155456 164148 155508
rect 164200 155496 164206 155508
rect 165614 155496 165620 155508
rect 164200 155468 165620 155496
rect 164200 155456 164206 155468
rect 165614 155456 165620 155468
rect 165672 155456 165678 155508
rect 166626 155456 166632 155508
rect 166684 155496 166690 155508
rect 186286 155496 186314 155536
rect 232314 155524 232320 155536
rect 232372 155524 232378 155576
rect 232498 155524 232504 155576
rect 232556 155564 232562 155576
rect 233142 155564 233148 155576
rect 232556 155536 233148 155564
rect 232556 155524 232562 155536
rect 233142 155524 233148 155536
rect 233200 155524 233206 155576
rect 233878 155524 233884 155576
rect 233936 155564 233942 155576
rect 272518 155564 272524 155576
rect 233936 155536 272524 155564
rect 233936 155524 233942 155536
rect 272518 155524 272524 155536
rect 272576 155524 272582 155576
rect 272702 155524 272708 155576
rect 272760 155564 272766 155576
rect 299566 155564 299572 155576
rect 272760 155536 299572 155564
rect 272760 155524 272766 155536
rect 299566 155524 299572 155536
rect 299624 155524 299630 155576
rect 306834 155524 306840 155576
rect 306892 155564 306898 155576
rect 325418 155564 325424 155576
rect 306892 155536 325424 155564
rect 306892 155524 306898 155536
rect 325418 155524 325424 155536
rect 325476 155524 325482 155576
rect 326614 155524 326620 155576
rect 326672 155564 326678 155576
rect 328638 155564 328644 155576
rect 326672 155536 328644 155564
rect 326672 155524 326678 155536
rect 328638 155524 328644 155536
rect 328696 155524 328702 155576
rect 328730 155524 328736 155576
rect 328788 155564 328794 155576
rect 336090 155564 336096 155576
rect 328788 155536 336096 155564
rect 328788 155524 328794 155536
rect 336090 155524 336096 155536
rect 336148 155524 336154 155576
rect 336182 155524 336188 155576
rect 336240 155564 336246 155576
rect 364978 155564 364984 155576
rect 336240 155536 364984 155564
rect 336240 155524 336246 155536
rect 364978 155524 364984 155536
rect 365036 155524 365042 155576
rect 365346 155524 365352 155576
rect 365404 155564 365410 155576
rect 375466 155564 375472 155576
rect 365404 155536 375472 155564
rect 365404 155524 365410 155536
rect 375466 155524 375472 155536
rect 375524 155524 375530 155576
rect 379054 155524 379060 155576
rect 379112 155564 379118 155576
rect 408770 155564 408776 155576
rect 379112 155536 408776 155564
rect 379112 155524 379118 155536
rect 408770 155524 408776 155536
rect 408828 155524 408834 155576
rect 410150 155524 410156 155576
rect 410208 155564 410214 155576
rect 417418 155564 417424 155576
rect 410208 155536 417424 155564
rect 410208 155524 410214 155536
rect 417418 155524 417424 155536
rect 417476 155524 417482 155576
rect 421098 155524 421104 155576
rect 421156 155564 421162 155576
rect 430574 155564 430580 155576
rect 421156 155536 430580 155564
rect 421156 155524 421162 155536
rect 430574 155524 430580 155536
rect 430632 155524 430638 155576
rect 431954 155524 431960 155576
rect 432012 155564 432018 155576
rect 445202 155564 445208 155576
rect 432012 155536 445208 155564
rect 432012 155524 432018 155536
rect 445202 155524 445208 155536
rect 445260 155524 445266 155576
rect 445312 155564 445340 155604
rect 446398 155592 446404 155644
rect 446456 155632 446462 155644
rect 451246 155632 451274 155672
rect 452838 155660 452844 155672
rect 452896 155660 452902 155712
rect 453850 155660 453856 155712
rect 453908 155700 453914 155712
rect 465534 155700 465540 155712
rect 453908 155672 465540 155700
rect 453908 155660 453914 155672
rect 465534 155660 465540 155672
rect 465592 155660 465598 155712
rect 465644 155700 465672 155808
rect 466454 155796 466460 155848
rect 466512 155836 466518 155848
rect 473078 155836 473084 155848
rect 466512 155808 473084 155836
rect 466512 155796 466518 155808
rect 473078 155796 473084 155808
rect 473136 155796 473142 155848
rect 480714 155796 480720 155848
rect 480772 155836 480778 155848
rect 486326 155836 486332 155848
rect 480772 155808 486332 155836
rect 480772 155796 480778 155808
rect 486326 155796 486332 155808
rect 486384 155796 486390 155848
rect 498378 155796 498384 155848
rect 498436 155836 498442 155848
rect 499574 155836 499580 155848
rect 498436 155808 499580 155836
rect 498436 155796 498442 155808
rect 499574 155796 499580 155808
rect 499632 155796 499638 155848
rect 469306 155768 469312 155780
rect 467852 155740 469312 155768
rect 467852 155700 467880 155740
rect 469306 155728 469312 155740
rect 469364 155728 469370 155780
rect 469766 155728 469772 155780
rect 469824 155768 469830 155780
rect 474734 155768 474740 155780
rect 469824 155740 474740 155768
rect 469824 155728 469830 155740
rect 474734 155728 474740 155740
rect 474792 155728 474798 155780
rect 479058 155728 479064 155780
rect 479116 155768 479122 155780
rect 484946 155768 484952 155780
rect 479116 155740 484952 155768
rect 479116 155728 479122 155740
rect 484946 155728 484952 155740
rect 485004 155728 485010 155780
rect 517330 155728 517336 155780
rect 517388 155768 517394 155780
rect 521010 155768 521016 155780
rect 517388 155740 521016 155768
rect 517388 155728 517394 155740
rect 521010 155728 521016 155740
rect 521068 155728 521074 155780
rect 465644 155672 467880 155700
rect 468110 155660 468116 155712
rect 468168 155700 468174 155712
rect 473630 155700 473636 155712
rect 468168 155672 473636 155700
rect 468168 155660 468174 155672
rect 473630 155660 473636 155672
rect 473688 155660 473694 155712
rect 475654 155660 475660 155712
rect 475712 155700 475718 155712
rect 480714 155700 480720 155712
rect 475712 155672 480720 155700
rect 475712 155660 475718 155672
rect 480714 155660 480720 155672
rect 480772 155660 480778 155712
rect 492490 155660 492496 155712
rect 492548 155700 492554 155712
rect 495342 155700 495348 155712
rect 492548 155672 495348 155700
rect 492548 155660 492554 155672
rect 495342 155660 495348 155672
rect 495400 155660 495406 155712
rect 515490 155660 515496 155712
rect 515548 155700 515554 155712
rect 518526 155700 518532 155712
rect 515548 155672 518532 155700
rect 515548 155660 515554 155672
rect 518526 155660 518532 155672
rect 518584 155660 518590 155712
rect 446456 155604 451274 155632
rect 446456 155592 446462 155604
rect 452102 155592 452108 155644
rect 452160 155632 452166 155644
rect 452160 155604 462820 155632
rect 452160 155592 452166 155604
rect 445312 155536 446628 155564
rect 166684 155468 186314 155496
rect 166684 155456 166690 155468
rect 186774 155456 186780 155508
rect 186832 155496 186838 155508
rect 191006 155496 191012 155508
rect 186832 155468 191012 155496
rect 186832 155456 186838 155468
rect 191006 155456 191012 155468
rect 191064 155456 191070 155508
rect 191098 155456 191104 155508
rect 191156 155496 191162 155508
rect 249058 155496 249064 155508
rect 191156 155468 249064 155496
rect 191156 155456 191162 155468
rect 249058 155456 249064 155468
rect 249116 155456 249122 155508
rect 249150 155456 249156 155508
rect 249208 155496 249214 155508
rect 254118 155496 254124 155508
rect 249208 155468 254124 155496
rect 249208 155456 249214 155468
rect 254118 155456 254124 155468
rect 254176 155456 254182 155508
rect 257338 155456 257344 155508
rect 257396 155496 257402 155508
rect 260558 155496 260564 155508
rect 257396 155468 260564 155496
rect 257396 155456 257402 155468
rect 260558 155456 260564 155468
rect 260616 155456 260622 155508
rect 260650 155456 260656 155508
rect 260708 155496 260714 155508
rect 311710 155496 311716 155508
rect 260708 155468 311716 155496
rect 260708 155456 260714 155468
rect 311710 155456 311716 155468
rect 311768 155456 311774 155508
rect 311802 155456 311808 155508
rect 311860 155496 311866 155508
rect 314562 155496 314568 155508
rect 311860 155468 314568 155496
rect 311860 155456 311866 155468
rect 314562 155456 314568 155468
rect 314620 155456 314626 155508
rect 315298 155456 315304 155508
rect 315356 155496 315362 155508
rect 321370 155496 321376 155508
rect 315356 155468 321376 155496
rect 315356 155456 315362 155468
rect 321370 155456 321376 155468
rect 321428 155456 321434 155508
rect 321462 155456 321468 155508
rect 321520 155496 321526 155508
rect 321520 155468 322428 155496
rect 321520 155456 321526 155468
rect 10410 155388 10416 155440
rect 10468 155428 10474 155440
rect 107746 155428 107752 155440
rect 10468 155400 107752 155428
rect 10468 155388 10474 155400
rect 107746 155388 107752 155400
rect 107804 155388 107810 155440
rect 107838 155388 107844 155440
rect 107896 155428 107902 155440
rect 108942 155428 108948 155440
rect 107896 155400 108948 155428
rect 107896 155388 107902 155400
rect 108942 155388 108948 155400
rect 109000 155388 109006 155440
rect 109034 155388 109040 155440
rect 109092 155428 109098 155440
rect 110138 155428 110144 155440
rect 109092 155400 110144 155428
rect 109092 155388 109098 155400
rect 110138 155388 110144 155400
rect 110196 155388 110202 155440
rect 111150 155388 111156 155440
rect 111208 155428 111214 155440
rect 111702 155428 111708 155440
rect 111208 155400 111708 155428
rect 111208 155388 111214 155400
rect 111702 155388 111708 155400
rect 111760 155388 111766 155440
rect 115382 155388 115388 155440
rect 115440 155428 115446 155440
rect 115842 155428 115848 155440
rect 115440 155400 115848 155428
rect 115440 155388 115446 155400
rect 115842 155388 115848 155400
rect 115900 155388 115906 155440
rect 116210 155388 116216 155440
rect 116268 155428 116274 155440
rect 117222 155428 117228 155440
rect 116268 155400 117228 155428
rect 116268 155388 116274 155400
rect 117222 155388 117228 155400
rect 117280 155388 117286 155440
rect 117866 155388 117872 155440
rect 117924 155428 117930 155440
rect 118602 155428 118608 155440
rect 117924 155400 118608 155428
rect 117924 155388 117930 155400
rect 118602 155388 118608 155400
rect 118660 155388 118666 155440
rect 120534 155388 120540 155440
rect 120592 155428 120598 155440
rect 122742 155428 122748 155440
rect 120592 155400 122748 155428
rect 120592 155388 120598 155400
rect 122742 155388 122748 155400
rect 122800 155388 122806 155440
rect 123478 155388 123484 155440
rect 123536 155428 123542 155440
rect 200758 155428 200764 155440
rect 123536 155400 200764 155428
rect 123536 155388 123542 155400
rect 200758 155388 200764 155400
rect 200816 155388 200822 155440
rect 200850 155388 200856 155440
rect 200908 155428 200914 155440
rect 209682 155428 209688 155440
rect 200908 155400 209688 155428
rect 200908 155388 200914 155400
rect 209682 155388 209688 155400
rect 209740 155388 209746 155440
rect 209774 155388 209780 155440
rect 209832 155428 209838 155440
rect 262858 155428 262864 155440
rect 209832 155400 262864 155428
rect 209832 155388 209838 155400
rect 262858 155388 262864 155400
rect 262916 155388 262922 155440
rect 264882 155388 264888 155440
rect 264940 155428 264946 155440
rect 266446 155428 266452 155440
rect 264940 155400 266452 155428
rect 264940 155388 264946 155400
rect 266446 155388 266452 155400
rect 266504 155388 266510 155440
rect 267366 155388 267372 155440
rect 267424 155428 267430 155440
rect 272518 155428 272524 155440
rect 267424 155400 272524 155428
rect 267424 155388 267430 155400
rect 272518 155388 272524 155400
rect 272576 155388 272582 155440
rect 272794 155388 272800 155440
rect 272852 155428 272858 155440
rect 273990 155428 273996 155440
rect 272852 155400 273996 155428
rect 272852 155388 272858 155400
rect 273990 155388 273996 155400
rect 274048 155388 274054 155440
rect 274082 155388 274088 155440
rect 274140 155428 274146 155440
rect 299658 155428 299664 155440
rect 274140 155400 299664 155428
rect 274140 155388 274146 155400
rect 299658 155388 299664 155400
rect 299716 155388 299722 155440
rect 299750 155388 299756 155440
rect 299808 155428 299814 155440
rect 316678 155428 316684 155440
rect 299808 155400 316684 155428
rect 299808 155388 299814 155400
rect 316678 155388 316684 155400
rect 316736 155388 316742 155440
rect 316770 155388 316776 155440
rect 316828 155428 316834 155440
rect 320266 155428 320272 155440
rect 316828 155400 320272 155428
rect 316828 155388 316834 155400
rect 320266 155388 320272 155400
rect 320324 155388 320330 155440
rect 322400 155428 322428 155468
rect 327258 155456 327264 155508
rect 327316 155496 327322 155508
rect 351638 155496 351644 155508
rect 327316 155468 351644 155496
rect 327316 155456 327322 155468
rect 351638 155456 351644 155468
rect 351696 155456 351702 155508
rect 351730 155456 351736 155508
rect 351788 155496 351794 155508
rect 355226 155496 355232 155508
rect 351788 155468 355232 155496
rect 351788 155456 351794 155468
rect 355226 155456 355232 155468
rect 355284 155456 355290 155508
rect 355318 155456 355324 155508
rect 355376 155496 355382 155508
rect 362678 155496 362684 155508
rect 355376 155468 362684 155496
rect 355376 155456 355382 155468
rect 362678 155456 362684 155468
rect 362736 155456 362742 155508
rect 369026 155456 369032 155508
rect 369084 155496 369090 155508
rect 401042 155496 401048 155508
rect 369084 155468 401048 155496
rect 369084 155456 369090 155468
rect 401042 155456 401048 155468
rect 401100 155456 401106 155508
rect 405918 155456 405924 155508
rect 405976 155496 405982 155508
rect 419166 155496 419172 155508
rect 405976 155468 419172 155496
rect 405976 155456 405982 155468
rect 419166 155456 419172 155468
rect 419224 155456 419230 155508
rect 426986 155456 426992 155508
rect 427044 155496 427050 155508
rect 445110 155496 445116 155508
rect 427044 155468 445116 155496
rect 427044 155456 427050 155468
rect 445110 155456 445116 155468
rect 445168 155456 445174 155508
rect 325234 155428 325240 155440
rect 322400 155400 325240 155428
rect 325234 155388 325240 155400
rect 325292 155388 325298 155440
rect 325418 155388 325424 155440
rect 325476 155428 325482 155440
rect 331214 155428 331220 155440
rect 325476 155400 331220 155428
rect 325476 155388 325482 155400
rect 331214 155388 331220 155400
rect 331272 155388 331278 155440
rect 331306 155388 331312 155440
rect 331364 155428 331370 155440
rect 335906 155428 335912 155440
rect 331364 155400 335912 155428
rect 331364 155388 331370 155400
rect 335906 155388 335912 155400
rect 335964 155388 335970 155440
rect 336090 155388 336096 155440
rect 336148 155428 336154 155440
rect 370222 155428 370228 155440
rect 336148 155400 370228 155428
rect 336148 155388 336154 155400
rect 370222 155388 370228 155400
rect 370280 155388 370286 155440
rect 375742 155388 375748 155440
rect 375800 155428 375806 155440
rect 406194 155428 406200 155440
rect 375800 155400 406200 155428
rect 375800 155388 375806 155400
rect 406194 155388 406200 155400
rect 406252 155388 406258 155440
rect 413554 155388 413560 155440
rect 413612 155428 413618 155440
rect 435082 155428 435088 155440
rect 413612 155400 435088 155428
rect 413612 155388 413618 155400
rect 435082 155388 435088 155400
rect 435140 155388 435146 155440
rect 438670 155388 438676 155440
rect 438728 155428 438734 155440
rect 446398 155428 446404 155440
rect 438728 155400 446404 155428
rect 438728 155388 438734 155400
rect 446398 155388 446404 155400
rect 446456 155388 446462 155440
rect 446600 155428 446628 155536
rect 449618 155524 449624 155576
rect 449676 155564 449682 155576
rect 462682 155564 462688 155576
rect 449676 155536 462688 155564
rect 449676 155524 449682 155536
rect 462682 155524 462688 155536
rect 462740 155524 462746 155576
rect 462792 155564 462820 155604
rect 463878 155592 463884 155644
rect 463936 155632 463942 155644
rect 473354 155632 473360 155644
rect 463936 155604 473360 155632
rect 463936 155592 463942 155604
rect 473354 155592 473360 155604
rect 473412 155592 473418 155644
rect 474826 155592 474832 155644
rect 474884 155632 474890 155644
rect 480806 155632 480812 155644
rect 474884 155604 480812 155632
rect 474884 155592 474890 155604
rect 480806 155592 480812 155604
rect 480864 155592 480870 155644
rect 481542 155592 481548 155644
rect 481600 155632 481606 155644
rect 487062 155632 487068 155644
rect 481600 155604 487068 155632
rect 481600 155592 481606 155604
rect 487062 155592 487068 155604
rect 487120 155592 487126 155644
rect 491662 155592 491668 155644
rect 491720 155632 491726 155644
rect 494606 155632 494612 155644
rect 491720 155604 494612 155632
rect 491720 155592 491726 155604
rect 494606 155592 494612 155604
rect 494664 155592 494670 155644
rect 513558 155592 513564 155644
rect 513616 155632 513622 155644
rect 515950 155632 515956 155644
rect 513616 155604 515956 155632
rect 513616 155592 513622 155604
rect 515950 155592 515956 155604
rect 516008 155592 516014 155644
rect 464614 155564 464620 155576
rect 462792 155536 464620 155564
rect 464614 155524 464620 155536
rect 464672 155524 464678 155576
rect 464706 155524 464712 155576
rect 464764 155564 464770 155576
rect 473906 155564 473912 155576
rect 464764 155536 473912 155564
rect 464764 155524 464770 155536
rect 473906 155524 473912 155536
rect 473964 155524 473970 155576
rect 483198 155524 483204 155576
rect 483256 155564 483262 155576
rect 485866 155564 485872 155576
rect 483256 155536 485872 155564
rect 483256 155524 483262 155536
rect 485866 155524 485872 155536
rect 485924 155524 485930 155576
rect 490742 155524 490748 155576
rect 490800 155564 490806 155576
rect 493962 155564 493968 155576
rect 490800 155536 493968 155564
rect 490800 155524 490806 155536
rect 493962 155524 493968 155536
rect 494020 155524 494026 155576
rect 494146 155524 494152 155576
rect 494204 155564 494210 155576
rect 496722 155564 496728 155576
rect 494204 155536 496728 155564
rect 494204 155524 494210 155536
rect 496722 155524 496728 155536
rect 496780 155524 496786 155576
rect 497458 155524 497464 155576
rect 497516 155564 497522 155576
rect 499298 155564 499304 155576
rect 497516 155536 499304 155564
rect 497516 155524 497522 155536
rect 499298 155524 499304 155536
rect 499356 155524 499362 155576
rect 501690 155524 501696 155576
rect 501748 155564 501754 155576
rect 502426 155564 502432 155576
rect 501748 155536 502432 155564
rect 501748 155524 501754 155536
rect 502426 155524 502432 155536
rect 502484 155524 502490 155576
rect 507762 155524 507768 155576
rect 507820 155564 507826 155576
rect 508406 155564 508412 155576
rect 507820 155536 508412 155564
rect 507820 155524 507826 155536
rect 508406 155524 508412 155536
rect 508464 155524 508470 155576
rect 510522 155524 510528 155576
rect 510580 155564 510586 155576
rect 511810 155564 511816 155576
rect 510580 155536 511816 155564
rect 510580 155524 510586 155536
rect 511810 155524 511816 155536
rect 511868 155524 511874 155576
rect 512270 155524 512276 155576
rect 512328 155564 512334 155576
rect 514294 155564 514300 155576
rect 512328 155536 514300 155564
rect 512328 155524 512334 155536
rect 514294 155524 514300 155536
rect 514352 155524 514358 155576
rect 514846 155524 514852 155576
rect 514904 155564 514910 155576
rect 517606 155564 517612 155576
rect 514904 155536 517612 155564
rect 514904 155524 514910 155536
rect 517606 155524 517612 155536
rect 517664 155524 517670 155576
rect 447962 155456 447968 155508
rect 448020 155496 448026 155508
rect 461394 155496 461400 155508
rect 448020 155468 461400 155496
rect 448020 155456 448026 155468
rect 461394 155456 461400 155468
rect 461452 155456 461458 155508
rect 464338 155456 464344 155508
rect 464396 155496 464402 155508
rect 467742 155496 467748 155508
rect 464396 155468 467748 155496
rect 464396 155456 464402 155468
rect 467742 155456 467748 155468
rect 467800 155456 467806 155508
rect 472342 155456 472348 155508
rect 472400 155496 472406 155508
rect 477586 155496 477592 155508
rect 472400 155468 477592 155496
rect 472400 155456 472406 155468
rect 477586 155456 477592 155468
rect 477644 155456 477650 155508
rect 482370 155456 482376 155508
rect 482428 155496 482434 155508
rect 487706 155496 487712 155508
rect 482428 155468 487712 155496
rect 482428 155456 482434 155468
rect 487706 155456 487712 155468
rect 487764 155456 487770 155508
rect 500034 155456 500040 155508
rect 500092 155496 500098 155508
rect 501230 155496 501236 155508
rect 500092 155468 501236 155496
rect 500092 155456 500098 155468
rect 501230 155456 501236 155468
rect 501288 155456 501294 155508
rect 514202 155456 514208 155508
rect 514260 155496 514266 155508
rect 516778 155496 516784 155508
rect 514260 155468 516784 155496
rect 514260 155456 514266 155468
rect 516778 155456 516784 155468
rect 516836 155456 516842 155508
rect 449986 155428 449992 155440
rect 446600 155400 449992 155428
rect 449986 155388 449992 155400
rect 450044 155388 450050 155440
rect 450446 155388 450452 155440
rect 450504 155428 450510 155440
rect 454586 155428 454592 155440
rect 450504 155400 454592 155428
rect 450504 155388 450510 155400
rect 454586 155388 454592 155400
rect 454644 155388 454650 155440
rect 454678 155388 454684 155440
rect 454736 155428 454742 155440
rect 466362 155428 466368 155440
rect 454736 155400 466368 155428
rect 454736 155388 454742 155400
rect 466362 155388 466368 155400
rect 466420 155388 466426 155440
rect 468938 155388 468944 155440
rect 468996 155428 469002 155440
rect 477494 155428 477500 155440
rect 468996 155400 477500 155428
rect 468996 155388 469002 155400
rect 477494 155388 477500 155400
rect 477552 155388 477558 155440
rect 478138 155388 478144 155440
rect 478196 155428 478202 155440
rect 484302 155428 484308 155440
rect 478196 155400 484308 155428
rect 478196 155388 478202 155400
rect 484302 155388 484308 155400
rect 484360 155388 484366 155440
rect 11238 155320 11244 155372
rect 11296 155360 11302 155372
rect 12342 155360 12348 155372
rect 11296 155332 12348 155360
rect 11296 155320 11302 155332
rect 12342 155320 12348 155332
rect 12400 155320 12406 155372
rect 36446 155320 36452 155372
rect 36504 155360 36510 155372
rect 50338 155360 50344 155372
rect 36504 155332 50344 155360
rect 36504 155320 36510 155332
rect 50338 155320 50344 155332
rect 50396 155320 50402 155372
rect 53282 155320 53288 155372
rect 53340 155360 53346 155372
rect 153930 155360 153936 155372
rect 53340 155332 153936 155360
rect 53340 155320 53346 155332
rect 153930 155320 153936 155332
rect 153988 155320 153994 155372
rect 154022 155320 154028 155372
rect 154080 155360 154086 155372
rect 160646 155360 160652 155372
rect 154080 155332 160652 155360
rect 154080 155320 154086 155332
rect 160646 155320 160652 155332
rect 160704 155320 160710 155372
rect 160738 155320 160744 155372
rect 160796 155360 160802 155372
rect 175918 155360 175924 155372
rect 160796 155332 175924 155360
rect 160796 155320 160802 155332
rect 175918 155320 175924 155332
rect 175976 155320 175982 155372
rect 176010 155320 176016 155372
rect 176068 155360 176074 155372
rect 242894 155360 242900 155372
rect 176068 155332 242900 155360
rect 176068 155320 176074 155332
rect 242894 155320 242900 155332
rect 242952 155320 242958 155372
rect 242986 155320 242992 155372
rect 243044 155360 243050 155372
rect 244642 155360 244648 155372
rect 243044 155332 244648 155360
rect 243044 155320 243050 155332
rect 244642 155320 244648 155332
rect 244700 155320 244706 155372
rect 244734 155320 244740 155372
rect 244792 155360 244798 155372
rect 252554 155360 252560 155372
rect 244792 155332 252560 155360
rect 244792 155320 244798 155332
rect 252554 155320 252560 155332
rect 252612 155320 252618 155372
rect 253934 155320 253940 155372
rect 253992 155360 253998 155372
rect 299566 155360 299572 155372
rect 253992 155332 299572 155360
rect 253992 155320 253998 155332
rect 299566 155320 299572 155332
rect 299624 155320 299630 155372
rect 299842 155320 299848 155372
rect 299900 155360 299906 155372
rect 311894 155360 311900 155372
rect 299900 155332 311900 155360
rect 299900 155320 299906 155332
rect 311894 155320 311900 155332
rect 311952 155320 311958 155372
rect 311986 155320 311992 155372
rect 312044 155360 312050 155372
rect 313182 155360 313188 155372
rect 312044 155332 313188 155360
rect 312044 155320 312050 155332
rect 313182 155320 313188 155332
rect 313240 155320 313246 155372
rect 314378 155320 314384 155372
rect 314436 155360 314442 155372
rect 314436 155332 357434 155360
rect 314436 155320 314442 155332
rect 39850 155252 39856 155304
rect 39908 155292 39914 155304
rect 132954 155292 132960 155304
rect 39908 155264 132960 155292
rect 39908 155252 39914 155264
rect 132954 155252 132960 155264
rect 133012 155252 133018 155304
rect 133046 155252 133052 155304
rect 133104 155292 133110 155304
rect 137002 155292 137008 155304
rect 133104 155264 137008 155292
rect 133104 155252 133110 155264
rect 137002 155252 137008 155264
rect 137060 155252 137066 155304
rect 137370 155252 137376 155304
rect 137428 155292 137434 155304
rect 140774 155292 140780 155304
rect 137428 155264 140780 155292
rect 137428 155252 137434 155264
rect 140774 155252 140780 155264
rect 140832 155252 140838 155304
rect 143074 155252 143080 155304
rect 143132 155292 143138 155304
rect 191006 155292 191012 155304
rect 143132 155264 156736 155292
rect 143132 155252 143138 155264
rect 17954 155184 17960 155236
rect 18012 155224 18018 155236
rect 19242 155224 19248 155236
rect 18012 155196 19248 155224
rect 18012 155184 18018 155196
rect 19242 155184 19248 155196
rect 19300 155184 19306 155236
rect 22186 155184 22192 155236
rect 22244 155224 22250 155236
rect 135898 155224 135904 155236
rect 22244 155196 135904 155224
rect 22244 155184 22250 155196
rect 135898 155184 135904 155196
rect 135956 155184 135962 155236
rect 137186 155184 137192 155236
rect 137244 155224 137250 155236
rect 142614 155224 142620 155236
rect 137244 155196 142620 155224
rect 137244 155184 137250 155196
rect 142614 155184 142620 155196
rect 142672 155184 142678 155236
rect 143902 155184 143908 155236
rect 143960 155224 143966 155236
rect 147582 155224 147588 155236
rect 143960 155196 147588 155224
rect 143960 155184 143966 155196
rect 147582 155184 147588 155196
rect 147640 155184 147646 155236
rect 149790 155184 149796 155236
rect 149848 155224 149854 155236
rect 156598 155224 156604 155236
rect 149848 155196 156604 155224
rect 149848 155184 149854 155196
rect 156598 155184 156604 155196
rect 156656 155184 156662 155236
rect 156708 155224 156736 155264
rect 160756 155264 191012 155292
rect 160756 155224 160784 155264
rect 191006 155252 191012 155264
rect 191064 155252 191070 155304
rect 191098 155252 191104 155304
rect 191156 155292 191162 155304
rect 230382 155292 230388 155304
rect 191156 155264 230388 155292
rect 191156 155252 191162 155264
rect 230382 155252 230388 155264
rect 230440 155252 230446 155304
rect 230474 155252 230480 155304
rect 230532 155292 230538 155304
rect 238662 155292 238668 155304
rect 230532 155264 238668 155292
rect 230532 155252 230538 155264
rect 238662 155252 238668 155264
rect 238720 155252 238726 155304
rect 238754 155252 238760 155304
rect 238812 155292 238818 155304
rect 245470 155292 245476 155304
rect 238812 155264 245476 155292
rect 238812 155252 238818 155264
rect 245470 155252 245476 155264
rect 245528 155252 245534 155304
rect 248046 155252 248052 155304
rect 248104 155292 248110 155304
rect 294046 155292 294052 155304
rect 248104 155264 294052 155292
rect 248104 155252 248110 155264
rect 294046 155252 294052 155264
rect 294104 155252 294110 155304
rect 299474 155292 299480 155304
rect 294156 155264 299480 155292
rect 156708 155196 160784 155224
rect 160830 155184 160836 155236
rect 160888 155224 160894 155236
rect 234614 155224 234620 155236
rect 160888 155196 234620 155224
rect 160888 155184 160894 155196
rect 234614 155184 234620 155196
rect 234672 155184 234678 155236
rect 237190 155184 237196 155236
rect 237248 155224 237254 155236
rect 240502 155224 240508 155236
rect 237248 155196 240508 155224
rect 237248 155184 237254 155196
rect 240502 155184 240508 155196
rect 240560 155184 240566 155236
rect 241330 155184 241336 155236
rect 241388 155224 241394 155236
rect 294156 155224 294184 155264
rect 299474 155252 299480 155264
rect 299532 155252 299538 155304
rect 302786 155252 302792 155304
rect 302844 155292 302850 155304
rect 307110 155292 307116 155304
rect 302844 155264 307116 155292
rect 302844 155252 302850 155264
rect 307110 155252 307116 155264
rect 307168 155252 307174 155304
rect 308490 155292 308496 155304
rect 307588 155264 308496 155292
rect 241388 155196 294184 155224
rect 241388 155184 241394 155196
rect 294230 155184 294236 155236
rect 294288 155224 294294 155236
rect 300854 155224 300860 155236
rect 294288 155196 300860 155224
rect 294288 155184 294294 155196
rect 300854 155184 300860 155196
rect 300912 155184 300918 155236
rect 300946 155184 300952 155236
rect 301004 155224 301010 155236
rect 302878 155224 302884 155236
rect 301004 155196 302884 155224
rect 301004 155184 301010 155196
rect 302878 155184 302884 155196
rect 302936 155184 302942 155236
rect 304350 155184 304356 155236
rect 304408 155224 304414 155236
rect 306374 155224 306380 155236
rect 304408 155196 306380 155224
rect 304408 155184 304414 155196
rect 306374 155184 306380 155196
rect 306432 155184 306438 155236
rect 306926 155184 306932 155236
rect 306984 155224 306990 155236
rect 307588 155224 307616 155264
rect 308490 155252 308496 155264
rect 308548 155252 308554 155304
rect 308582 155252 308588 155304
rect 308640 155292 308646 155304
rect 341058 155292 341064 155304
rect 308640 155264 341064 155292
rect 308640 155252 308646 155264
rect 341058 155252 341064 155264
rect 341116 155252 341122 155304
rect 348786 155292 348792 155304
rect 341168 155264 348792 155292
rect 306984 155196 307616 155224
rect 306984 155184 306990 155196
rect 307662 155184 307668 155236
rect 307720 155224 307726 155236
rect 341168 155224 341196 155264
rect 348786 155252 348792 155264
rect 348844 155252 348850 155304
rect 351270 155252 351276 155304
rect 351328 155292 351334 155304
rect 355410 155292 355416 155304
rect 351328 155264 355416 155292
rect 351328 155252 351334 155264
rect 355410 155252 355416 155264
rect 355468 155252 355474 155304
rect 357406 155292 357434 155332
rect 362310 155320 362316 155372
rect 362368 155360 362374 155372
rect 394878 155360 394884 155372
rect 362368 155332 394884 155360
rect 362368 155320 362374 155332
rect 394878 155320 394884 155332
rect 394936 155320 394942 155372
rect 406838 155320 406844 155372
rect 406896 155360 406902 155372
rect 422662 155360 422668 155372
rect 406896 155332 422668 155360
rect 406896 155320 406902 155332
rect 422662 155320 422668 155332
rect 422720 155320 422726 155372
rect 422754 155320 422760 155372
rect 422812 155360 422818 155372
rect 424962 155360 424968 155372
rect 422812 155332 424968 155360
rect 422812 155320 422818 155332
rect 424962 155320 424968 155332
rect 425020 155320 425026 155372
rect 437014 155320 437020 155372
rect 437072 155360 437078 155372
rect 451274 155360 451280 155372
rect 437072 155332 451280 155360
rect 437072 155320 437078 155332
rect 451274 155320 451280 155332
rect 451332 155320 451338 155372
rect 452856 155332 453068 155360
rect 358446 155292 358452 155304
rect 357406 155264 358452 155292
rect 358446 155252 358452 155264
rect 358504 155252 358510 155304
rect 364702 155252 364708 155304
rect 364760 155292 364766 155304
rect 392394 155292 392400 155304
rect 364760 155264 392400 155292
rect 364760 155252 364766 155264
rect 392394 155252 392400 155264
rect 392452 155252 392458 155304
rect 395062 155252 395068 155304
rect 395120 155292 395126 155304
rect 405642 155292 405648 155304
rect 395120 155264 405648 155292
rect 395120 155252 395126 155264
rect 405642 155252 405648 155264
rect 405700 155252 405706 155304
rect 420270 155252 420276 155304
rect 420328 155292 420334 155304
rect 440234 155292 440240 155304
rect 420328 155264 440240 155292
rect 420328 155252 420334 155264
rect 440234 155252 440240 155264
rect 440292 155252 440298 155304
rect 442902 155252 442908 155304
rect 442960 155292 442966 155304
rect 452856 155292 452884 155332
rect 442960 155264 452884 155292
rect 453040 155292 453068 155332
rect 453114 155320 453120 155372
rect 453172 155360 453178 155372
rect 465074 155360 465080 155372
rect 453172 155332 465080 155360
rect 453172 155320 453178 155332
rect 465074 155320 465080 155332
rect 465132 155320 465138 155372
rect 465626 155320 465632 155372
rect 465684 155360 465690 155372
rect 474918 155360 474924 155372
rect 465684 155332 474924 155360
rect 465684 155320 465690 155332
rect 474918 155320 474924 155332
rect 474976 155320 474982 155372
rect 489914 155320 489920 155372
rect 489972 155360 489978 155372
rect 493226 155360 493232 155372
rect 489972 155332 493232 155360
rect 489972 155320 489978 155332
rect 493226 155320 493232 155332
rect 493284 155320 493290 155372
rect 495802 155320 495808 155372
rect 495860 155360 495866 155372
rect 496906 155360 496912 155372
rect 495860 155332 496912 155360
rect 495860 155320 495866 155332
rect 496906 155320 496912 155332
rect 496964 155320 496970 155372
rect 518066 155320 518072 155372
rect 518124 155360 518130 155372
rect 521838 155360 521844 155372
rect 518124 155332 521844 155360
rect 518124 155320 518130 155332
rect 521838 155320 521844 155332
rect 521896 155320 521902 155372
rect 456794 155292 456800 155304
rect 453040 155264 456800 155292
rect 442960 155252 442966 155264
rect 456794 155252 456800 155264
rect 456852 155252 456858 155304
rect 462222 155252 462228 155304
rect 462280 155292 462286 155304
rect 472342 155292 472348 155304
rect 462280 155264 472348 155292
rect 462280 155252 462286 155264
rect 472342 155252 472348 155264
rect 472400 155252 472406 155304
rect 473170 155252 473176 155304
rect 473228 155292 473234 155304
rect 477678 155292 477684 155304
rect 473228 155264 477684 155292
rect 473228 155252 473234 155264
rect 477678 155252 477684 155264
rect 477736 155252 477742 155304
rect 479886 155252 479892 155304
rect 479944 155292 479950 155304
rect 485682 155292 485688 155304
rect 479944 155264 485688 155292
rect 479944 155252 479950 155264
rect 485682 155252 485688 155264
rect 485740 155252 485746 155304
rect 487430 155252 487436 155304
rect 487488 155292 487494 155304
rect 491202 155292 491208 155304
rect 487488 155264 491208 155292
rect 487488 155252 487494 155264
rect 491202 155252 491208 155264
rect 491260 155252 491266 155304
rect 494974 155252 494980 155304
rect 495032 155292 495038 155304
rect 497366 155292 497372 155304
rect 495032 155264 497372 155292
rect 495032 155252 495038 155264
rect 497366 155252 497372 155264
rect 497424 155252 497430 155304
rect 512914 155252 512920 155304
rect 512972 155292 512978 155304
rect 515122 155292 515128 155304
rect 512972 155264 515128 155292
rect 512972 155252 512978 155264
rect 515122 155252 515128 155264
rect 515180 155252 515186 155304
rect 518802 155252 518808 155304
rect 518860 155292 518866 155304
rect 522666 155292 522672 155304
rect 518860 155264 522672 155292
rect 518860 155252 518866 155264
rect 522666 155252 522672 155264
rect 522724 155252 522730 155304
rect 307720 155196 341196 155224
rect 307720 155184 307726 155196
rect 341242 155184 341248 155236
rect 341300 155224 341306 155236
rect 344922 155224 344928 155236
rect 341300 155196 344928 155224
rect 341300 155184 341306 155196
rect 344922 155184 344928 155196
rect 344980 155184 344986 155236
rect 355594 155184 355600 155236
rect 355652 155224 355658 155236
rect 390738 155224 390744 155236
rect 355652 155196 390744 155224
rect 355652 155184 355658 155196
rect 390738 155184 390744 155196
rect 390796 155184 390802 155236
rect 404262 155184 404268 155236
rect 404320 155224 404326 155236
rect 427722 155224 427728 155236
rect 404320 155196 427728 155224
rect 404320 155184 404326 155196
rect 427722 155184 427728 155196
rect 427780 155184 427786 155236
rect 434530 155184 434536 155236
rect 434588 155224 434594 155236
rect 448514 155224 448520 155236
rect 434588 155196 448520 155224
rect 434588 155184 434594 155196
rect 448514 155184 448520 155196
rect 448572 155184 448578 155236
rect 454586 155184 454592 155236
rect 454644 155224 454650 155236
rect 462314 155224 462320 155236
rect 454644 155196 462320 155224
rect 454644 155184 454650 155196
rect 462314 155184 462320 155196
rect 462372 155184 462378 155236
rect 467282 155184 467288 155236
rect 467340 155224 467346 155236
rect 476206 155224 476212 155236
rect 467340 155196 476212 155224
rect 467340 155184 467346 155196
rect 476206 155184 476212 155196
rect 476264 155184 476270 155236
rect 493318 155184 493324 155236
rect 493376 155224 493382 155236
rect 495802 155224 495808 155236
rect 493376 155196 495808 155224
rect 493376 155184 493382 155196
rect 495802 155184 495808 155196
rect 495860 155184 495866 155236
rect 503346 155184 503352 155236
rect 503404 155224 503410 155236
rect 503806 155224 503812 155236
rect 503404 155196 503812 155224
rect 503404 155184 503410 155196
rect 503806 155184 503812 155196
rect 503864 155184 503870 155236
rect 510982 155184 510988 155236
rect 511040 155224 511046 155236
rect 512638 155224 512644 155236
rect 511040 155196 512644 155224
rect 511040 155184 511046 155196
rect 512638 155184 512644 155196
rect 512696 155184 512702 155236
rect 516778 155184 516784 155236
rect 516836 155224 516842 155236
rect 520182 155224 520188 155236
rect 516836 155196 520188 155224
rect 516836 155184 516842 155196
rect 520182 155184 520188 155196
rect 520240 155184 520246 155236
rect 521838 155184 521844 155236
rect 521896 155224 521902 155236
rect 523494 155224 523500 155236
rect 521896 155196 523500 155224
rect 521896 155184 521902 155196
rect 523494 155184 523500 155196
rect 523552 155184 523558 155236
rect 90174 155116 90180 155168
rect 90232 155156 90238 155168
rect 175826 155156 175832 155168
rect 90232 155128 175832 155156
rect 90232 155116 90238 155128
rect 175826 155116 175832 155128
rect 175884 155116 175890 155168
rect 175918 155116 175924 155168
rect 175976 155156 175982 155168
rect 191098 155156 191104 155168
rect 175976 155128 191104 155156
rect 175976 155116 175982 155128
rect 191098 155116 191104 155128
rect 191156 155116 191162 155168
rect 191190 155116 191196 155168
rect 191248 155156 191254 155168
rect 249150 155156 249156 155168
rect 191248 155128 249156 155156
rect 191248 155116 191254 155128
rect 249150 155116 249156 155128
rect 249208 155116 249214 155168
rect 253106 155116 253112 155168
rect 253164 155156 253170 155168
rect 272610 155156 272616 155168
rect 253164 155128 272616 155156
rect 253164 155116 253170 155128
rect 272610 155116 272616 155128
rect 272668 155116 272674 155168
rect 273254 155116 273260 155168
rect 273312 155156 273318 155168
rect 282086 155156 282092 155168
rect 273312 155128 282092 155156
rect 273312 155116 273318 155128
rect 282086 155116 282092 155128
rect 282144 155116 282150 155168
rect 282178 155116 282184 155168
rect 282236 155156 282242 155168
rect 283282 155156 283288 155168
rect 282236 155128 283288 155156
rect 282236 155116 282242 155128
rect 283282 155116 283288 155128
rect 283340 155116 283346 155168
rect 283374 155116 283380 155168
rect 283432 155156 283438 155168
rect 284294 155156 284300 155168
rect 283432 155128 284300 155156
rect 283432 155116 283438 155128
rect 284294 155116 284300 155128
rect 284352 155116 284358 155168
rect 286686 155116 286692 155168
rect 286744 155156 286750 155168
rect 292298 155156 292304 155168
rect 286744 155128 292304 155156
rect 286744 155116 286750 155128
rect 292298 155116 292304 155128
rect 292356 155116 292362 155168
rect 292574 155116 292580 155168
rect 292632 155156 292638 155168
rect 295610 155156 295616 155168
rect 292632 155128 295616 155156
rect 292632 155116 292638 155128
rect 295610 155116 295616 155128
rect 295668 155116 295674 155168
rect 295702 155116 295708 155168
rect 295760 155156 295766 155168
rect 326430 155156 326436 155168
rect 295760 155128 326436 155156
rect 295760 155116 295766 155128
rect 326430 155116 326436 155128
rect 326488 155116 326494 155168
rect 326982 155116 326988 155168
rect 327040 155156 327046 155168
rect 351270 155156 351276 155168
rect 327040 155128 351276 155156
rect 327040 155116 327046 155128
rect 351270 155116 351276 155128
rect 351328 155116 351334 155168
rect 351822 155116 351828 155168
rect 351880 155156 351886 155168
rect 387610 155156 387616 155168
rect 351880 155128 387616 155156
rect 351880 155116 351886 155128
rect 387610 155116 387616 155128
rect 387668 155116 387674 155168
rect 391658 155116 391664 155168
rect 391716 155156 391722 155168
rect 404170 155156 404176 155168
rect 391716 155128 404176 155156
rect 391716 155116 391722 155128
rect 404170 155116 404176 155128
rect 404228 155116 404234 155168
rect 416038 155116 416044 155168
rect 416096 155156 416102 155168
rect 422570 155156 422576 155168
rect 416096 155128 422576 155156
rect 416096 155116 416102 155128
rect 422570 155116 422576 155128
rect 422628 155116 422634 155168
rect 422662 155116 422668 155168
rect 422720 155156 422726 155168
rect 429930 155156 429936 155168
rect 422720 155128 429936 155156
rect 422720 155116 422726 155128
rect 429930 155116 429936 155128
rect 429988 155116 429994 155168
rect 437842 155116 437848 155168
rect 437900 155156 437906 155168
rect 453206 155156 453212 155168
rect 437900 155128 453212 155156
rect 437900 155116 437906 155128
rect 453206 155116 453212 155128
rect 453264 155116 453270 155168
rect 457990 155116 457996 155168
rect 458048 155156 458054 155168
rect 468018 155156 468024 155168
rect 458048 155128 468024 155156
rect 458048 155116 458054 155128
rect 468018 155116 468024 155128
rect 468076 155116 468082 155168
rect 484854 155116 484860 155168
rect 484912 155156 484918 155168
rect 488442 155156 488448 155168
rect 484912 155128 488448 155156
rect 484912 155116 484918 155128
rect 488442 155116 488448 155128
rect 488500 155116 488506 155168
rect 489086 155116 489092 155168
rect 489144 155156 489150 155168
rect 492582 155156 492588 155168
rect 489144 155128 492588 155156
rect 489144 155116 489150 155128
rect 492582 155116 492588 155128
rect 492640 155116 492646 155168
rect 84194 155048 84200 155100
rect 84252 155088 84258 155100
rect 91094 155088 91100 155100
rect 84252 155060 91100 155088
rect 84252 155048 84258 155060
rect 91094 155048 91100 155060
rect 91152 155048 91158 155100
rect 96890 155048 96896 155100
rect 96948 155088 96954 155100
rect 184198 155088 184204 155100
rect 96948 155060 184204 155088
rect 96948 155048 96954 155060
rect 184198 155048 184204 155060
rect 184256 155048 184262 155100
rect 184290 155048 184296 155100
rect 184348 155088 184354 155100
rect 186130 155088 186136 155100
rect 184348 155060 186136 155088
rect 184348 155048 184354 155060
rect 186130 155048 186136 155060
rect 186188 155048 186194 155100
rect 187510 155048 187516 155100
rect 187568 155088 187574 155100
rect 190822 155088 190828 155100
rect 187568 155060 190828 155088
rect 187568 155048 187574 155060
rect 190822 155048 190828 155060
rect 190880 155048 190886 155100
rect 191006 155048 191012 155100
rect 191064 155088 191070 155100
rect 200482 155088 200488 155100
rect 191064 155060 200488 155088
rect 191064 155048 191070 155060
rect 200482 155048 200488 155060
rect 200540 155048 200546 155100
rect 200758 155048 200764 155100
rect 200816 155088 200822 155100
rect 260190 155088 260196 155100
rect 200816 155060 260196 155088
rect 200816 155048 200822 155060
rect 260190 155048 260196 155060
rect 260248 155048 260254 155100
rect 261386 155048 261392 155100
rect 261444 155088 261450 155100
rect 262766 155088 262772 155100
rect 261444 155060 262772 155088
rect 261444 155048 261450 155060
rect 262766 155048 262772 155060
rect 262824 155048 262830 155100
rect 262858 155048 262864 155100
rect 262916 155088 262922 155100
rect 269022 155088 269028 155100
rect 262916 155060 269028 155088
rect 262916 155048 262922 155060
rect 269022 155048 269028 155060
rect 269080 155048 269086 155100
rect 269942 155048 269948 155100
rect 270000 155088 270006 155100
rect 299382 155088 299388 155100
rect 270000 155060 299388 155088
rect 270000 155048 270006 155060
rect 299382 155048 299388 155060
rect 299440 155048 299446 155100
rect 300854 155048 300860 155100
rect 300912 155088 300918 155100
rect 335998 155088 336004 155100
rect 300912 155060 336004 155088
rect 300912 155048 300918 155060
rect 335998 155048 336004 155060
rect 336056 155048 336062 155100
rect 336090 155048 336096 155100
rect 336148 155088 336154 155100
rect 341150 155088 341156 155100
rect 336148 155060 341156 155088
rect 336148 155048 336154 155060
rect 341150 155048 341156 155060
rect 341208 155048 341214 155100
rect 341334 155048 341340 155100
rect 341392 155088 341398 155100
rect 342070 155088 342076 155100
rect 341392 155060 342076 155088
rect 341392 155048 341398 155060
rect 342070 155048 342076 155060
rect 342128 155048 342134 155100
rect 343818 155048 343824 155100
rect 343876 155088 343882 155100
rect 377214 155088 377220 155100
rect 343876 155060 377220 155088
rect 343876 155048 343882 155060
rect 377214 155048 377220 155060
rect 377272 155048 377278 155100
rect 380802 155048 380808 155100
rect 380860 155088 380866 155100
rect 384482 155088 384488 155100
rect 380860 155060 384488 155088
rect 380860 155048 380866 155060
rect 384482 155048 384488 155060
rect 384540 155048 384546 155100
rect 384574 155048 384580 155100
rect 384632 155088 384638 155100
rect 395430 155088 395436 155100
rect 384632 155060 395436 155088
rect 384632 155048 384638 155060
rect 395430 155048 395436 155060
rect 395488 155048 395494 155100
rect 408494 155048 408500 155100
rect 408552 155088 408558 155100
rect 411714 155088 411720 155100
rect 408552 155060 411720 155088
rect 408552 155048 408558 155060
rect 411714 155048 411720 155060
rect 411772 155048 411778 155100
rect 436186 155048 436192 155100
rect 436244 155088 436250 155100
rect 451366 155088 451372 155100
rect 436244 155060 451372 155088
rect 436244 155048 436250 155060
rect 451366 155048 451372 155060
rect 451424 155048 451430 155100
rect 451458 155048 451464 155100
rect 451516 155088 451522 155100
rect 463694 155088 463700 155100
rect 451516 155060 463700 155088
rect 451516 155048 451522 155060
rect 463694 155048 463700 155060
rect 463752 155048 463758 155100
rect 470686 155048 470692 155100
rect 470744 155088 470750 155100
rect 477402 155088 477408 155100
rect 470744 155060 477408 155088
rect 470744 155048 470750 155060
rect 477402 155048 477408 155060
rect 477460 155048 477466 155100
rect 64138 154980 64144 155032
rect 64196 155020 64202 155032
rect 64196 154992 113312 155020
rect 64196 154980 64202 154992
rect 57422 154912 57428 154964
rect 57480 154952 57486 154964
rect 103514 154952 103520 154964
rect 57480 154924 103520 154952
rect 57480 154912 57486 154924
rect 103514 154912 103520 154924
rect 103572 154912 103578 154964
rect 103606 154912 103612 154964
rect 103664 154952 103670 154964
rect 111794 154952 111800 154964
rect 103664 154924 111800 154952
rect 103664 154912 103670 154924
rect 111794 154912 111800 154924
rect 111852 154912 111858 154964
rect 113284 154952 113312 154992
rect 114554 154980 114560 155032
rect 114612 155020 114618 155032
rect 115750 155020 115756 155032
rect 114612 154992 115756 155020
rect 114612 154980 114618 154992
rect 115750 154980 115756 154992
rect 115808 154980 115814 155032
rect 115934 154980 115940 155032
rect 115992 155020 115998 155032
rect 117130 155020 117136 155032
rect 115992 154992 117136 155020
rect 115992 154980 115998 154992
rect 117130 154980 117136 154992
rect 117188 154980 117194 155032
rect 117222 154980 117228 155032
rect 117280 155020 117286 155032
rect 120626 155020 120632 155032
rect 117280 154992 120632 155020
rect 117280 154980 117286 154992
rect 120626 154980 120632 154992
rect 120684 154980 120690 155032
rect 123386 155020 123392 155032
rect 120736 154992 123392 155020
rect 120736 154952 120764 154992
rect 123386 154980 123392 154992
rect 123444 154980 123450 155032
rect 123754 154980 123760 155032
rect 123812 155020 123818 155032
rect 128262 155020 128268 155032
rect 123812 154992 128268 155020
rect 123812 154980 123818 154992
rect 128262 154980 128268 154992
rect 128320 154980 128326 155032
rect 130470 154980 130476 155032
rect 130528 155020 130534 155032
rect 133230 155020 133236 155032
rect 130528 154992 133236 155020
rect 130528 154980 130534 154992
rect 133230 154980 133236 154992
rect 133288 154980 133294 155032
rect 133874 154980 133880 155032
rect 133932 155020 133938 155032
rect 133932 154992 137232 155020
rect 133932 154980 133938 154992
rect 128538 154952 128544 154964
rect 113284 154924 120764 154952
rect 122208 154924 128544 154952
rect 79318 154844 79324 154896
rect 79376 154884 79382 154896
rect 113174 154884 113180 154896
rect 79376 154856 113180 154884
rect 79376 154844 79382 154856
rect 113174 154844 113180 154856
rect 113232 154844 113238 154896
rect 116578 154884 116584 154896
rect 113284 154856 116584 154884
rect 86034 154776 86040 154828
rect 86092 154816 86098 154828
rect 113284 154816 113312 154856
rect 116578 154844 116584 154856
rect 116636 154844 116642 154896
rect 117038 154844 117044 154896
rect 117096 154884 117102 154896
rect 122208 154884 122236 154924
rect 128538 154912 128544 154924
rect 128596 154912 128602 154964
rect 134610 154912 134616 154964
rect 134668 154952 134674 154964
rect 136910 154952 136916 154964
rect 134668 154924 136916 154952
rect 134668 154912 134674 154924
rect 136910 154912 136916 154924
rect 136968 154912 136974 154964
rect 137204 154952 137232 154992
rect 137646 154980 137652 155032
rect 137704 155020 137710 155032
rect 213086 155020 213092 155032
rect 137704 154992 213092 155020
rect 137704 154980 137710 154992
rect 213086 154980 213092 154992
rect 213144 154980 213150 155032
rect 213638 154980 213644 155032
rect 213696 155020 213702 155032
rect 216490 155020 216496 155032
rect 213696 154992 216496 155020
rect 213696 154980 213702 154992
rect 216490 154980 216496 154992
rect 216548 154980 216554 155032
rect 221182 154980 221188 155032
rect 221240 155020 221246 155032
rect 279878 155020 279884 155032
rect 221240 154992 279884 155020
rect 221240 154980 221246 154992
rect 279878 154980 279884 154992
rect 279936 154980 279942 155032
rect 279970 154980 279976 155032
rect 280028 155020 280034 155032
rect 287698 155020 287704 155032
rect 280028 154992 287704 155020
rect 280028 154980 280034 154992
rect 287698 154980 287704 154992
rect 287756 154980 287762 155032
rect 288342 154980 288348 155032
rect 288400 155020 288406 155032
rect 321922 155020 321928 155032
rect 288400 154992 321928 155020
rect 288400 154980 288406 154992
rect 321922 154980 321928 154992
rect 321980 154980 321986 155032
rect 322106 154980 322112 155032
rect 322164 155020 322170 155032
rect 325970 155020 325976 155032
rect 322164 154992 325976 155020
rect 322164 154980 322170 154992
rect 325970 154980 325976 154992
rect 326028 154980 326034 155032
rect 326338 154980 326344 155032
rect 326396 155020 326402 155032
rect 355226 155020 355232 155032
rect 326396 154992 340736 155020
rect 326396 154980 326402 154992
rect 211890 154952 211896 154964
rect 137204 154924 211896 154952
rect 211890 154912 211896 154924
rect 211948 154912 211954 154964
rect 211982 154912 211988 154964
rect 212040 154952 212046 154964
rect 212442 154952 212448 154964
rect 212040 154924 212448 154952
rect 212040 154912 212046 154924
rect 212442 154912 212448 154924
rect 212500 154912 212506 154964
rect 212534 154912 212540 154964
rect 212592 154952 212598 154964
rect 214374 154952 214380 154964
rect 212592 154924 214380 154952
rect 212592 154912 212598 154924
rect 214374 154912 214380 154924
rect 214432 154912 214438 154964
rect 214558 154912 214564 154964
rect 214616 154952 214622 154964
rect 232038 154952 232044 154964
rect 214616 154924 232044 154952
rect 214616 154912 214622 154924
rect 232038 154912 232044 154924
rect 232096 154912 232102 154964
rect 232314 154912 232320 154964
rect 232372 154952 232378 154964
rect 241422 154952 241428 154964
rect 232372 154924 241428 154952
rect 232372 154912 232378 154924
rect 241422 154912 241428 154924
rect 241480 154912 241486 154964
rect 243538 154912 243544 154964
rect 243596 154952 243602 154964
rect 292390 154952 292396 154964
rect 243596 154924 292396 154952
rect 243596 154912 243602 154924
rect 292390 154912 292396 154924
rect 292448 154912 292454 154964
rect 294046 154912 294052 154964
rect 294104 154952 294110 154964
rect 306926 154952 306932 154964
rect 294104 154924 306932 154952
rect 294104 154912 294110 154924
rect 306926 154912 306932 154924
rect 306984 154912 306990 154964
rect 307202 154912 307208 154964
rect 307260 154952 307266 154964
rect 321830 154952 321836 154964
rect 307260 154924 321836 154952
rect 307260 154912 307266 154924
rect 321830 154912 321836 154924
rect 321888 154912 321894 154964
rect 322198 154912 322204 154964
rect 322256 154952 322262 154964
rect 340506 154952 340512 154964
rect 322256 154924 340512 154952
rect 322256 154912 322262 154924
rect 340506 154912 340512 154924
rect 340564 154912 340570 154964
rect 340708 154952 340736 154992
rect 340984 154992 355232 155020
rect 340984 154952 341012 154992
rect 355226 154980 355232 154992
rect 355284 154980 355290 155032
rect 355410 154980 355416 155032
rect 355468 155020 355474 155032
rect 357434 155020 357440 155032
rect 355468 154992 357440 155020
rect 355468 154980 355474 154992
rect 357434 154980 357440 154992
rect 357492 154980 357498 155032
rect 371510 154980 371516 155032
rect 371568 155020 371574 155032
rect 396442 155020 396448 155032
rect 371568 154992 383654 155020
rect 371568 154980 371574 154992
rect 340708 154924 341012 154952
rect 341058 154912 341064 154964
rect 341116 154952 341122 154964
rect 348786 154952 348792 154964
rect 341116 154924 348792 154952
rect 341116 154912 341122 154924
rect 348786 154912 348792 154924
rect 348844 154912 348850 154964
rect 355318 154952 355324 154964
rect 351564 154924 355324 154952
rect 117096 154856 122236 154884
rect 117096 154844 117102 154856
rect 127158 154844 127164 154896
rect 127216 154884 127222 154896
rect 137370 154884 137376 154896
rect 127216 154856 137376 154884
rect 127216 154844 127222 154856
rect 137370 154844 137376 154856
rect 137428 154844 137434 154896
rect 137554 154844 137560 154896
rect 137612 154884 137618 154896
rect 144822 154884 144828 154896
rect 137612 154856 144828 154884
rect 137612 154844 137618 154856
rect 144822 154844 144828 154856
rect 144880 154844 144886 154896
rect 146938 154844 146944 154896
rect 146996 154884 147002 154896
rect 155862 154884 155868 154896
rect 146996 154856 155868 154884
rect 146996 154844 147002 154856
rect 155862 154844 155868 154856
rect 155920 154844 155926 154896
rect 161198 154884 161204 154896
rect 155972 154856 161204 154884
rect 86092 154788 113312 154816
rect 86092 154776 86098 154788
rect 113450 154776 113456 154828
rect 113508 154816 113514 154828
rect 120534 154816 120540 154828
rect 113508 154788 120540 154816
rect 113508 154776 113514 154788
rect 120534 154776 120540 154788
rect 120592 154776 120598 154828
rect 120626 154776 120632 154828
rect 120684 154816 120690 154828
rect 153010 154816 153016 154828
rect 120684 154788 153016 154816
rect 120684 154776 120690 154788
rect 153010 154776 153016 154788
rect 153068 154776 153074 154828
rect 153102 154776 153108 154828
rect 153160 154816 153166 154828
rect 155972 154816 156000 154856
rect 161198 154844 161204 154856
rect 161256 154844 161262 154896
rect 161290 154844 161296 154896
rect 161348 154884 161354 154896
rect 164234 154884 164240 154896
rect 161348 154856 164240 154884
rect 161348 154844 161354 154856
rect 164234 154844 164240 154856
rect 164292 154844 164298 154896
rect 164326 154844 164332 154896
rect 164384 154884 164390 154896
rect 233694 154884 233700 154896
rect 164384 154856 233700 154884
rect 164384 154844 164390 154856
rect 233694 154844 233700 154856
rect 233752 154844 233758 154896
rect 233786 154844 233792 154896
rect 233844 154884 233850 154896
rect 233844 154856 237972 154884
rect 233844 154844 233850 154856
rect 153160 154788 156000 154816
rect 153160 154776 153166 154788
rect 156598 154776 156604 154828
rect 156656 154816 156662 154828
rect 220722 154816 220728 154828
rect 156656 154788 161428 154816
rect 156656 154776 156662 154788
rect 103514 154708 103520 154760
rect 103572 154748 103578 154760
rect 109126 154748 109132 154760
rect 103572 154720 109132 154748
rect 103572 154708 103578 154720
rect 109126 154708 109132 154720
rect 109184 154708 109190 154760
rect 109402 154708 109408 154760
rect 109460 154748 109466 154760
rect 161290 154748 161296 154760
rect 109460 154720 161296 154748
rect 109460 154708 109466 154720
rect 161290 154708 161296 154720
rect 161348 154708 161354 154760
rect 161400 154748 161428 154788
rect 161952 154788 220728 154816
rect 161952 154748 161980 154788
rect 220722 154776 220728 154788
rect 220780 154776 220786 154828
rect 223758 154776 223764 154828
rect 223816 154816 223822 154828
rect 226978 154816 226984 154828
rect 223816 154788 226984 154816
rect 223816 154776 223822 154788
rect 226978 154776 226984 154788
rect 227036 154776 227042 154828
rect 227070 154776 227076 154828
rect 227128 154816 227134 154828
rect 233878 154816 233884 154828
rect 227128 154788 233884 154816
rect 227128 154776 227134 154788
rect 233878 154776 233884 154788
rect 233936 154776 233942 154828
rect 233970 154776 233976 154828
rect 234028 154816 234034 154828
rect 237374 154816 237380 154828
rect 234028 154788 237380 154816
rect 234028 154776 234034 154788
rect 237374 154776 237380 154788
rect 237432 154776 237438 154828
rect 237944 154816 237972 154856
rect 238018 154844 238024 154896
rect 238076 154884 238082 154896
rect 238754 154884 238760 154896
rect 238076 154856 238760 154884
rect 238076 154844 238082 154856
rect 238754 154844 238760 154856
rect 238812 154844 238818 154896
rect 238846 154844 238852 154896
rect 238904 154884 238910 154896
rect 247126 154884 247132 154896
rect 238904 154856 247132 154884
rect 238904 154844 238910 154856
rect 247126 154844 247132 154856
rect 247184 154844 247190 154896
rect 247218 154844 247224 154896
rect 247276 154884 247282 154896
rect 247276 154856 293356 154884
rect 247276 154844 247282 154856
rect 238570 154816 238576 154828
rect 237944 154788 238576 154816
rect 238570 154776 238576 154788
rect 238628 154776 238634 154828
rect 238662 154776 238668 154828
rect 238720 154816 238726 154828
rect 238720 154788 238984 154816
rect 238720 154776 238726 154788
rect 161400 154720 161980 154748
rect 162118 154708 162124 154760
rect 162176 154748 162182 154760
rect 167638 154748 167644 154760
rect 162176 154720 167644 154748
rect 162176 154708 162182 154720
rect 167638 154708 167644 154720
rect 167696 154708 167702 154760
rect 175826 154708 175832 154760
rect 175884 154748 175890 154760
rect 183278 154748 183284 154760
rect 175884 154720 183284 154748
rect 175884 154708 175890 154720
rect 183278 154708 183284 154720
rect 183336 154708 183342 154760
rect 184198 154708 184204 154760
rect 184256 154748 184262 154760
rect 184256 154720 185072 154748
rect 184256 154708 184262 154720
rect 99466 154640 99472 154692
rect 99524 154680 99530 154692
rect 116762 154680 116768 154692
rect 99524 154652 116768 154680
rect 99524 154640 99530 154652
rect 116762 154640 116768 154652
rect 116820 154640 116826 154692
rect 116854 154640 116860 154692
rect 116912 154680 116918 154692
rect 121270 154680 121276 154692
rect 116912 154652 121276 154680
rect 116912 154640 116918 154652
rect 121270 154640 121276 154652
rect 121328 154640 121334 154692
rect 122926 154640 122932 154692
rect 122984 154680 122990 154692
rect 122984 154652 128354 154680
rect 122984 154640 122990 154652
rect 92750 154572 92756 154624
rect 92808 154612 92814 154624
rect 113634 154612 113640 154624
rect 92808 154584 113640 154612
rect 92808 154572 92814 154584
rect 113634 154572 113640 154584
rect 113692 154572 113698 154624
rect 113726 154572 113732 154624
rect 113784 154612 113790 154624
rect 123478 154612 123484 154624
rect 113784 154584 123484 154612
rect 113784 154572 113790 154584
rect 123478 154572 123484 154584
rect 123536 154572 123542 154624
rect 128326 154612 128354 154652
rect 128814 154640 128820 154692
rect 128872 154680 128878 154692
rect 129550 154680 129556 154692
rect 128872 154652 129556 154680
rect 128872 154640 128878 154652
rect 129550 154640 129556 154652
rect 129608 154640 129614 154692
rect 129642 154640 129648 154692
rect 129700 154680 129706 154692
rect 184934 154680 184940 154692
rect 129700 154652 184940 154680
rect 129700 154640 129706 154652
rect 184934 154640 184940 154652
rect 184992 154640 184998 154692
rect 184842 154612 184848 154624
rect 128326 154584 184848 154612
rect 184842 154572 184848 154584
rect 184900 154572 184906 154624
rect 185044 154612 185072 154720
rect 185486 154708 185492 154760
rect 185544 154748 185550 154760
rect 238754 154748 238760 154760
rect 185544 154720 238760 154748
rect 185544 154708 185550 154720
rect 238754 154708 238760 154720
rect 238812 154708 238818 154760
rect 238956 154748 238984 154788
rect 239030 154776 239036 154828
rect 239088 154816 239094 154828
rect 282178 154816 282184 154828
rect 239088 154788 282184 154816
rect 239088 154776 239094 154788
rect 282178 154776 282184 154788
rect 282236 154776 282242 154828
rect 285030 154776 285036 154828
rect 285088 154816 285094 154828
rect 287054 154816 287060 154828
rect 285088 154788 287060 154816
rect 285088 154776 285094 154788
rect 287054 154776 287060 154788
rect 287112 154776 287118 154828
rect 287514 154776 287520 154828
rect 287572 154816 287578 154828
rect 291194 154816 291200 154828
rect 287572 154788 291200 154816
rect 287572 154776 287578 154788
rect 291194 154776 291200 154788
rect 291252 154776 291258 154828
rect 292114 154776 292120 154828
rect 292172 154816 292178 154828
rect 293126 154816 293132 154828
rect 292172 154788 293132 154816
rect 292172 154776 292178 154788
rect 293126 154776 293132 154788
rect 293184 154776 293190 154828
rect 293328 154816 293356 154856
rect 293402 154844 293408 154896
rect 293460 154884 293466 154896
rect 321370 154884 321376 154896
rect 293460 154856 321376 154884
rect 293460 154844 293466 154856
rect 321370 154844 321376 154856
rect 321428 154844 321434 154896
rect 321922 154844 321928 154896
rect 321980 154884 321986 154896
rect 326522 154884 326528 154896
rect 321980 154856 326528 154884
rect 321980 154844 321986 154856
rect 326522 154844 326528 154856
rect 326580 154844 326586 154896
rect 326614 154844 326620 154896
rect 326672 154884 326678 154896
rect 351564 154884 351592 154924
rect 355318 154912 355324 154924
rect 355376 154912 355382 154964
rect 357250 154912 357256 154964
rect 357308 154952 357314 154964
rect 380986 154952 380992 154964
rect 357308 154924 380992 154952
rect 357308 154912 357314 154924
rect 380986 154912 380992 154924
rect 381044 154912 381050 154964
rect 383626 154952 383654 154992
rect 384592 154992 396448 155020
rect 384592 154952 384620 154992
rect 396442 154980 396448 154992
rect 396500 154980 396506 155032
rect 441246 154980 441252 155032
rect 441304 155020 441310 155032
rect 455414 155020 455420 155032
rect 441304 154992 455420 155020
rect 441304 154980 441310 154992
rect 455414 154980 455420 154992
rect 455472 154980 455478 155032
rect 455506 154980 455512 155032
rect 455564 155020 455570 155032
rect 455564 154992 457116 155020
rect 455564 154980 455570 154992
rect 383626 154924 384620 154952
rect 384666 154912 384672 154964
rect 384724 154952 384730 154964
rect 388530 154952 388536 154964
rect 384724 154924 388536 154952
rect 384724 154912 384730 154924
rect 388530 154912 388536 154924
rect 388588 154912 388594 154964
rect 392486 154912 392492 154964
rect 392544 154952 392550 154964
rect 415486 154952 415492 154964
rect 392544 154924 415492 154952
rect 392544 154912 392550 154924
rect 415486 154912 415492 154924
rect 415544 154912 415550 154964
rect 440418 154912 440424 154964
rect 440476 154952 440482 154964
rect 455690 154952 455696 154964
rect 440476 154924 455696 154952
rect 440476 154912 440482 154924
rect 455690 154912 455696 154924
rect 455748 154912 455754 154964
rect 457088 154952 457116 154992
rect 457162 154980 457168 155032
rect 457220 155020 457226 155032
rect 468478 155020 468484 155032
rect 457220 154992 468484 155020
rect 457220 154980 457226 154992
rect 468478 154980 468484 154992
rect 468536 154980 468542 155032
rect 473998 154980 474004 155032
rect 474056 155020 474062 155032
rect 479518 155020 479524 155032
rect 474056 154992 479524 155020
rect 474056 154980 474062 154992
rect 479518 154980 479524 154992
rect 479576 154980 479582 155032
rect 511626 154980 511632 155032
rect 511684 155020 511690 155032
rect 513466 155020 513472 155032
rect 511684 154992 513472 155020
rect 511684 154980 511690 154992
rect 513466 154980 513472 154992
rect 513524 154980 513530 155032
rect 467006 154952 467012 154964
rect 457088 154924 467012 154952
rect 467006 154912 467012 154924
rect 467064 154912 467070 154964
rect 326672 154856 351592 154884
rect 326672 154844 326678 154856
rect 351638 154844 351644 154896
rect 351696 154884 351702 154896
rect 364242 154884 364248 154896
rect 351696 154856 364248 154884
rect 351696 154844 351702 154856
rect 364242 154844 364248 154856
rect 364300 154844 364306 154896
rect 364978 154844 364984 154896
rect 365036 154884 365042 154896
rect 373994 154884 374000 154896
rect 365036 154856 374000 154884
rect 365036 154844 365042 154856
rect 373994 154844 374000 154856
rect 374052 154844 374058 154896
rect 374914 154844 374920 154896
rect 374972 154884 374978 154896
rect 398098 154884 398104 154896
rect 374972 154856 398104 154884
rect 374972 154844 374978 154856
rect 398098 154844 398104 154856
rect 398156 154844 398162 154896
rect 446306 154844 446312 154896
rect 446364 154884 446370 154896
rect 459646 154884 459652 154896
rect 446364 154856 459652 154884
rect 446364 154844 446370 154856
rect 459646 154844 459652 154856
rect 459704 154844 459710 154896
rect 294322 154816 294328 154828
rect 293328 154788 294328 154816
rect 294322 154776 294328 154788
rect 294380 154776 294386 154828
rect 306926 154816 306932 154828
rect 294616 154788 306932 154816
rect 281442 154748 281448 154760
rect 238956 154720 281448 154748
rect 281442 154708 281448 154720
rect 281500 154708 281506 154760
rect 282086 154708 282092 154760
rect 282144 154748 282150 154760
rect 294616 154748 294644 154788
rect 306926 154776 306932 154788
rect 306984 154776 306990 154828
rect 310238 154776 310244 154828
rect 310296 154816 310302 154828
rect 340322 154816 340328 154828
rect 310296 154788 340328 154816
rect 310296 154776 310302 154788
rect 340322 154776 340328 154788
rect 340380 154776 340386 154828
rect 363874 154816 363880 154828
rect 340708 154788 363880 154816
rect 282144 154720 294644 154748
rect 282144 154708 282150 154720
rect 294690 154708 294696 154760
rect 294748 154748 294754 154760
rect 301038 154748 301044 154760
rect 294748 154720 301044 154748
rect 294748 154708 294754 154720
rect 301038 154708 301044 154720
rect 301096 154708 301102 154760
rect 301866 154708 301872 154760
rect 301924 154748 301930 154760
rect 307018 154748 307024 154760
rect 301924 154720 307024 154748
rect 301924 154708 301930 154720
rect 307018 154708 307024 154720
rect 307076 154708 307082 154760
rect 307110 154708 307116 154760
rect 307168 154748 307174 154760
rect 307168 154720 311756 154748
rect 307168 154708 307174 154720
rect 185118 154640 185124 154692
rect 185176 154680 185182 154692
rect 193214 154680 193220 154692
rect 185176 154652 193220 154680
rect 185176 154640 185182 154652
rect 193214 154640 193220 154652
rect 193272 154640 193278 154692
rect 193490 154640 193496 154692
rect 193548 154680 193554 154692
rect 200758 154680 200764 154692
rect 193548 154652 200764 154680
rect 193548 154640 193554 154652
rect 200758 154640 200764 154652
rect 200816 154640 200822 154692
rect 200942 154640 200948 154692
rect 201000 154680 201006 154692
rect 209590 154680 209596 154692
rect 201000 154652 209596 154680
rect 201000 154640 201006 154652
rect 209590 154640 209596 154652
rect 209648 154640 209654 154692
rect 209682 154640 209688 154692
rect 209740 154680 209746 154692
rect 263594 154680 263600 154692
rect 209740 154652 263600 154680
rect 209740 154640 209746 154652
rect 263594 154640 263600 154652
rect 263652 154640 263658 154692
rect 263686 154640 263692 154692
rect 263744 154680 263750 154692
rect 264514 154680 264520 154692
rect 263744 154652 264520 154680
rect 263744 154640 263750 154652
rect 264514 154640 264520 154652
rect 264572 154640 264578 154692
rect 266538 154640 266544 154692
rect 266596 154680 266602 154692
rect 266596 154652 272564 154680
rect 266596 154640 266602 154652
rect 188982 154612 188988 154624
rect 185044 154584 188988 154612
rect 188982 154572 188988 154584
rect 189040 154572 189046 154624
rect 190914 154572 190920 154624
rect 190972 154612 190978 154624
rect 191834 154612 191840 154624
rect 190972 154584 191840 154612
rect 190972 154572 190978 154584
rect 191834 154572 191840 154584
rect 191892 154572 191898 154624
rect 192018 154572 192024 154624
rect 192076 154612 192082 154624
rect 194594 154612 194600 154624
rect 192076 154584 194600 154612
rect 192076 154572 192082 154584
rect 194594 154572 194600 154584
rect 194652 154572 194658 154624
rect 197722 154572 197728 154624
rect 197780 154612 197786 154624
rect 214558 154612 214564 154624
rect 197780 154584 214564 154612
rect 197780 154572 197786 154584
rect 214558 154572 214564 154584
rect 214616 154572 214622 154624
rect 216490 154572 216496 154624
rect 216548 154612 216554 154624
rect 271506 154612 271512 154624
rect 216548 154584 271512 154612
rect 216548 154572 216554 154584
rect 271506 154572 271512 154584
rect 271564 154572 271570 154624
rect 272536 154612 272564 154652
rect 272610 154640 272616 154692
rect 272668 154680 272674 154692
rect 278682 154680 278688 154692
rect 272668 154652 278688 154680
rect 272668 154640 272674 154652
rect 278682 154640 278688 154652
rect 278740 154640 278746 154692
rect 280798 154640 280804 154692
rect 280856 154680 280862 154692
rect 280856 154652 287652 154680
rect 280856 154640 280862 154652
rect 287514 154612 287520 154624
rect 272536 154584 287520 154612
rect 287514 154572 287520 154584
rect 287572 154572 287578 154624
rect 287624 154612 287652 154652
rect 287698 154640 287704 154692
rect 287756 154680 287762 154692
rect 311434 154680 311440 154692
rect 287756 154652 311440 154680
rect 287756 154640 287762 154652
rect 311434 154640 311440 154652
rect 311492 154640 311498 154692
rect 311728 154680 311756 154720
rect 311802 154708 311808 154760
rect 311860 154748 311866 154760
rect 313458 154748 313464 154760
rect 311860 154720 313464 154748
rect 311860 154708 311866 154720
rect 313458 154708 313464 154720
rect 313516 154708 313522 154760
rect 313550 154708 313556 154760
rect 313608 154748 313614 154760
rect 340230 154748 340236 154760
rect 313608 154720 340236 154748
rect 313608 154708 313614 154720
rect 340230 154708 340236 154720
rect 340288 154708 340294 154760
rect 311728 154652 321968 154680
rect 292206 154612 292212 154624
rect 287624 154584 292212 154612
rect 292206 154572 292212 154584
rect 292264 154572 292270 154624
rect 292482 154572 292488 154624
rect 292540 154612 292546 154624
rect 316586 154612 316592 154624
rect 292540 154584 316592 154612
rect 292540 154572 292546 154584
rect 316586 154572 316592 154584
rect 316644 154572 316650 154624
rect 316678 154572 316684 154624
rect 316736 154612 316742 154624
rect 321830 154612 321836 154624
rect 316736 154584 321836 154612
rect 316736 154572 316742 154584
rect 321830 154572 321836 154584
rect 321888 154572 321894 154624
rect 321940 154612 321968 154652
rect 322014 154640 322020 154692
rect 322072 154680 322078 154692
rect 326614 154680 326620 154692
rect 322072 154652 326620 154680
rect 322072 154640 322078 154652
rect 326614 154640 326620 154652
rect 326672 154640 326678 154692
rect 327902 154640 327908 154692
rect 327960 154680 327966 154692
rect 340708 154680 340736 154788
rect 363874 154776 363880 154788
rect 363932 154776 363938 154828
rect 363966 154776 363972 154828
rect 364024 154816 364030 154828
rect 386230 154816 386236 154828
rect 364024 154788 386236 154816
rect 364024 154776 364030 154788
rect 386230 154776 386236 154788
rect 386288 154776 386294 154828
rect 444558 154776 444564 154828
rect 444616 154816 444622 154828
rect 458358 154816 458364 154828
rect 444616 154788 458364 154816
rect 444616 154776 444622 154788
rect 458358 154776 458364 154788
rect 458416 154776 458422 154828
rect 463050 154776 463056 154828
rect 463108 154816 463114 154828
rect 471974 154816 471980 154828
rect 463108 154788 471980 154816
rect 463108 154776 463114 154788
rect 471974 154776 471980 154788
rect 472032 154776 472038 154828
rect 484026 154776 484032 154828
rect 484084 154816 484090 154828
rect 488994 154816 489000 154828
rect 484084 154788 489000 154816
rect 484084 154776 484090 154788
rect 488994 154776 489000 154788
rect 489052 154776 489058 154828
rect 509694 154776 509700 154828
rect 509752 154816 509758 154828
rect 510890 154816 510896 154828
rect 509752 154788 510896 154816
rect 509752 154776 509758 154788
rect 510890 154776 510896 154788
rect 510948 154776 510954 154828
rect 340874 154708 340880 154760
rect 340932 154748 340938 154760
rect 351822 154748 351828 154760
rect 340932 154720 351828 154748
rect 340932 154708 340938 154720
rect 351822 154708 351828 154720
rect 351880 154708 351886 154760
rect 353846 154708 353852 154760
rect 353904 154748 353910 154760
rect 380894 154748 380900 154760
rect 353904 154720 380900 154748
rect 353904 154708 353910 154720
rect 380894 154708 380900 154720
rect 380952 154708 380958 154760
rect 385678 154748 385684 154760
rect 383626 154720 385684 154748
rect 327960 154652 340736 154680
rect 327960 154640 327966 154652
rect 341150 154640 341156 154692
rect 341208 154680 341214 154692
rect 367094 154680 367100 154692
rect 341208 154652 367100 154680
rect 341208 154640 341214 154652
rect 367094 154640 367100 154652
rect 367152 154640 367158 154692
rect 367370 154640 367376 154692
rect 367428 154680 367434 154692
rect 383626 154680 383654 154720
rect 385678 154708 385684 154720
rect 385736 154708 385742 154760
rect 385770 154708 385776 154760
rect 385828 154748 385834 154760
rect 413186 154748 413192 154760
rect 385828 154720 413192 154748
rect 385828 154708 385834 154720
rect 413186 154708 413192 154720
rect 413244 154708 413250 154760
rect 445386 154708 445392 154760
rect 445444 154748 445450 154760
rect 458726 154748 458732 154760
rect 445444 154720 458732 154748
rect 445444 154708 445450 154720
rect 458726 154708 458732 154720
rect 458784 154708 458790 154760
rect 461486 154708 461492 154760
rect 461544 154748 461550 154760
rect 471698 154748 471704 154760
rect 461544 154720 471704 154748
rect 461544 154708 461550 154720
rect 471698 154708 471704 154720
rect 471756 154708 471762 154760
rect 485774 154708 485780 154760
rect 485832 154748 485838 154760
rect 488902 154748 488908 154760
rect 485832 154720 488908 154748
rect 485832 154708 485838 154720
rect 488902 154708 488908 154720
rect 488960 154708 488966 154760
rect 496630 154708 496636 154760
rect 496688 154748 496694 154760
rect 498194 154748 498200 154760
rect 496688 154720 498200 154748
rect 496688 154708 496694 154720
rect 498194 154708 498200 154720
rect 498252 154708 498258 154760
rect 367428 154652 383654 154680
rect 367428 154640 367434 154652
rect 387518 154640 387524 154692
rect 387576 154680 387582 154692
rect 390922 154680 390928 154692
rect 387576 154652 390928 154680
rect 387576 154640 387582 154652
rect 390922 154640 390928 154652
rect 390980 154640 390986 154692
rect 445202 154640 445208 154692
rect 445260 154680 445266 154692
rect 447226 154680 447232 154692
rect 445260 154652 447232 154680
rect 445260 154640 445266 154652
rect 447226 154640 447232 154652
rect 447284 154640 447290 154692
rect 448790 154640 448796 154692
rect 448848 154680 448854 154692
rect 459554 154680 459560 154692
rect 448848 154652 459560 154680
rect 448848 154640 448854 154652
rect 459554 154640 459560 154652
rect 459612 154640 459618 154692
rect 477310 154640 477316 154692
rect 477368 154680 477374 154692
rect 481726 154680 481732 154692
rect 477368 154652 481732 154680
rect 477368 154640 477374 154652
rect 481726 154640 481732 154652
rect 481784 154640 481790 154692
rect 326062 154612 326068 154624
rect 321940 154584 326068 154612
rect 326062 154572 326068 154584
rect 326120 154572 326126 154624
rect 326154 154572 326160 154624
rect 326212 154612 326218 154624
rect 332502 154612 332508 154624
rect 326212 154584 332508 154612
rect 326212 154572 326218 154584
rect 332502 154572 332508 154584
rect 332560 154572 332566 154624
rect 334618 154572 334624 154624
rect 334676 154612 334682 154624
rect 368474 154612 368480 154624
rect 334676 154584 368480 154612
rect 334676 154572 334682 154584
rect 368474 154572 368480 154584
rect 368532 154572 368538 154624
rect 374086 154572 374092 154624
rect 374144 154612 374150 154624
rect 388438 154612 388444 154624
rect 374144 154584 388444 154612
rect 374144 154572 374150 154584
rect 388438 154572 388444 154584
rect 388496 154572 388502 154624
rect 390830 154572 390836 154624
rect 390888 154612 390894 154624
rect 392302 154612 392308 154624
rect 390888 154584 392308 154612
rect 390888 154572 390894 154584
rect 392302 154572 392308 154584
rect 392360 154572 392366 154624
rect 447134 154572 447140 154624
rect 447192 154612 447198 154624
rect 458174 154612 458180 154624
rect 447192 154584 458180 154612
rect 447192 154572 447198 154584
rect 458174 154572 458180 154584
rect 458232 154572 458238 154624
rect 459738 154572 459744 154624
rect 459796 154612 459802 154624
rect 470410 154612 470416 154624
rect 459796 154584 470416 154612
rect 459796 154572 459802 154584
rect 470410 154572 470416 154584
rect 470468 154572 470474 154624
rect 486602 154572 486608 154624
rect 486660 154612 486666 154624
rect 488534 154612 488540 154624
rect 486660 154584 488540 154612
rect 486660 154572 486666 154584
rect 488534 154572 488540 154584
rect 488592 154572 488598 154624
rect 51534 154504 51540 154556
rect 51592 154544 51598 154556
rect 158346 154544 158352 154556
rect 51592 154516 158352 154544
rect 51592 154504 51598 154516
rect 158346 154504 158352 154516
rect 158404 154504 158410 154556
rect 159082 154504 159088 154556
rect 159140 154544 159146 154556
rect 238018 154544 238024 154556
rect 159140 154516 238024 154544
rect 159140 154504 159146 154516
rect 238018 154504 238024 154516
rect 238076 154504 238082 154556
rect 243078 154544 243084 154556
rect 238128 154516 243084 154544
rect 54938 154436 54944 154488
rect 54996 154476 55002 154488
rect 160922 154476 160928 154488
rect 54996 154448 160928 154476
rect 54996 154436 55002 154448
rect 160922 154436 160928 154448
rect 160980 154436 160986 154488
rect 162026 154436 162032 154488
rect 162084 154476 162090 154488
rect 238128 154476 238156 154516
rect 243078 154504 243084 154516
rect 243136 154504 243142 154556
rect 245562 154504 245568 154556
rect 245620 154544 245626 154556
rect 248782 154544 248788 154556
rect 245620 154516 248788 154544
rect 245620 154504 245626 154516
rect 248782 154504 248788 154516
rect 248840 154504 248846 154556
rect 248874 154504 248880 154556
rect 248932 154544 248938 154556
rect 248932 154516 306880 154544
rect 248932 154504 248938 154516
rect 162084 154448 238156 154476
rect 162084 154436 162090 154448
rect 238938 154436 238944 154488
rect 238996 154476 239002 154488
rect 249058 154476 249064 154488
rect 238996 154448 249064 154476
rect 238996 154436 239002 154448
rect 249058 154436 249064 154448
rect 249116 154436 249122 154488
rect 249150 154436 249156 154488
rect 249208 154476 249214 154488
rect 249208 154448 297404 154476
rect 249208 154436 249214 154448
rect 48222 154368 48228 154420
rect 48280 154408 48286 154420
rect 155586 154408 155592 154420
rect 48280 154380 155592 154408
rect 48280 154368 48286 154380
rect 155586 154368 155592 154380
rect 155644 154368 155650 154420
rect 155770 154368 155776 154420
rect 155828 154408 155834 154420
rect 235258 154408 235264 154420
rect 155828 154380 232084 154408
rect 155828 154368 155834 154380
rect 41506 154300 41512 154352
rect 41564 154340 41570 154352
rect 150618 154340 150624 154352
rect 41564 154312 150624 154340
rect 41564 154300 41570 154312
rect 150618 154300 150624 154312
rect 150676 154300 150682 154352
rect 152366 154300 152372 154352
rect 152424 154340 152430 154352
rect 232056 154340 232084 154380
rect 233068 154380 235264 154408
rect 232958 154340 232964 154352
rect 152424 154312 231992 154340
rect 232056 154312 232964 154340
rect 152424 154300 152430 154312
rect 34790 154232 34796 154284
rect 34848 154272 34854 154284
rect 145558 154272 145564 154284
rect 34848 154244 145564 154272
rect 34848 154232 34854 154244
rect 145558 154232 145564 154244
rect 145616 154232 145622 154284
rect 145650 154232 145656 154284
rect 145708 154272 145714 154284
rect 230290 154272 230296 154284
rect 145708 154244 230296 154272
rect 145708 154232 145714 154244
rect 230290 154232 230296 154244
rect 230348 154232 230354 154284
rect 231964 154272 231992 154312
rect 232958 154300 232964 154312
rect 233016 154300 233022 154352
rect 233068 154272 233096 154380
rect 235258 154368 235264 154380
rect 235316 154368 235322 154420
rect 235350 154368 235356 154420
rect 235408 154408 235414 154420
rect 238110 154408 238116 154420
rect 235408 154380 238116 154408
rect 235408 154368 235414 154380
rect 238110 154368 238116 154380
rect 238168 154368 238174 154420
rect 238202 154368 238208 154420
rect 238260 154408 238266 154420
rect 240594 154408 240600 154420
rect 238260 154380 240600 154408
rect 238260 154368 238266 154380
rect 240594 154368 240600 154380
rect 240652 154368 240658 154420
rect 242158 154368 242164 154420
rect 242216 154408 242222 154420
rect 297376 154408 297404 154448
rect 299474 154436 299480 154488
rect 299532 154476 299538 154488
rect 306852 154476 306880 154516
rect 306926 154504 306932 154556
rect 306984 154544 306990 154556
rect 316402 154544 316408 154556
rect 306984 154516 316408 154544
rect 306984 154504 306990 154516
rect 316402 154504 316408 154516
rect 316460 154504 316466 154556
rect 316494 154504 316500 154556
rect 316552 154544 316558 154556
rect 360654 154544 360660 154556
rect 316552 154516 360660 154544
rect 316552 154504 316558 154516
rect 360654 154504 360660 154516
rect 360712 154504 360718 154556
rect 363874 154504 363880 154556
rect 363932 154544 363938 154556
rect 369578 154544 369584 154556
rect 363932 154516 369584 154544
rect 363932 154504 363938 154516
rect 369578 154504 369584 154516
rect 369636 154504 369642 154556
rect 369854 154504 369860 154556
rect 369912 154544 369918 154556
rect 401686 154544 401692 154556
rect 369912 154516 401692 154544
rect 369912 154504 369918 154516
rect 401686 154504 401692 154516
rect 401744 154504 401750 154556
rect 299532 154448 306788 154476
rect 306852 154448 307064 154476
rect 299532 154436 299538 154448
rect 306650 154408 306656 154420
rect 242216 154380 296024 154408
rect 297376 154380 306656 154408
rect 242216 154368 242222 154380
rect 233694 154300 233700 154352
rect 233752 154340 233758 154352
rect 236178 154340 236184 154352
rect 233752 154312 236184 154340
rect 233752 154300 233758 154312
rect 236178 154300 236184 154312
rect 236236 154300 236242 154352
rect 236362 154300 236368 154352
rect 236420 154340 236426 154352
rect 292666 154340 292672 154352
rect 236420 154312 292672 154340
rect 236420 154300 236426 154312
rect 292666 154300 292672 154312
rect 292724 154300 292730 154352
rect 295996 154340 296024 154380
rect 306650 154368 306656 154380
rect 306708 154368 306714 154420
rect 306760 154408 306788 154448
rect 306926 154408 306932 154420
rect 306760 154380 306932 154408
rect 306926 154368 306932 154380
rect 306984 154368 306990 154420
rect 307036 154408 307064 154448
rect 307110 154436 307116 154488
rect 307168 154476 307174 154488
rect 311434 154476 311440 154488
rect 307168 154448 311440 154476
rect 307168 154436 307174 154448
rect 311434 154436 311440 154448
rect 311492 154436 311498 154488
rect 312722 154436 312728 154488
rect 312780 154476 312786 154488
rect 358078 154476 358084 154488
rect 312780 154448 358084 154476
rect 312780 154436 312786 154448
rect 358078 154436 358084 154448
rect 358136 154436 358142 154488
rect 363138 154436 363144 154488
rect 363196 154476 363202 154488
rect 396534 154476 396540 154488
rect 363196 154448 396540 154476
rect 363196 154436 363202 154448
rect 396534 154436 396540 154448
rect 396592 154436 396598 154488
rect 403434 154436 403440 154488
rect 403492 154476 403498 154488
rect 427354 154476 427360 154488
rect 403492 154448 427360 154476
rect 403492 154436 403498 154448
rect 427354 154436 427360 154448
rect 427412 154436 427418 154488
rect 309226 154408 309232 154420
rect 307036 154380 309232 154408
rect 309226 154368 309232 154380
rect 309284 154368 309290 154420
rect 309410 154368 309416 154420
rect 309468 154408 309474 154420
rect 355502 154408 355508 154420
rect 309468 154380 355508 154408
rect 309468 154368 309474 154380
rect 355502 154368 355508 154380
rect 355560 154368 355566 154420
rect 358446 154368 358452 154420
rect 358504 154408 358510 154420
rect 359366 154408 359372 154420
rect 358504 154380 359372 154408
rect 358504 154368 358510 154380
rect 359366 154368 359372 154380
rect 359424 154368 359430 154420
rect 366450 154368 366456 154420
rect 366508 154408 366514 154420
rect 399110 154408 399116 154420
rect 366508 154380 399116 154408
rect 366508 154368 366514 154380
rect 399110 154368 399116 154380
rect 399168 154368 399174 154420
rect 400950 154368 400956 154420
rect 401008 154408 401014 154420
rect 425514 154408 425520 154420
rect 401008 154380 425520 154408
rect 401008 154368 401014 154380
rect 425514 154368 425520 154380
rect 425572 154368 425578 154420
rect 304074 154340 304080 154352
rect 295996 154312 304080 154340
rect 304074 154300 304080 154312
rect 304132 154300 304138 154352
rect 306006 154300 306012 154352
rect 306064 154340 306070 154352
rect 352834 154340 352840 154352
rect 306064 154312 352840 154340
rect 306064 154300 306070 154312
rect 352834 154300 352840 154312
rect 352892 154300 352898 154352
rect 358722 154340 358728 154352
rect 352990 154312 358728 154340
rect 231964 154244 233096 154272
rect 233142 154232 233148 154284
rect 233200 154272 233206 154284
rect 292298 154272 292304 154284
rect 233200 154244 292304 154272
rect 233200 154232 233206 154244
rect 292298 154232 292304 154244
rect 292356 154232 292362 154284
rect 295978 154232 295984 154284
rect 296036 154272 296042 154284
rect 336090 154272 336096 154284
rect 296036 154244 336096 154272
rect 296036 154232 296042 154244
rect 336090 154232 336096 154244
rect 336148 154232 336154 154284
rect 336182 154232 336188 154284
rect 336240 154272 336246 154284
rect 340138 154272 340144 154284
rect 336240 154244 340144 154272
rect 336240 154232 336246 154244
rect 340138 154232 340144 154244
rect 340196 154232 340202 154284
rect 340414 154232 340420 154284
rect 340472 154272 340478 154284
rect 345658 154272 345664 154284
rect 340472 154244 345664 154272
rect 340472 154232 340478 154244
rect 345658 154232 345664 154244
rect 345716 154232 345722 154284
rect 345750 154232 345756 154284
rect 345808 154272 345814 154284
rect 350350 154272 350356 154284
rect 345808 154244 350356 154272
rect 345808 154232 345814 154244
rect 350350 154232 350356 154244
rect 350408 154232 350414 154284
rect 38102 154164 38108 154216
rect 38160 154204 38166 154216
rect 148134 154204 148140 154216
rect 38160 154176 148140 154204
rect 38160 154164 38166 154176
rect 148134 154164 148140 154176
rect 148192 154164 148198 154216
rect 148962 154164 148968 154216
rect 149020 154204 149026 154216
rect 232866 154204 232872 154216
rect 149020 154176 232872 154204
rect 149020 154164 149026 154176
rect 232866 154164 232872 154176
rect 232924 154164 232930 154216
rect 232958 154164 232964 154216
rect 233016 154204 233022 154216
rect 235350 154204 235356 154216
rect 233016 154176 235356 154204
rect 233016 154164 233022 154176
rect 235350 154164 235356 154176
rect 235408 154164 235414 154216
rect 235442 154164 235448 154216
rect 235500 154204 235506 154216
rect 287146 154204 287152 154216
rect 235500 154176 287152 154204
rect 235500 154164 235506 154176
rect 287146 154164 287152 154176
rect 287204 154164 287210 154216
rect 287790 154164 287796 154216
rect 287848 154204 287854 154216
rect 292482 154204 292488 154216
rect 287848 154176 292488 154204
rect 287848 154164 287854 154176
rect 292482 154164 292488 154176
rect 292540 154164 292546 154216
rect 292942 154164 292948 154216
rect 293000 154204 293006 154216
rect 293000 154176 302234 154204
rect 293000 154164 293006 154176
rect 30558 154096 30564 154148
rect 30616 154136 30622 154148
rect 142338 154136 142344 154148
rect 30616 154108 142344 154136
rect 30616 154096 30622 154108
rect 142338 154096 142344 154108
rect 142396 154096 142402 154148
rect 142430 154096 142436 154148
rect 142488 154136 142494 154148
rect 227714 154136 227720 154148
rect 142488 154108 227720 154136
rect 142488 154096 142494 154108
rect 227714 154096 227720 154108
rect 227772 154096 227778 154148
rect 228726 154096 228732 154148
rect 228784 154136 228790 154148
rect 287606 154136 287612 154148
rect 228784 154108 287612 154136
rect 228784 154096 228790 154108
rect 287606 154096 287612 154108
rect 287664 154096 287670 154148
rect 291194 154096 291200 154148
rect 291252 154136 291258 154148
rect 297358 154136 297364 154148
rect 291252 154108 297364 154136
rect 291252 154096 291258 154108
rect 297358 154096 297364 154108
rect 297416 154096 297422 154148
rect 301590 154136 301596 154148
rect 299216 154108 301596 154136
rect 13814 154028 13820 154080
rect 13872 154068 13878 154080
rect 129458 154068 129464 154080
rect 13872 154040 129464 154068
rect 13872 154028 13878 154040
rect 129458 154028 129464 154040
rect 129516 154028 129522 154080
rect 129550 154028 129556 154080
rect 129608 154068 129614 154080
rect 217410 154068 217416 154080
rect 129608 154040 217416 154068
rect 129608 154028 129614 154040
rect 217410 154028 217416 154040
rect 217468 154028 217474 154080
rect 217502 154028 217508 154080
rect 217560 154068 217566 154080
rect 221918 154068 221924 154080
rect 217560 154040 221924 154068
rect 217560 154028 217566 154040
rect 221918 154028 221924 154040
rect 221976 154028 221982 154080
rect 222010 154028 222016 154080
rect 222068 154068 222074 154080
rect 225322 154068 225328 154080
rect 222068 154040 225328 154068
rect 222068 154028 222074 154040
rect 225322 154028 225328 154040
rect 225380 154028 225386 154080
rect 225414 154028 225420 154080
rect 225472 154068 225478 154080
rect 286962 154068 286968 154080
rect 225472 154040 286968 154068
rect 225472 154028 225478 154040
rect 286962 154028 286968 154040
rect 287020 154028 287026 154080
rect 287146 154028 287152 154080
rect 287204 154068 287210 154080
rect 292390 154068 292396 154080
rect 287204 154040 292396 154068
rect 287204 154028 287210 154040
rect 292390 154028 292396 154040
rect 292448 154028 292454 154080
rect 292666 154028 292672 154080
rect 292724 154068 292730 154080
rect 296438 154068 296444 154080
rect 292724 154040 296444 154068
rect 292724 154028 292730 154040
rect 296438 154028 296444 154040
rect 296496 154028 296502 154080
rect 297266 154028 297272 154080
rect 297324 154068 297330 154080
rect 299216 154068 299244 154108
rect 301590 154096 301596 154108
rect 301648 154096 301654 154148
rect 302206 154136 302234 154176
rect 302694 154164 302700 154216
rect 302752 154204 302758 154216
rect 342714 154204 342720 154216
rect 302752 154176 342720 154204
rect 302752 154164 302758 154176
rect 342714 154164 342720 154176
rect 342772 154164 342778 154216
rect 342806 154164 342812 154216
rect 342864 154204 342870 154216
rect 348510 154204 348516 154216
rect 342864 154176 348516 154204
rect 342864 154164 342870 154176
rect 348510 154164 348516 154176
rect 348568 154164 348574 154216
rect 351822 154164 351828 154216
rect 351880 154204 351886 154216
rect 352990 154204 353018 154312
rect 358722 154300 358728 154312
rect 358780 154300 358786 154352
rect 359734 154300 359740 154352
rect 359792 154340 359798 154352
rect 394050 154340 394056 154352
rect 359792 154312 394056 154340
rect 359792 154300 359798 154312
rect 394050 154300 394056 154312
rect 394108 154300 394114 154352
rect 400122 154300 400128 154352
rect 400180 154340 400186 154352
rect 424870 154340 424876 154352
rect 400180 154312 424876 154340
rect 400180 154300 400186 154312
rect 424870 154300 424876 154312
rect 424928 154300 424934 154352
rect 355318 154232 355324 154284
rect 355376 154272 355382 154284
rect 365714 154272 365720 154284
rect 355376 154244 365720 154272
rect 355376 154232 355382 154244
rect 365714 154232 365720 154244
rect 365772 154232 365778 154284
rect 393406 154232 393412 154284
rect 393464 154272 393470 154284
rect 419718 154272 419724 154284
rect 393464 154244 419724 154272
rect 393464 154232 393470 154244
rect 419718 154232 419724 154244
rect 419776 154232 419782 154284
rect 351880 154176 353018 154204
rect 351880 154164 351886 154176
rect 353110 154164 353116 154216
rect 353168 154204 353174 154216
rect 388898 154204 388904 154216
rect 353168 154176 388904 154204
rect 353168 154164 353174 154176
rect 388898 154164 388904 154176
rect 388956 154164 388962 154216
rect 396718 154164 396724 154216
rect 396776 154204 396782 154216
rect 422294 154204 422300 154216
rect 396776 154176 422300 154204
rect 396776 154164 396782 154176
rect 422294 154164 422300 154176
rect 422352 154164 422358 154216
rect 335998 154136 336004 154148
rect 302206 154108 336004 154136
rect 335998 154096 336004 154108
rect 336056 154096 336062 154148
rect 336090 154096 336096 154148
rect 336148 154136 336154 154148
rect 345198 154136 345204 154148
rect 336148 154108 345204 154136
rect 336148 154096 336154 154108
rect 345198 154096 345204 154108
rect 345256 154096 345262 154148
rect 346302 154096 346308 154148
rect 346360 154136 346366 154148
rect 383746 154136 383752 154148
rect 346360 154108 383752 154136
rect 346360 154096 346366 154108
rect 383746 154096 383752 154108
rect 383804 154096 383810 154148
rect 386598 154096 386604 154148
rect 386656 154136 386662 154148
rect 414566 154136 414572 154148
rect 386656 154108 414572 154136
rect 386656 154096 386662 154108
rect 414566 154096 414572 154108
rect 414624 154096 414630 154148
rect 417418 154096 417424 154148
rect 417476 154136 417482 154148
rect 432506 154136 432512 154148
rect 417476 154108 432512 154136
rect 417476 154096 417482 154108
rect 432506 154096 432512 154108
rect 432564 154096 432570 154148
rect 297324 154040 299244 154068
rect 297324 154028 297330 154040
rect 299290 154028 299296 154080
rect 299348 154068 299354 154080
rect 347774 154068 347780 154080
rect 299348 154040 347780 154068
rect 299348 154028 299354 154040
rect 347774 154028 347780 154040
rect 347832 154028 347838 154080
rect 349706 154028 349712 154080
rect 349764 154068 349770 154080
rect 386322 154068 386328 154080
rect 349764 154040 386328 154068
rect 349764 154028 349770 154040
rect 386322 154028 386328 154040
rect 386380 154028 386386 154080
rect 390002 154028 390008 154080
rect 390060 154068 390066 154080
rect 417142 154068 417148 154080
rect 390060 154040 417148 154068
rect 390060 154028 390066 154040
rect 417142 154028 417148 154040
rect 417200 154028 417206 154080
rect 427814 154028 427820 154080
rect 427872 154068 427878 154080
rect 446030 154068 446036 154080
rect 427872 154040 446036 154068
rect 427872 154028 427878 154040
rect 446030 154028 446036 154040
rect 446088 154028 446094 154080
rect 17126 153960 17132 154012
rect 17184 154000 17190 154012
rect 132034 154000 132040 154012
rect 17184 153972 132040 154000
rect 17184 153960 17190 153972
rect 132034 153960 132040 153972
rect 132092 153960 132098 154012
rect 132218 153960 132224 154012
rect 132276 154000 132282 154012
rect 219986 154000 219992 154012
rect 132276 153972 219992 154000
rect 132276 153960 132282 153972
rect 219986 153960 219992 153972
rect 220044 153960 220050 154012
rect 220722 153960 220728 154012
rect 220780 154000 220786 154012
rect 228266 154000 228272 154012
rect 220780 153972 228272 154000
rect 220780 153960 220786 153972
rect 228266 153960 228272 153972
rect 228324 153960 228330 154012
rect 228358 153960 228364 154012
rect 228416 154000 228422 154012
rect 288710 154000 288716 154012
rect 228416 153972 288716 154000
rect 228416 153960 228422 153972
rect 288710 153960 288716 153972
rect 288768 153960 288774 154012
rect 289262 153960 289268 154012
rect 289320 154000 289326 154012
rect 335906 154000 335912 154012
rect 289320 153972 335912 154000
rect 289320 153960 289326 153972
rect 335906 153960 335912 153972
rect 335964 153960 335970 154012
rect 335998 153960 336004 154012
rect 336056 154000 336062 154012
rect 342622 154000 342628 154012
rect 336056 153972 342628 154000
rect 336056 153960 336062 153972
rect 342622 153960 342628 153972
rect 342680 153960 342686 154012
rect 342990 153960 342996 154012
rect 343048 154000 343054 154012
rect 381170 154000 381176 154012
rect 343048 153972 381176 154000
rect 343048 153960 343054 153972
rect 381170 153960 381176 153972
rect 381228 153960 381234 154012
rect 383286 153960 383292 154012
rect 383344 154000 383350 154012
rect 411990 154000 411996 154012
rect 383344 153972 411996 154000
rect 383344 153960 383350 153972
rect 411990 153960 411996 153972
rect 412048 153960 412054 154012
rect 423582 153960 423588 154012
rect 423640 154000 423646 154012
rect 442810 154000 442816 154012
rect 423640 153972 442816 154000
rect 423640 153960 423646 153972
rect 442810 153960 442816 153972
rect 442868 153960 442874 154012
rect 4522 153892 4528 153944
rect 4580 153932 4586 153944
rect 122374 153932 122380 153944
rect 4580 153904 122380 153932
rect 4580 153892 4586 153904
rect 122374 153892 122380 153904
rect 122432 153892 122438 153944
rect 212258 153932 212264 153944
rect 122484 153904 212264 153932
rect 1210 153824 1216 153876
rect 1268 153864 1274 153876
rect 119798 153864 119804 153876
rect 1268 153836 119804 153864
rect 1268 153824 1274 153836
rect 119798 153824 119804 153836
rect 119856 153824 119862 153876
rect 122098 153824 122104 153876
rect 122156 153864 122162 153876
rect 122484 153864 122512 153904
rect 212258 153892 212264 153904
rect 212316 153892 212322 153944
rect 212810 153892 212816 153944
rect 212868 153932 212874 153944
rect 217502 153932 217508 153944
rect 212868 153904 217508 153932
rect 212868 153892 212874 153904
rect 217502 153892 217508 153904
rect 217560 153892 217566 153944
rect 217594 153892 217600 153944
rect 217652 153932 217658 153944
rect 280982 153932 280988 153944
rect 217652 153904 280988 153932
rect 217652 153892 217658 153904
rect 280982 153892 280988 153904
rect 281040 153892 281046 153944
rect 282546 153892 282552 153944
rect 282604 153932 282610 153944
rect 282604 153904 326200 153932
rect 282604 153892 282610 153904
rect 122156 153836 122512 153864
rect 122156 153824 122162 153836
rect 125502 153824 125508 153876
rect 125560 153864 125566 153876
rect 214834 153864 214840 153876
rect 125560 153836 214840 153864
rect 125560 153824 125566 153836
rect 214834 153824 214840 153836
rect 214892 153824 214898 153876
rect 215294 153824 215300 153876
rect 215352 153864 215358 153876
rect 217686 153864 217692 153876
rect 215352 153836 217692 153864
rect 215352 153824 215358 153836
rect 217686 153824 217692 153836
rect 217744 153824 217750 153876
rect 218698 153824 218704 153876
rect 218756 153864 218762 153876
rect 286134 153864 286140 153876
rect 218756 153836 286140 153864
rect 218756 153824 218762 153836
rect 286134 153824 286140 153836
rect 286192 153824 286198 153876
rect 286226 153824 286232 153876
rect 286284 153864 286290 153876
rect 326062 153864 326068 153876
rect 286284 153836 326068 153864
rect 286284 153824 286290 153836
rect 326062 153824 326068 153836
rect 326120 153824 326126 153876
rect 58250 153756 58256 153808
rect 58308 153796 58314 153808
rect 163498 153796 163504 153808
rect 58308 153768 163504 153796
rect 58308 153756 58314 153768
rect 163498 153756 163504 153768
rect 163556 153756 163562 153808
rect 165798 153756 165804 153808
rect 165856 153796 165862 153808
rect 245654 153796 245660 153808
rect 165856 153768 245660 153796
rect 165856 153756 165862 153768
rect 245654 153756 245660 153768
rect 245712 153756 245718 153808
rect 246960 153768 252232 153796
rect 68370 153688 68376 153740
rect 68428 153728 68434 153740
rect 171226 153728 171232 153740
rect 68428 153700 171232 153728
rect 68428 153688 68434 153700
rect 171226 153688 171232 153700
rect 171284 153688 171290 153740
rect 175734 153688 175740 153740
rect 175792 153728 175798 153740
rect 246960 153728 246988 153768
rect 248230 153728 248236 153740
rect 175792 153700 246988 153728
rect 247052 153700 248236 153728
rect 175792 153688 175798 153700
rect 64966 153620 64972 153672
rect 65024 153660 65030 153672
rect 168650 153660 168656 153672
rect 65024 153632 168656 153660
rect 65024 153620 65030 153632
rect 168650 153620 168656 153632
rect 168708 153620 168714 153672
rect 169110 153620 169116 153672
rect 169168 153660 169174 153672
rect 247052 153660 247080 153700
rect 248230 153688 248236 153700
rect 248288 153688 248294 153740
rect 252204 153728 252232 153768
rect 252278 153756 252284 153808
rect 252336 153796 252342 153808
rect 306926 153796 306932 153808
rect 252336 153768 306932 153796
rect 252336 153756 252342 153768
rect 306926 153756 306932 153768
rect 306984 153756 306990 153808
rect 307018 153756 307024 153808
rect 307076 153796 307082 153808
rect 325326 153796 325332 153808
rect 307076 153768 325332 153796
rect 307076 153756 307082 153768
rect 325326 153756 325332 153768
rect 325384 153756 325390 153808
rect 326172 153796 326200 153904
rect 326246 153892 326252 153944
rect 326304 153932 326310 153944
rect 326304 153904 336228 153932
rect 326304 153892 326310 153904
rect 326430 153824 326436 153876
rect 326488 153864 326494 153876
rect 335538 153864 335544 153876
rect 326488 153836 335544 153864
rect 326488 153824 326494 153836
rect 335538 153824 335544 153836
rect 335596 153824 335602 153876
rect 336200 153864 336228 153904
rect 336274 153892 336280 153944
rect 336332 153932 336338 153944
rect 376018 153932 376024 153944
rect 336332 153904 376024 153932
rect 336332 153892 336338 153904
rect 376018 153892 376024 153904
rect 376076 153892 376082 153944
rect 376570 153892 376576 153944
rect 376628 153932 376634 153944
rect 406838 153932 406844 153944
rect 376628 153904 406844 153932
rect 376628 153892 376634 153904
rect 406838 153892 406844 153904
rect 406896 153892 406902 153944
rect 407666 153892 407672 153944
rect 407724 153932 407730 153944
rect 430482 153932 430488 153944
rect 407724 153904 430488 153932
rect 407724 153892 407730 153904
rect 430482 153892 430488 153904
rect 430540 153892 430546 153944
rect 430574 153892 430580 153944
rect 430632 153932 430638 153944
rect 440878 153932 440884 153944
rect 430632 153904 440884 153932
rect 430632 153892 430638 153904
rect 440878 153892 440884 153904
rect 440936 153892 440942 153944
rect 337470 153864 337476 153876
rect 336200 153836 337476 153864
rect 337470 153824 337476 153836
rect 337528 153824 337534 153876
rect 339586 153824 339592 153876
rect 339644 153864 339650 153876
rect 378594 153864 378600 153876
rect 339644 153836 378600 153864
rect 339644 153824 339650 153836
rect 378594 153824 378600 153836
rect 378652 153824 378658 153876
rect 379882 153824 379888 153876
rect 379940 153864 379946 153876
rect 409414 153864 409420 153876
rect 379940 153836 409420 153864
rect 379940 153824 379946 153836
rect 409414 153824 409420 153836
rect 409472 153824 409478 153876
rect 416866 153824 416872 153876
rect 416924 153864 416930 153876
rect 437658 153864 437664 153876
rect 416924 153836 437664 153864
rect 416924 153824 416930 153836
rect 437658 153824 437664 153836
rect 437716 153824 437722 153876
rect 326522 153796 326528 153808
rect 326172 153768 326528 153796
rect 326522 153756 326528 153768
rect 326580 153756 326586 153808
rect 326614 153756 326620 153808
rect 326672 153796 326678 153808
rect 350718 153796 350724 153808
rect 326672 153768 350724 153796
rect 326672 153756 326678 153768
rect 350718 153756 350724 153768
rect 350776 153756 350782 153808
rect 363230 153796 363236 153808
rect 350828 153768 363236 153796
rect 253382 153728 253388 153740
rect 252204 153700 253388 153728
rect 253382 153688 253388 153700
rect 253440 153688 253446 153740
rect 255590 153688 255596 153740
rect 255648 153728 255654 153740
rect 311710 153728 311716 153740
rect 255648 153700 311716 153728
rect 255648 153688 255654 153700
rect 311710 153688 311716 153700
rect 311768 153688 311774 153740
rect 311802 153688 311808 153740
rect 311860 153728 311866 153740
rect 312354 153728 312360 153740
rect 311860 153700 312360 153728
rect 311860 153688 311866 153700
rect 312354 153688 312360 153700
rect 312412 153688 312418 153740
rect 312722 153688 312728 153740
rect 312780 153728 312786 153740
rect 324682 153728 324688 153740
rect 312780 153700 324688 153728
rect 312780 153688 312786 153700
rect 324682 153688 324688 153700
rect 324740 153688 324746 153740
rect 326338 153688 326344 153740
rect 326396 153728 326402 153740
rect 350828 153728 350856 153768
rect 363230 153756 363236 153768
rect 363288 153756 363294 153808
rect 367094 153756 367100 153808
rect 367152 153796 367158 153808
rect 372154 153796 372160 153808
rect 367152 153768 372160 153796
rect 367152 153756 367158 153768
rect 372154 153756 372160 153768
rect 372212 153756 372218 153808
rect 373166 153756 373172 153808
rect 373224 153796 373230 153808
rect 404262 153796 404268 153808
rect 373224 153768 404268 153796
rect 373224 153756 373230 153768
rect 404262 153756 404268 153768
rect 404320 153756 404326 153808
rect 326396 153700 350856 153728
rect 326396 153688 326402 153700
rect 350902 153688 350908 153740
rect 350960 153728 350966 153740
rect 355318 153728 355324 153740
rect 350960 153700 355324 153728
rect 350960 153688 350966 153700
rect 355318 153688 355324 153700
rect 355376 153688 355382 153740
rect 357434 153688 357440 153740
rect 357492 153728 357498 153740
rect 368934 153728 368940 153740
rect 357492 153700 368940 153728
rect 357492 153688 357498 153700
rect 368934 153688 368940 153700
rect 368992 153688 368998 153740
rect 169168 153632 247080 153660
rect 169168 153620 169174 153632
rect 247126 153620 247132 153672
rect 247184 153660 247190 153672
rect 256510 153660 256516 153672
rect 247184 153632 256516 153660
rect 247184 153620 247190 153632
rect 256510 153620 256516 153632
rect 256568 153620 256574 153672
rect 258994 153620 259000 153672
rect 259052 153660 259058 153672
rect 316310 153660 316316 153672
rect 259052 153632 316316 153660
rect 259052 153620 259058 153632
rect 316310 153620 316316 153632
rect 316368 153620 316374 153672
rect 316402 153620 316408 153672
rect 316460 153660 316466 153672
rect 327902 153660 327908 153672
rect 316460 153632 327908 153660
rect 316460 153620 316466 153632
rect 327902 153620 327908 153632
rect 327960 153620 327966 153672
rect 329558 153620 329564 153672
rect 329616 153660 329622 153672
rect 370866 153660 370872 153672
rect 329616 153632 370872 153660
rect 329616 153620 329622 153632
rect 370866 153620 370872 153632
rect 370924 153620 370930 153672
rect 8754 153552 8760 153604
rect 8812 153592 8818 153604
rect 109034 153592 109040 153604
rect 8812 153564 109040 153592
rect 8812 153552 8818 153564
rect 109034 153552 109040 153564
rect 109092 153552 109098 153604
rect 112070 153552 112076 153604
rect 112128 153592 112134 153604
rect 204622 153592 204628 153604
rect 112128 153564 204628 153592
rect 112128 153552 112134 153564
rect 204622 153552 204628 153564
rect 204680 153552 204686 153604
rect 208578 153552 208584 153604
rect 208636 153592 208642 153604
rect 278406 153592 278412 153604
rect 208636 153564 278412 153592
rect 208636 153552 208642 153564
rect 278406 153552 278412 153564
rect 278464 153552 278470 153604
rect 279142 153552 279148 153604
rect 279200 153592 279206 153604
rect 332410 153592 332416 153604
rect 279200 153564 312492 153592
rect 279200 153552 279206 153564
rect 75086 153484 75092 153536
rect 75144 153524 75150 153536
rect 176378 153524 176384 153536
rect 75144 153496 176384 153524
rect 75144 153484 75150 153496
rect 176378 153484 176384 153496
rect 176436 153484 176442 153536
rect 182542 153484 182548 153536
rect 182600 153524 182606 153536
rect 258534 153524 258540 153536
rect 182600 153496 258540 153524
rect 182600 153484 182606 153496
rect 258534 153484 258540 153496
rect 258592 153484 258598 153536
rect 269114 153484 269120 153536
rect 269172 153524 269178 153536
rect 312354 153524 312360 153536
rect 269172 153496 312360 153524
rect 269172 153484 269178 153496
rect 312354 153484 312360 153496
rect 312412 153484 312418 153536
rect 312464 153524 312492 153564
rect 312648 153564 332416 153592
rect 312648 153524 312676 153564
rect 332410 153552 332416 153564
rect 332468 153552 332474 153604
rect 332870 153552 332876 153604
rect 332928 153592 332934 153604
rect 373442 153592 373448 153604
rect 332928 153564 373448 153592
rect 332928 153552 332934 153564
rect 373442 153552 373448 153564
rect 373500 153552 373506 153604
rect 322750 153524 322756 153536
rect 312464 153496 312676 153524
rect 312740 153496 322756 153524
rect 27246 153416 27252 153468
rect 27304 153456 27310 153468
rect 125686 153456 125692 153468
rect 27304 153428 125692 153456
rect 27304 153416 27310 153428
rect 125686 153416 125692 153428
rect 125744 153416 125750 153468
rect 135530 153416 135536 153468
rect 135588 153456 135594 153468
rect 222562 153456 222568 153468
rect 135588 153428 222568 153456
rect 135588 153416 135594 153428
rect 222562 153416 222568 153428
rect 222620 153416 222626 153468
rect 225322 153416 225328 153468
rect 225380 153456 225386 153468
rect 228358 153456 228364 153468
rect 225380 153428 228364 153456
rect 225380 153416 225386 153428
rect 228358 153416 228364 153428
rect 228416 153416 228422 153468
rect 228450 153416 228456 153468
rect 228508 153456 228514 153468
rect 236086 153456 236092 153468
rect 228508 153428 236092 153456
rect 228508 153416 228514 153428
rect 236086 153416 236092 153428
rect 236144 153416 236150 153468
rect 236178 153416 236184 153468
rect 236236 153456 236242 153468
rect 241238 153456 241244 153468
rect 236236 153428 241244 153456
rect 236236 153416 236242 153428
rect 241238 153416 241244 153428
rect 241296 153416 241302 153468
rect 241422 153416 241428 153468
rect 241480 153456 241486 153468
rect 246298 153456 246304 153468
rect 241480 153428 246304 153456
rect 241480 153416 241486 153428
rect 246298 153416 246304 153428
rect 246356 153416 246362 153468
rect 249058 153416 249064 153468
rect 249116 153456 249122 153468
rect 297266 153456 297272 153468
rect 249116 153428 297272 153456
rect 249116 153416 249122 153428
rect 297266 153416 297272 153428
rect 297324 153416 297330 153468
rect 297358 153416 297364 153468
rect 297416 153456 297422 153468
rect 312740 153456 312768 153496
rect 322750 153484 322756 153496
rect 322808 153484 322814 153536
rect 322842 153484 322848 153536
rect 322900 153524 322906 153536
rect 326614 153524 326620 153536
rect 322900 153496 326620 153524
rect 322900 153484 322906 153496
rect 326614 153484 326620 153496
rect 326672 153484 326678 153536
rect 364886 153524 364892 153536
rect 327460 153496 364892 153524
rect 327258 153456 327264 153468
rect 297416 153428 312768 153456
rect 312832 153428 327264 153456
rect 297416 153416 297422 153428
rect 85114 153348 85120 153400
rect 85172 153388 85178 153400
rect 184014 153388 184020 153400
rect 85172 153360 184020 153388
rect 85172 153348 85178 153360
rect 184014 153348 184020 153360
rect 184072 153348 184078 153400
rect 184842 153348 184848 153400
rect 184900 153388 184906 153400
rect 184900 153360 188660 153388
rect 184900 153348 184906 153360
rect 88518 153280 88524 153332
rect 88576 153320 88582 153332
rect 186590 153320 186596 153332
rect 88576 153292 186596 153320
rect 88576 153280 88582 153292
rect 186590 153280 186596 153292
rect 186648 153280 186654 153332
rect 188632 153320 188660 153360
rect 189258 153348 189264 153400
rect 189316 153388 189322 153400
rect 263686 153388 263692 153400
rect 189316 153360 263692 153388
rect 189316 153348 189322 153360
rect 263686 153348 263692 153360
rect 263744 153348 263750 153400
rect 272426 153348 272432 153400
rect 272484 153388 272490 153400
rect 312832 153388 312860 153428
rect 327258 153416 327264 153428
rect 327316 153416 327322 153468
rect 272484 153360 312860 153388
rect 272484 153348 272490 153360
rect 312906 153348 312912 153400
rect 312964 153388 312970 153400
rect 317598 153388 317604 153400
rect 312964 153360 317604 153388
rect 312964 153348 312970 153360
rect 317598 153348 317604 153360
rect 317656 153348 317662 153400
rect 317782 153348 317788 153400
rect 317840 153388 317846 153400
rect 319346 153388 319352 153400
rect 317840 153360 319352 153388
rect 317840 153348 317846 153360
rect 319346 153348 319352 153360
rect 319404 153348 319410 153400
rect 319438 153348 319444 153400
rect 319496 153388 319502 153400
rect 326338 153388 326344 153400
rect 319496 153360 326344 153388
rect 319496 153348 319502 153360
rect 326338 153348 326344 153360
rect 326396 153348 326402 153400
rect 326706 153348 326712 153400
rect 326764 153388 326770 153400
rect 327460 153388 327488 153496
rect 364886 153484 364892 153496
rect 364944 153484 364950 153536
rect 376662 153524 376668 153536
rect 365088 153496 376668 153524
rect 327626 153416 327632 153468
rect 327684 153456 327690 153468
rect 327684 153428 343404 153456
rect 327684 153416 327690 153428
rect 326764 153360 327488 153388
rect 326764 153348 326770 153360
rect 327534 153348 327540 153400
rect 327592 153388 327598 153400
rect 331398 153388 331404 153400
rect 327592 153360 331404 153388
rect 327592 153348 327598 153360
rect 331398 153348 331404 153360
rect 331456 153348 331462 153400
rect 334894 153388 334900 153400
rect 331508 153360 334900 153388
rect 212902 153320 212908 153332
rect 188632 153292 212908 153320
rect 212902 153280 212908 153292
rect 212960 153280 212966 153332
rect 212994 153280 213000 153332
rect 213052 153320 213058 153332
rect 217594 153320 217600 153332
rect 213052 153292 217600 153320
rect 213052 153280 213058 153292
rect 217594 153280 217600 153292
rect 217652 153280 217658 153332
rect 217686 153280 217692 153332
rect 217744 153320 217750 153332
rect 217744 153292 220860 153320
rect 217744 153280 217750 153292
rect 105354 153212 105360 153264
rect 105412 153252 105418 153264
rect 199470 153252 199476 153264
rect 105412 153224 199476 153252
rect 105412 153212 105418 153224
rect 199470 153212 199476 153224
rect 199528 153212 199534 153264
rect 200482 153212 200488 153264
rect 200540 153252 200546 153264
rect 220722 153252 220728 153264
rect 200540 153224 220728 153252
rect 200540 153212 200546 153224
rect 220722 153212 220728 153224
rect 220780 153212 220786 153264
rect 220832 153252 220860 153292
rect 221918 153280 221924 153332
rect 221976 153320 221982 153332
rect 281626 153320 281632 153332
rect 221976 153292 281632 153320
rect 221976 153280 221982 153292
rect 281626 153280 281632 153292
rect 281684 153280 281690 153332
rect 283006 153280 283012 153332
rect 283064 153320 283070 153332
rect 286870 153320 286876 153332
rect 283064 153292 286876 153320
rect 283064 153280 283070 153292
rect 286870 153280 286876 153292
rect 286928 153280 286934 153332
rect 286962 153280 286968 153332
rect 287020 153320 287026 153332
rect 291286 153320 291292 153332
rect 287020 153292 291292 153320
rect 287020 153280 287026 153292
rect 291286 153280 291292 153292
rect 291344 153280 291350 153332
rect 326430 153320 326436 153332
rect 291396 153292 326436 153320
rect 283558 153252 283564 153264
rect 220832 153224 283564 153252
rect 283558 153212 283564 153224
rect 283616 153212 283622 153264
rect 284294 153212 284300 153264
rect 284352 153252 284358 153264
rect 291396 153252 291424 153292
rect 326430 153280 326436 153292
rect 326488 153280 326494 153332
rect 326522 153280 326528 153332
rect 326580 153320 326586 153332
rect 331508 153320 331536 153360
rect 334894 153348 334900 153360
rect 334952 153348 334958 153400
rect 335262 153348 335268 153400
rect 335320 153388 335326 153400
rect 337010 153388 337016 153400
rect 335320 153360 337016 153388
rect 335320 153348 335326 153360
rect 337010 153348 337016 153360
rect 337068 153348 337074 153400
rect 337102 153348 337108 153400
rect 337160 153388 337166 153400
rect 342898 153388 342904 153400
rect 337160 153360 342904 153388
rect 337160 153348 337166 153360
rect 342898 153348 342904 153360
rect 342956 153348 342962 153400
rect 326580 153292 331536 153320
rect 326580 153280 326586 153292
rect 331582 153280 331588 153332
rect 331640 153320 331646 153332
rect 343266 153320 343272 153332
rect 331640 153292 343272 153320
rect 331640 153280 331646 153292
rect 343266 153280 343272 153292
rect 343324 153280 343330 153332
rect 343376 153320 343404 153428
rect 345658 153416 345664 153468
rect 345716 153456 345722 153468
rect 364978 153456 364984 153468
rect 345716 153428 364984 153456
rect 345716 153416 345722 153428
rect 364978 153416 364984 153428
rect 365036 153416 365042 153468
rect 345382 153348 345388 153400
rect 345440 153388 345446 153400
rect 365088 153388 365116 153496
rect 376662 153484 376668 153496
rect 376720 153484 376726 153536
rect 365162 153416 365168 153468
rect 365220 153456 365226 153468
rect 379238 153456 379244 153468
rect 365220 153428 379244 153456
rect 365220 153416 365226 153428
rect 379238 153416 379244 153428
rect 379296 153416 379302 153468
rect 345440 153360 365116 153388
rect 345440 153348 345446 153360
rect 368474 153348 368480 153400
rect 368532 153388 368538 153400
rect 374730 153388 374736 153400
rect 368532 153360 374736 153388
rect 368532 153348 368538 153360
rect 374730 153348 374736 153360
rect 374788 153348 374794 153400
rect 348418 153320 348424 153332
rect 343376 153292 348424 153320
rect 348418 153280 348424 153292
rect 348476 153280 348482 153332
rect 348510 153280 348516 153332
rect 348568 153320 348574 153332
rect 356146 153320 356152 153332
rect 348568 153292 356152 153320
rect 348568 153280 348574 153292
rect 356146 153280 356152 153292
rect 356204 153280 356210 153332
rect 363874 153320 363880 153332
rect 356256 153292 363880 153320
rect 284352 153224 291424 153252
rect 284352 153212 284358 153224
rect 291470 153212 291476 153264
rect 291528 153252 291534 153264
rect 311802 153252 311808 153264
rect 291528 153224 311808 153252
rect 291528 153212 291534 153224
rect 311802 153212 311808 153224
rect 311860 153212 311866 153264
rect 311894 153212 311900 153264
rect 311952 153252 311958 153264
rect 314378 153252 314384 153264
rect 311952 153224 314384 153252
rect 311952 153212 311958 153224
rect 314378 153212 314384 153224
rect 314436 153212 314442 153264
rect 314562 153212 314568 153264
rect 314620 153252 314626 153264
rect 316218 153252 316224 153264
rect 314620 153224 316224 153252
rect 314620 153212 314626 153224
rect 316218 153212 316224 153224
rect 316276 153212 316282 153264
rect 316310 153212 316316 153264
rect 316368 153252 316374 153264
rect 316954 153252 316960 153264
rect 316368 153224 316960 153252
rect 316368 153212 316374 153224
rect 316954 153212 316960 153224
rect 317012 153212 317018 153264
rect 317138 153212 317144 153264
rect 317196 153252 317202 153264
rect 333054 153252 333060 153264
rect 317196 153224 333060 153252
rect 317196 153212 317202 153224
rect 333054 153212 333060 153224
rect 333112 153212 333118 153264
rect 335906 153212 335912 153264
rect 335964 153252 335970 153264
rect 340046 153252 340052 153264
rect 335964 153224 340052 153252
rect 335964 153212 335970 153224
rect 340046 153212 340052 153224
rect 340104 153212 340110 153264
rect 340138 153212 340144 153264
rect 340196 153252 340202 153264
rect 353570 153252 353576 153264
rect 340196 153224 353576 153252
rect 340196 153212 340202 153224
rect 353570 153212 353576 153224
rect 353628 153212 353634 153264
rect 355226 153212 355232 153264
rect 355284 153252 355290 153264
rect 356256 153252 356284 153292
rect 363874 153280 363880 153292
rect 363932 153280 363938 153332
rect 364886 153280 364892 153332
rect 364944 153320 364950 153332
rect 368290 153320 368296 153332
rect 364944 153292 368296 153320
rect 364944 153280 364950 153292
rect 368290 153280 368296 153292
rect 368348 153280 368354 153332
rect 355284 153224 356284 153252
rect 355284 153212 355290 153224
rect 356422 153212 356428 153264
rect 356480 153252 356486 153264
rect 391474 153252 391480 153264
rect 356480 153224 391480 153252
rect 356480 153212 356486 153224
rect 391474 153212 391480 153224
rect 391532 153212 391538 153264
rect 437474 153212 437480 153264
rect 437532 153252 437538 153264
rect 443454 153252 443460 153264
rect 437532 153224 443460 153252
rect 437532 153212 437538 153224
rect 443454 153212 443460 153224
rect 443512 153212 443518 153264
rect 80146 153144 80152 153196
rect 80204 153184 80210 153196
rect 180242 153184 180248 153196
rect 80204 153156 180248 153184
rect 80204 153144 80210 153156
rect 180242 153144 180248 153156
rect 180300 153144 180306 153196
rect 183278 153144 183284 153196
rect 183336 153184 183342 153196
rect 187878 153184 187884 153196
rect 183336 153156 187884 153184
rect 183336 153144 183342 153156
rect 187878 153144 187884 153156
rect 187936 153144 187942 153196
rect 190086 153144 190092 153196
rect 190144 153184 190150 153196
rect 264422 153184 264428 153196
rect 190144 153156 264428 153184
rect 190144 153144 190150 153156
rect 264422 153144 264428 153156
rect 264480 153144 264486 153196
rect 264514 153144 264520 153196
rect 264572 153184 264578 153196
rect 315666 153184 315672 153196
rect 264572 153156 315672 153184
rect 264572 153144 264578 153156
rect 315666 153144 315672 153156
rect 315724 153144 315730 153196
rect 315942 153144 315948 153196
rect 316000 153184 316006 153196
rect 318242 153184 318248 153196
rect 316000 153156 318248 153184
rect 316000 153144 316006 153156
rect 318242 153144 318248 153156
rect 318300 153144 318306 153196
rect 318610 153144 318616 153196
rect 318668 153184 318674 153196
rect 362586 153184 362592 153196
rect 318668 153156 362592 153184
rect 318668 153144 318674 153156
rect 362586 153144 362592 153156
rect 362644 153144 362650 153196
rect 365622 153144 365628 153196
rect 365680 153184 365686 153196
rect 398466 153184 398472 153196
rect 365680 153156 398472 153184
rect 365680 153144 365686 153156
rect 398466 153144 398472 153156
rect 398524 153144 398530 153196
rect 404170 153144 404176 153196
rect 404228 153184 404234 153196
rect 418430 153184 418436 153196
rect 404228 153156 418436 153184
rect 404228 153144 404234 153156
rect 418430 153144 418436 153156
rect 418488 153144 418494 153196
rect 418522 153144 418528 153196
rect 418580 153184 418586 153196
rect 438946 153184 438952 153196
rect 418580 153156 438952 153184
rect 418580 153144 418586 153156
rect 438946 153144 438952 153156
rect 439004 153144 439010 153196
rect 448514 153144 448520 153196
rect 448572 153184 448578 153196
rect 451182 153184 451188 153196
rect 448572 153156 451188 153184
rect 448572 153144 448578 153156
rect 451182 153144 451188 153156
rect 451240 153144 451246 153196
rect 451274 153144 451280 153196
rect 451332 153184 451338 153196
rect 453114 153184 453120 153196
rect 451332 153156 453120 153184
rect 451332 153144 451338 153156
rect 453114 153144 453120 153156
rect 453172 153144 453178 153196
rect 458174 153144 458180 153196
rect 458232 153184 458238 153196
rect 460750 153184 460756 153196
rect 458232 153156 460756 153184
rect 458232 153144 458238 153156
rect 460750 153144 460756 153156
rect 460808 153144 460814 153196
rect 473078 153144 473084 153196
rect 473136 153184 473142 153196
rect 475562 153184 475568 153196
rect 473136 153156 475568 153184
rect 473136 153144 473142 153156
rect 475562 153144 475568 153156
rect 475620 153144 475626 153196
rect 477402 153144 477408 153196
rect 477460 153184 477466 153196
rect 478782 153184 478788 153196
rect 477460 153156 478788 153184
rect 477460 153144 477466 153156
rect 478782 153144 478788 153156
rect 478840 153144 478846 153196
rect 480806 153144 480812 153196
rect 480864 153184 480870 153196
rect 482002 153184 482008 153196
rect 480864 153156 482008 153184
rect 480864 153144 480870 153156
rect 482002 153144 482008 153156
rect 482060 153144 482066 153196
rect 490374 153144 490380 153196
rect 490432 153184 490438 153196
rect 492214 153184 492220 153196
rect 490432 153156 492220 153184
rect 490432 153144 490438 153156
rect 492214 153144 492220 153156
rect 492272 153144 492278 153196
rect 73430 153076 73436 153128
rect 73488 153116 73494 153128
rect 175090 153116 175096 153128
rect 73488 153088 175096 153116
rect 73488 153076 73494 153088
rect 175090 153076 175096 153088
rect 175148 153076 175154 153128
rect 176654 153076 176660 153128
rect 176712 153116 176718 153128
rect 176712 153088 185624 153116
rect 176712 153076 176718 153088
rect 63310 153008 63316 153060
rect 63368 153048 63374 153060
rect 167362 153048 167368 153060
rect 63368 153020 167368 153048
rect 63368 153008 63374 153020
rect 167362 153008 167368 153020
rect 167420 153008 167426 153060
rect 169754 153008 169760 153060
rect 169812 153048 169818 153060
rect 177666 153048 177672 153060
rect 169812 153020 177672 153048
rect 169812 153008 169818 153020
rect 177666 153008 177672 153020
rect 177724 153008 177730 153060
rect 177758 153008 177764 153060
rect 177816 153048 177822 153060
rect 182726 153048 182732 153060
rect 177816 153020 182732 153048
rect 177816 153008 177822 153020
rect 182726 153008 182732 153020
rect 182784 153008 182790 153060
rect 185596 153048 185624 153088
rect 186130 153076 186136 153128
rect 186188 153116 186194 153128
rect 259822 153116 259828 153128
rect 186188 153088 259828 153116
rect 186188 153076 186194 153088
rect 259822 153076 259828 153088
rect 259880 153076 259886 153128
rect 260190 153076 260196 153128
rect 260248 153116 260254 153128
rect 266906 153116 266912 153128
rect 260248 153088 266912 153116
rect 260248 153076 260254 153088
rect 266906 153076 266912 153088
rect 266964 153076 266970 153128
rect 271874 153076 271880 153128
rect 271932 153116 271938 153128
rect 271932 153088 274496 153116
rect 271932 153076 271938 153088
rect 254026 153048 254032 153060
rect 185596 153020 254032 153048
rect 254026 153008 254032 153020
rect 254084 153008 254090 153060
rect 254118 153008 254124 153060
rect 254176 153048 254182 153060
rect 261754 153048 261760 153060
rect 254176 153020 261760 153048
rect 254176 153008 254182 153020
rect 261754 153008 261760 153020
rect 261812 153008 261818 153060
rect 263594 153008 263600 153060
rect 263652 153048 263658 153060
rect 272058 153048 272064 153060
rect 263652 153020 272064 153048
rect 263652 153008 263658 153020
rect 272058 153008 272064 153020
rect 272116 153008 272122 153060
rect 274468 153048 274496 153088
rect 276658 153076 276664 153128
rect 276716 153116 276722 153128
rect 330478 153116 330484 153128
rect 276716 153088 330484 153116
rect 276716 153076 276722 153088
rect 330478 153076 330484 153088
rect 330536 153076 330542 153128
rect 330754 153076 330760 153128
rect 330812 153116 330818 153128
rect 371510 153116 371516 153128
rect 330812 153088 371516 153116
rect 330812 153076 330818 153088
rect 371510 153076 371516 153088
rect 371568 153076 371574 153128
rect 377398 153076 377404 153128
rect 377456 153116 377462 153128
rect 407482 153116 407488 153128
rect 377456 153088 407488 153116
rect 377456 153076 377462 153088
rect 407482 153076 407488 153088
rect 407540 153076 407546 153128
rect 414382 153076 414388 153128
rect 414440 153116 414446 153128
rect 435726 153116 435732 153128
rect 414440 153088 435732 153116
rect 414440 153076 414446 153088
rect 435726 153076 435732 153088
rect 435784 153076 435790 153128
rect 447226 153076 447232 153128
rect 447284 153116 447290 153128
rect 449250 153116 449256 153128
rect 447284 153088 449256 153116
rect 447284 153076 447290 153088
rect 449250 153076 449256 153088
rect 449308 153076 449314 153128
rect 452838 153076 452844 153128
rect 452896 153116 452902 153128
rect 454402 153116 454408 153128
rect 452896 153088 454408 153116
rect 452896 153076 452902 153088
rect 454402 153076 454408 153088
rect 454460 153076 454466 153128
rect 473630 153076 473636 153128
rect 473688 153116 473694 153128
rect 476942 153116 476948 153128
rect 473688 153088 476948 153116
rect 473688 153076 473694 153088
rect 476942 153076 476948 153088
rect 477000 153076 477006 153128
rect 481726 153076 481732 153128
rect 481784 153116 481790 153128
rect 483934 153116 483940 153128
rect 481784 153088 483940 153116
rect 481784 153076 481790 153088
rect 483934 153076 483940 153088
rect 483992 153076 483998 153128
rect 326614 153048 326620 153060
rect 274468 153020 326620 153048
rect 326614 153008 326620 153020
rect 326672 153008 326678 153060
rect 367646 153048 367652 153060
rect 326724 153020 367652 153048
rect 56594 152940 56600 152992
rect 56652 152980 56658 152992
rect 162210 152980 162216 152992
rect 56652 152952 162216 152980
rect 56652 152940 56658 152952
rect 162210 152940 162216 152952
rect 162268 152940 162274 152992
rect 169938 152940 169944 152992
rect 169996 152980 170002 152992
rect 248874 152980 248880 152992
rect 169996 152952 248880 152980
rect 169996 152940 170002 152952
rect 248874 152940 248880 152952
rect 248932 152940 248938 152992
rect 250622 152940 250628 152992
rect 250680 152980 250686 152992
rect 254302 152980 254308 152992
rect 250680 152952 254308 152980
rect 250680 152940 250686 152952
rect 254302 152940 254308 152952
rect 254360 152940 254366 152992
rect 266722 152940 266728 152992
rect 266780 152980 266786 152992
rect 320818 152980 320824 152992
rect 266780 152952 320824 152980
rect 266780 152940 266786 152952
rect 320818 152940 320824 152952
rect 320876 152940 320882 152992
rect 321554 152940 321560 152992
rect 321612 152980 321618 152992
rect 324038 152980 324044 152992
rect 321612 152952 324044 152980
rect 321612 152940 321618 152952
rect 324038 152940 324044 152952
rect 324096 152940 324102 152992
rect 325694 152940 325700 152992
rect 325752 152980 325758 152992
rect 326724 152980 326752 153020
rect 367646 153008 367652 153020
rect 367704 153008 367710 153060
rect 370682 153008 370688 153060
rect 370740 153048 370746 153060
rect 402330 153048 402336 153060
rect 370740 153020 402336 153048
rect 370740 153008 370746 153020
rect 402330 153008 402336 153020
rect 402388 153008 402394 153060
rect 413922 153008 413928 153060
rect 413980 153048 413986 153060
rect 433794 153048 433800 153060
rect 413980 153020 433800 153048
rect 413980 153008 413986 153020
rect 433794 153008 433800 153020
rect 433852 153008 433858 153060
rect 448606 153008 448612 153060
rect 448664 153048 448670 153060
rect 450630 153048 450636 153060
rect 448664 153020 450636 153048
rect 448664 153008 448670 153020
rect 450630 153008 450636 153020
rect 450688 153008 450694 153060
rect 474734 153008 474740 153060
rect 474792 153048 474798 153060
rect 478138 153048 478144 153060
rect 474792 153020 478144 153048
rect 474792 153008 474798 153020
rect 478138 153008 478144 153020
rect 478196 153008 478202 153060
rect 480714 153008 480720 153060
rect 480772 153048 480778 153060
rect 482646 153048 482652 153060
rect 480772 153020 482652 153048
rect 480772 153008 480778 153020
rect 482646 153008 482652 153020
rect 482704 153008 482710 153060
rect 325752 152952 326752 152980
rect 325752 152940 325758 152952
rect 326798 152940 326804 152992
rect 326856 152980 326862 152992
rect 366358 152980 366364 152992
rect 326856 152952 366364 152980
rect 326856 152940 326862 152952
rect 366358 152940 366364 152952
rect 366416 152940 366422 152992
rect 372338 152940 372344 152992
rect 372396 152980 372402 152992
rect 403618 152980 403624 152992
rect 372396 152952 403624 152980
rect 372396 152940 372402 152952
rect 403618 152940 403624 152952
rect 403676 152940 403682 152992
rect 410978 152940 410984 152992
rect 411036 152980 411042 152992
rect 433150 152980 433156 152992
rect 411036 152952 433156 152980
rect 411036 152940 411042 152952
rect 433150 152940 433156 152952
rect 433208 152940 433214 152992
rect 46566 152872 46572 152924
rect 46624 152912 46630 152924
rect 154482 152912 154488 152924
rect 46624 152884 154488 152912
rect 46624 152872 46630 152884
rect 154482 152872 154488 152884
rect 154540 152872 154546 152924
rect 156690 152872 156696 152924
rect 156748 152912 156754 152924
rect 164786 152912 164792 152924
rect 156748 152884 164792 152912
rect 156748 152872 156754 152884
rect 164786 152872 164792 152884
rect 164844 152872 164850 152924
rect 165614 152872 165620 152924
rect 165672 152912 165678 152924
rect 244366 152912 244372 152924
rect 165672 152884 244372 152912
rect 165672 152872 165678 152884
rect 244366 152872 244372 152884
rect 244424 152872 244430 152924
rect 245470 152872 245476 152924
rect 245528 152912 245534 152924
rect 300946 152912 300952 152924
rect 245528 152884 300952 152912
rect 245528 152872 245534 152884
rect 300946 152872 300952 152884
rect 301004 152872 301010 152924
rect 301038 152872 301044 152924
rect 301096 152912 301102 152924
rect 307938 152912 307944 152924
rect 301096 152884 307944 152912
rect 301096 152872 301102 152884
rect 307938 152872 307944 152884
rect 307996 152872 308002 152924
rect 309134 152872 309140 152924
rect 309192 152912 309198 152924
rect 313090 152912 313096 152924
rect 309192 152884 313096 152912
rect 309192 152872 309198 152884
rect 313090 152872 313096 152884
rect 313148 152872 313154 152924
rect 313182 152872 313188 152924
rect 313240 152912 313246 152924
rect 313826 152912 313832 152924
rect 313240 152884 313832 152912
rect 313240 152872 313246 152884
rect 313826 152872 313832 152884
rect 313884 152872 313890 152924
rect 316678 152872 316684 152924
rect 316736 152912 316742 152924
rect 351638 152912 351644 152924
rect 316736 152884 351644 152912
rect 316736 152872 316742 152884
rect 351638 152872 351644 152884
rect 351696 152872 351702 152924
rect 354766 152872 354772 152924
rect 354824 152912 354830 152924
rect 390186 152912 390192 152924
rect 354824 152884 390192 152912
rect 354824 152872 354830 152884
rect 390186 152872 390192 152884
rect 390244 152872 390250 152924
rect 394234 152872 394240 152924
rect 394292 152912 394298 152924
rect 420362 152912 420368 152924
rect 394292 152884 420368 152912
rect 394292 152872 394298 152884
rect 420362 152872 420368 152884
rect 420420 152872 420426 152924
rect 421926 152872 421932 152924
rect 421984 152912 421990 152924
rect 441522 152912 441528 152924
rect 421984 152884 441528 152912
rect 421984 152872 421990 152884
rect 441522 152872 441528 152884
rect 441580 152872 441586 152924
rect 502518 152872 502524 152924
rect 502576 152912 502582 152924
rect 503162 152912 503168 152924
rect 502576 152884 503168 152912
rect 502576 152872 502582 152884
rect 503162 152872 503168 152884
rect 503220 152872 503226 152924
rect 43162 152804 43168 152856
rect 43220 152844 43226 152856
rect 151906 152844 151912 152856
rect 43220 152816 151912 152844
rect 43220 152804 43226 152816
rect 151906 152804 151912 152816
rect 151964 152804 151970 152856
rect 153930 152804 153936 152856
rect 153988 152844 153994 152856
rect 159634 152844 159640 152856
rect 153988 152816 159640 152844
rect 153988 152804 153994 152816
rect 159634 152804 159640 152816
rect 159692 152804 159698 152856
rect 163222 152804 163228 152856
rect 163280 152844 163286 152856
rect 243722 152844 243728 152856
rect 163280 152816 243728 152844
rect 163280 152804 163286 152816
rect 243722 152804 243728 152816
rect 243780 152804 243786 152856
rect 251450 152804 251456 152856
rect 251508 152844 251514 152856
rect 251508 152816 258074 152844
rect 251508 152804 251514 152816
rect 33134 152736 33140 152788
rect 33192 152776 33198 152788
rect 144270 152776 144276 152788
rect 33192 152748 144276 152776
rect 33192 152736 33198 152748
rect 144270 152736 144276 152748
rect 144328 152736 144334 152788
rect 144822 152736 144828 152788
rect 144880 152776 144886 152788
rect 157058 152776 157064 152788
rect 144880 152748 157064 152776
rect 144880 152736 144886 152748
rect 157058 152736 157064 152748
rect 157116 152736 157122 152788
rect 157334 152736 157340 152788
rect 157392 152776 157398 152788
rect 239306 152776 239312 152788
rect 157392 152748 239312 152776
rect 157392 152736 157398 152748
rect 239306 152736 239312 152748
rect 239364 152736 239370 152788
rect 242894 152736 242900 152788
rect 242952 152776 242958 152788
rect 246942 152776 246948 152788
rect 242952 152748 246948 152776
rect 242952 152736 242958 152748
rect 246942 152736 246948 152748
rect 247000 152736 247006 152788
rect 258046 152776 258074 152816
rect 258166 152804 258172 152856
rect 258224 152844 258230 152856
rect 316310 152844 316316 152856
rect 258224 152816 316316 152844
rect 258224 152804 258230 152816
rect 316310 152804 316316 152816
rect 316368 152804 316374 152856
rect 317046 152804 317052 152856
rect 317104 152844 317110 152856
rect 361298 152844 361304 152856
rect 317104 152816 361304 152844
rect 317104 152804 317110 152816
rect 361298 152804 361304 152816
rect 361356 152804 361362 152856
rect 368198 152804 368204 152856
rect 368256 152844 368262 152856
rect 400398 152844 400404 152856
rect 368256 152816 400404 152844
rect 368256 152804 368262 152816
rect 400398 152804 400404 152816
rect 400456 152804 400462 152856
rect 409322 152804 409328 152856
rect 409380 152844 409386 152856
rect 430574 152844 430580 152856
rect 409380 152816 430580 152844
rect 409380 152804 409386 152816
rect 430574 152804 430580 152816
rect 430632 152804 430638 152856
rect 431126 152804 431132 152856
rect 431184 152844 431190 152856
rect 448606 152844 448612 152856
rect 431184 152816 448612 152844
rect 431184 152804 431190 152816
rect 448606 152804 448612 152816
rect 448664 152804 448670 152856
rect 488442 152804 488448 152856
rect 488500 152844 488506 152856
rect 489638 152844 489644 152856
rect 488500 152816 489644 152844
rect 488500 152804 488506 152816
rect 489638 152804 489644 152816
rect 489696 152804 489702 152856
rect 311158 152776 311164 152788
rect 258046 152748 311164 152776
rect 311158 152736 311164 152748
rect 311216 152736 311222 152788
rect 311526 152736 311532 152788
rect 311584 152776 311590 152788
rect 356790 152776 356796 152788
rect 311584 152748 356796 152776
rect 311584 152736 311590 152748
rect 356790 152736 356796 152748
rect 356848 152736 356854 152788
rect 356882 152736 356888 152788
rect 356940 152776 356946 152788
rect 356940 152748 360194 152776
rect 356940 152736 356946 152748
rect 26326 152668 26332 152720
rect 26384 152708 26390 152720
rect 139118 152708 139124 152720
rect 26384 152680 139124 152708
rect 26384 152668 26390 152680
rect 139118 152668 139124 152680
rect 139176 152668 139182 152720
rect 139762 152668 139768 152720
rect 139820 152708 139826 152720
rect 141786 152708 141792 152720
rect 139820 152680 141792 152708
rect 139820 152668 139826 152680
rect 141786 152668 141792 152680
rect 141844 152668 141850 152720
rect 147582 152668 147588 152720
rect 147640 152708 147646 152720
rect 229002 152708 229008 152720
rect 147640 152680 229008 152708
rect 147640 152668 147646 152680
rect 229002 152668 229008 152680
rect 229060 152668 229066 152720
rect 233234 152668 233240 152720
rect 233292 152708 233298 152720
rect 233970 152708 233976 152720
rect 233292 152680 233976 152708
rect 233292 152668 233298 152680
rect 233970 152668 233976 152680
rect 234028 152668 234034 152720
rect 234614 152668 234620 152720
rect 234672 152708 234678 152720
rect 236730 152708 236736 152720
rect 234672 152680 236736 152708
rect 234672 152668 234678 152680
rect 236730 152668 236736 152680
rect 236788 152668 236794 152720
rect 240502 152668 240508 152720
rect 240560 152708 240566 152720
rect 300302 152708 300308 152720
rect 240560 152680 300308 152708
rect 240560 152668 240566 152680
rect 300302 152668 300308 152680
rect 300360 152668 300366 152720
rect 310514 152708 310520 152720
rect 302206 152680 310520 152708
rect 32214 152600 32220 152652
rect 32272 152640 32278 152652
rect 143626 152640 143632 152652
rect 32272 152612 143632 152640
rect 32272 152600 32278 152612
rect 143626 152600 143632 152612
rect 143684 152600 143690 152652
rect 146478 152600 146484 152652
rect 146536 152640 146542 152652
rect 146536 152612 149560 152640
rect 146536 152600 146542 152612
rect 25498 152532 25504 152584
rect 25556 152572 25562 152584
rect 138474 152572 138480 152584
rect 25556 152544 138480 152572
rect 25556 152532 25562 152544
rect 138474 152532 138480 152544
rect 138532 152532 138538 152584
rect 140774 152532 140780 152584
rect 140832 152572 140838 152584
rect 149422 152572 149428 152584
rect 140832 152544 149428 152572
rect 140832 152532 140838 152544
rect 149422 152532 149428 152544
rect 149480 152532 149486 152584
rect 149532 152572 149560 152612
rect 150710 152600 150716 152652
rect 150768 152640 150774 152652
rect 234154 152640 234160 152652
rect 150768 152612 234160 152640
rect 150768 152600 150774 152612
rect 234154 152600 234160 152612
rect 234212 152600 234218 152652
rect 244274 152600 244280 152652
rect 244332 152640 244338 152652
rect 244332 152612 253934 152640
rect 244332 152600 244338 152612
rect 230934 152572 230940 152584
rect 149532 152544 230940 152572
rect 230934 152532 230940 152544
rect 230992 152532 230998 152584
rect 237374 152532 237380 152584
rect 237432 152572 237438 152584
rect 241882 152572 241888 152584
rect 237432 152544 241888 152572
rect 237432 152532 237438 152544
rect 241882 152532 241888 152544
rect 241940 152532 241946 152584
rect 243538 152532 243544 152584
rect 243596 152572 243602 152584
rect 249518 152572 249524 152584
rect 243596 152544 249524 152572
rect 243596 152532 243602 152544
rect 249518 152532 249524 152544
rect 249576 152532 249582 152584
rect 253906 152572 253934 152612
rect 254302 152600 254308 152652
rect 254360 152640 254366 152652
rect 302206 152640 302234 152680
rect 310514 152668 310520 152680
rect 310572 152668 310578 152720
rect 350994 152708 351000 152720
rect 311866 152680 351000 152708
rect 304994 152640 305000 152652
rect 254360 152612 302234 152640
rect 302436 152612 305000 152640
rect 254360 152600 254366 152612
rect 302436 152572 302464 152612
rect 304994 152600 305000 152612
rect 305052 152600 305058 152652
rect 311866 152640 311894 152680
rect 350994 152668 351000 152680
rect 351052 152668 351058 152720
rect 352190 152668 352196 152720
rect 352248 152708 352254 152720
rect 360166 152708 360194 152748
rect 360746 152736 360752 152788
rect 360804 152776 360810 152788
rect 394694 152776 394700 152788
rect 360804 152748 394700 152776
rect 360804 152736 360810 152748
rect 394694 152736 394700 152748
rect 394752 152736 394758 152788
rect 397546 152736 397552 152788
rect 397604 152776 397610 152788
rect 422938 152776 422944 152788
rect 397604 152748 422944 152776
rect 397604 152736 397610 152748
rect 422938 152736 422944 152748
rect 422996 152736 423002 152788
rect 424962 152736 424968 152788
rect 425020 152776 425026 152788
rect 442166 152776 442172 152788
rect 425020 152748 442172 152776
rect 425020 152736 425026 152748
rect 442166 152736 442172 152748
rect 442224 152736 442230 152788
rect 476114 152736 476120 152788
rect 476172 152776 476178 152788
rect 479426 152776 479432 152788
rect 476172 152748 479432 152776
rect 476172 152736 476178 152748
rect 479426 152736 479432 152748
rect 479484 152736 479490 152788
rect 386966 152708 386972 152720
rect 352248 152680 357572 152708
rect 360166 152680 386972 152708
rect 352248 152668 352254 152680
rect 305104 152612 311894 152640
rect 253906 152544 302464 152572
rect 302510 152532 302516 152584
rect 302568 152572 302574 152584
rect 302568 152544 303108 152572
rect 302568 152532 302574 152544
rect 12894 152464 12900 152516
rect 12952 152504 12958 152516
rect 128814 152504 128820 152516
rect 12952 152476 128820 152504
rect 12952 152464 12958 152476
rect 128814 152464 128820 152476
rect 128872 152464 128878 152516
rect 137002 152464 137008 152516
rect 137060 152504 137066 152516
rect 137278 152504 137284 152516
rect 137060 152476 137284 152504
rect 137060 152464 137066 152476
rect 137278 152464 137284 152476
rect 137336 152464 137342 152516
rect 138014 152464 138020 152516
rect 138072 152504 138078 152516
rect 141694 152504 141700 152516
rect 138072 152476 141700 152504
rect 138072 152464 138078 152476
rect 141694 152464 141700 152476
rect 141752 152464 141758 152516
rect 141786 152464 141792 152516
rect 141844 152504 141850 152516
rect 225782 152504 225788 152516
rect 141844 152476 225788 152504
rect 141844 152464 141850 152476
rect 225782 152464 225788 152476
rect 225840 152464 225846 152516
rect 231302 152464 231308 152516
rect 231360 152504 231366 152516
rect 295794 152504 295800 152516
rect 231360 152476 295800 152504
rect 231360 152464 231366 152476
rect 295794 152464 295800 152476
rect 295852 152464 295858 152516
rect 299566 152464 299572 152516
rect 299624 152504 299630 152516
rect 302878 152504 302884 152516
rect 299624 152476 302884 152504
rect 299624 152464 299630 152476
rect 302878 152464 302884 152476
rect 302936 152464 302942 152516
rect 303080 152504 303108 152544
rect 303430 152532 303436 152584
rect 303488 152572 303494 152584
rect 305104 152572 305132 152612
rect 313458 152600 313464 152652
rect 313516 152640 313522 152652
rect 318886 152640 318892 152652
rect 313516 152612 318892 152640
rect 313516 152600 313522 152612
rect 318886 152600 318892 152612
rect 318944 152600 318950 152652
rect 318978 152600 318984 152652
rect 319036 152640 319042 152652
rect 357434 152640 357440 152652
rect 319036 152612 357440 152640
rect 319036 152600 319042 152612
rect 357434 152600 357440 152612
rect 357492 152600 357498 152652
rect 303488 152544 305132 152572
rect 303488 152532 303494 152544
rect 305178 152532 305184 152584
rect 305236 152572 305242 152584
rect 352282 152572 352288 152584
rect 305236 152544 352288 152572
rect 305236 152532 305242 152544
rect 352282 152532 352288 152544
rect 352340 152532 352346 152584
rect 356882 152572 356888 152584
rect 352392 152544 356888 152572
rect 346486 152504 346492 152516
rect 303080 152476 346492 152504
rect 346486 152464 346492 152476
rect 346544 152464 346550 152516
rect 350534 152464 350540 152516
rect 350592 152504 350598 152516
rect 352392 152504 352420 152544
rect 356882 152532 356888 152544
rect 356940 152532 356946 152584
rect 357544 152572 357572 152680
rect 386966 152668 386972 152680
rect 387024 152668 387030 152720
rect 389174 152668 389180 152720
rect 389232 152708 389238 152720
rect 416498 152708 416504 152720
rect 389232 152680 416504 152708
rect 389232 152668 389238 152680
rect 416498 152668 416504 152680
rect 416556 152668 416562 152720
rect 417694 152668 417700 152720
rect 417752 152708 417758 152720
rect 438302 152708 438308 152720
rect 417752 152680 438308 152708
rect 417752 152668 417758 152680
rect 438302 152668 438308 152680
rect 438360 152668 438366 152720
rect 485866 152668 485872 152720
rect 485924 152708 485930 152720
rect 488442 152708 488448 152720
rect 485924 152680 488448 152708
rect 485924 152668 485930 152680
rect 488442 152668 488448 152680
rect 488500 152668 488506 152720
rect 357986 152600 357992 152652
rect 358044 152640 358050 152652
rect 360010 152640 360016 152652
rect 358044 152612 360016 152640
rect 358044 152600 358050 152612
rect 360010 152600 360016 152612
rect 360068 152600 360074 152652
rect 361482 152600 361488 152652
rect 361540 152640 361546 152652
rect 395338 152640 395344 152652
rect 361540 152612 395344 152640
rect 361540 152600 361546 152612
rect 395338 152600 395344 152612
rect 395396 152600 395402 152652
rect 395430 152600 395436 152652
rect 395488 152640 395494 152652
rect 397822 152640 397828 152652
rect 395488 152612 397828 152640
rect 395488 152600 395494 152612
rect 397822 152600 397828 152612
rect 397880 152600 397886 152652
rect 402606 152600 402612 152652
rect 402664 152640 402670 152652
rect 426802 152640 426808 152652
rect 402664 152612 426808 152640
rect 402664 152600 402670 152612
rect 426802 152600 426808 152612
rect 426860 152600 426866 152652
rect 430298 152600 430304 152652
rect 430356 152640 430362 152652
rect 447962 152640 447968 152652
rect 430356 152612 447968 152640
rect 430356 152600 430362 152612
rect 447962 152600 447968 152612
rect 448020 152600 448026 152652
rect 388254 152572 388260 152584
rect 357544 152544 388260 152572
rect 388254 152532 388260 152544
rect 388312 152532 388318 152584
rect 395890 152532 395896 152584
rect 395948 152572 395954 152584
rect 421650 152572 421656 152584
rect 395948 152544 421656 152572
rect 395948 152532 395954 152544
rect 421650 152532 421656 152544
rect 421708 152532 421714 152584
rect 426158 152532 426164 152584
rect 426216 152572 426222 152584
rect 444742 152572 444748 152584
rect 426216 152544 444748 152572
rect 426216 152532 426222 152544
rect 444742 152532 444748 152544
rect 444800 152532 444806 152584
rect 350592 152476 352420 152504
rect 350592 152464 350598 152476
rect 355226 152464 355232 152516
rect 355284 152504 355290 152516
rect 384390 152504 384396 152516
rect 355284 152476 384396 152504
rect 355284 152464 355290 152476
rect 384390 152464 384396 152476
rect 384448 152464 384454 152516
rect 384942 152464 384948 152516
rect 385000 152504 385006 152516
rect 413094 152504 413100 152516
rect 385000 152476 413100 152504
rect 385000 152464 385006 152476
rect 413094 152464 413100 152476
rect 413152 152464 413158 152516
rect 415210 152464 415216 152516
rect 415268 152504 415274 152516
rect 436370 152504 436376 152516
rect 415268 152476 436376 152504
rect 415268 152464 415274 152476
rect 436370 152464 436376 152476
rect 436428 152464 436434 152516
rect 477586 152464 477592 152516
rect 477644 152504 477650 152516
rect 480070 152504 480076 152516
rect 477644 152476 480076 152504
rect 477644 152464 477650 152476
rect 480070 152464 480076 152476
rect 480128 152464 480134 152516
rect 86862 152396 86868 152448
rect 86920 152436 86926 152448
rect 185302 152436 185308 152448
rect 86920 152408 185308 152436
rect 86920 152396 86926 152408
rect 185302 152396 185308 152408
rect 185360 152396 185366 152448
rect 188982 152396 188988 152448
rect 189040 152436 189046 152448
rect 193030 152436 193036 152448
rect 189040 152408 193036 152436
rect 189040 152396 189046 152408
rect 193030 152396 193036 152408
rect 193088 152396 193094 152448
rect 195974 152396 195980 152448
rect 196032 152436 196038 152448
rect 198182 152436 198188 152448
rect 196032 152408 198188 152436
rect 196032 152396 196038 152408
rect 198182 152396 198188 152408
rect 198240 152396 198246 152448
rect 203610 152396 203616 152448
rect 203668 152436 203674 152448
rect 274542 152436 274548 152448
rect 203668 152408 274548 152436
rect 203668 152396 203674 152408
rect 274542 152396 274548 152408
rect 274600 152396 274606 152448
rect 274634 152396 274640 152448
rect 274692 152436 274698 152448
rect 282270 152436 282276 152448
rect 274692 152408 282276 152436
rect 274692 152396 274698 152408
rect 282270 152396 282276 152408
rect 282328 152396 282334 152448
rect 282914 152396 282920 152448
rect 282972 152436 282978 152448
rect 288066 152436 288072 152448
rect 282972 152408 288072 152436
rect 282972 152396 282978 152408
rect 288066 152396 288072 152408
rect 288124 152396 288130 152448
rect 288158 152396 288164 152448
rect 288216 152436 288222 152448
rect 336182 152436 336188 152448
rect 288216 152408 336188 152436
rect 288216 152396 288222 152408
rect 336182 152396 336188 152408
rect 336240 152396 336246 152448
rect 338758 152396 338764 152448
rect 338816 152436 338822 152448
rect 377950 152436 377956 152448
rect 338816 152408 377956 152436
rect 338816 152396 338822 152408
rect 377950 152396 377956 152408
rect 378008 152396 378014 152448
rect 378226 152396 378232 152448
rect 378284 152436 378290 152448
rect 408126 152436 408132 152448
rect 378284 152408 408132 152436
rect 378284 152396 378290 152408
rect 408126 152396 408132 152408
rect 408184 152396 408190 152448
rect 408862 152396 408868 152448
rect 408920 152436 408926 152448
rect 428642 152436 428648 152448
rect 408920 152408 428648 152436
rect 408920 152396 408926 152408
rect 428642 152396 428648 152408
rect 428700 152396 428706 152448
rect 428734 152396 428740 152448
rect 428792 152436 428798 152448
rect 446674 152436 446680 152448
rect 428792 152408 446680 152436
rect 428792 152396 428798 152408
rect 446674 152396 446680 152408
rect 446732 152396 446738 152448
rect 50338 152328 50344 152380
rect 50396 152368 50402 152380
rect 146754 152368 146760 152380
rect 50396 152340 146760 152368
rect 50396 152328 50402 152340
rect 146754 152328 146760 152340
rect 146812 152328 146818 152380
rect 161198 152328 161204 152380
rect 161256 152368 161262 152380
rect 169938 152368 169944 152380
rect 161256 152340 169944 152368
rect 161256 152328 161262 152340
rect 169938 152328 169944 152340
rect 169996 152328 170002 152380
rect 173250 152328 173256 152380
rect 173308 152368 173314 152380
rect 243538 152368 243544 152380
rect 173308 152340 243544 152368
rect 173308 152328 173314 152340
rect 243538 152328 243544 152340
rect 243596 152328 243602 152380
rect 248138 152328 248144 152380
rect 248196 152368 248202 152380
rect 252094 152368 252100 152380
rect 248196 152340 252100 152368
rect 248196 152328 248202 152340
rect 252094 152328 252100 152340
rect 252152 152328 252158 152380
rect 252554 152328 252560 152380
rect 252612 152368 252618 152380
rect 306006 152368 306012 152380
rect 252612 152340 306012 152368
rect 252612 152328 252618 152340
rect 306006 152328 306012 152340
rect 306064 152328 306070 152380
rect 310606 152328 310612 152380
rect 310664 152368 310670 152380
rect 313734 152368 313740 152380
rect 310664 152340 313740 152368
rect 310664 152328 310670 152340
rect 313734 152328 313740 152340
rect 313792 152328 313798 152380
rect 313826 152328 313832 152380
rect 313884 152368 313890 152380
rect 318978 152368 318984 152380
rect 313884 152340 318984 152368
rect 313884 152328 313890 152340
rect 318978 152328 318984 152340
rect 319036 152328 319042 152380
rect 319346 152328 319352 152380
rect 319404 152368 319410 152380
rect 361942 152368 361948 152380
rect 319404 152340 361948 152368
rect 319404 152328 319410 152340
rect 361942 152328 361948 152340
rect 362000 152328 362006 152380
rect 362678 152328 362684 152380
rect 362736 152368 362742 152380
rect 365162 152368 365168 152380
rect 362736 152340 365168 152368
rect 362736 152328 362742 152340
rect 365162 152328 365168 152340
rect 365220 152328 365226 152380
rect 377214 152328 377220 152380
rect 377272 152368 377278 152380
rect 381814 152368 381820 152380
rect 377272 152340 381820 152368
rect 377272 152328 377278 152340
rect 381814 152328 381820 152340
rect 381872 152328 381878 152380
rect 384114 152328 384120 152380
rect 384172 152368 384178 152380
rect 412634 152368 412640 152380
rect 384172 152340 412640 152368
rect 384172 152328 384178 152340
rect 412634 152328 412640 152340
rect 412692 152328 412698 152380
rect 415486 152328 415492 152380
rect 415544 152368 415550 152380
rect 419074 152368 419080 152380
rect 415544 152340 419080 152368
rect 415544 152328 415550 152340
rect 419074 152328 419080 152340
rect 419132 152328 419138 152380
rect 419166 152328 419172 152380
rect 419224 152368 419230 152380
rect 429286 152368 429292 152380
rect 419224 152340 429292 152368
rect 419224 152328 419230 152340
rect 429286 152328 429292 152340
rect 429344 152328 429350 152380
rect 429470 152328 429476 152380
rect 429528 152368 429534 152380
rect 447318 152368 447324 152380
rect 429528 152340 447324 152368
rect 429528 152328 429534 152340
rect 447318 152328 447324 152340
rect 447376 152328 447382 152380
rect 100294 152260 100300 152312
rect 100352 152300 100358 152312
rect 195606 152300 195612 152312
rect 100352 152272 195612 152300
rect 100352 152260 100358 152272
rect 195606 152260 195612 152272
rect 195664 152260 195670 152312
rect 204438 152260 204444 152312
rect 204496 152300 204502 152312
rect 275186 152300 275192 152312
rect 204496 152272 275192 152300
rect 204496 152260 204502 152272
rect 275186 152260 275192 152272
rect 275244 152260 275250 152312
rect 279510 152260 279516 152312
rect 279568 152300 279574 152312
rect 282914 152300 282920 152312
rect 279568 152272 282920 152300
rect 279568 152260 279574 152272
rect 282914 152260 282920 152272
rect 282972 152260 282978 152312
rect 292758 152300 292764 152312
rect 283208 152272 292764 152300
rect 107010 152192 107016 152244
rect 107068 152232 107074 152244
rect 200758 152232 200764 152244
rect 107068 152204 200764 152232
rect 107068 152192 107074 152204
rect 200758 152192 200764 152204
rect 200816 152192 200822 152244
rect 213086 152192 213092 152244
rect 213144 152232 213150 152244
rect 216122 152232 216128 152244
rect 213144 152204 216128 152232
rect 213144 152192 213150 152204
rect 216122 152192 216128 152204
rect 216180 152192 216186 152244
rect 280338 152232 280344 152244
rect 216232 152204 280344 152232
rect 110322 152124 110328 152176
rect 110380 152164 110386 152176
rect 203334 152164 203340 152176
rect 110380 152136 203340 152164
rect 110380 152124 110386 152136
rect 203334 152124 203340 152136
rect 203392 152124 203398 152176
rect 210326 152124 210332 152176
rect 210384 152164 210390 152176
rect 210384 152136 211108 152164
rect 210384 152124 210390 152136
rect 6086 152056 6092 152108
rect 6144 152096 6150 152108
rect 80606 152096 80612 152108
rect 6144 152068 80612 152096
rect 6144 152056 6150 152068
rect 80606 152056 80612 152068
rect 80664 152056 80670 152108
rect 81710 152056 81716 152108
rect 81768 152096 81774 152108
rect 92474 152096 92480 152108
rect 81768 152068 92480 152096
rect 81768 152056 81774 152068
rect 92474 152056 92480 152068
rect 92532 152056 92538 152108
rect 105814 152056 105820 152108
rect 105872 152096 105878 152108
rect 116486 152096 116492 152108
rect 105872 152068 116492 152096
rect 105872 152056 105878 152068
rect 116486 152056 116492 152068
rect 116544 152056 116550 152108
rect 119614 152056 119620 152108
rect 119672 152096 119678 152108
rect 210418 152096 210424 152108
rect 119672 152068 210424 152096
rect 119672 152056 119678 152068
rect 210418 152056 210424 152068
rect 210476 152056 210482 152108
rect 211080 152096 211108 152136
rect 211154 152124 211160 152176
rect 211212 152164 211218 152176
rect 216232 152164 216260 152204
rect 280338 152192 280344 152204
rect 280396 152192 280402 152244
rect 281442 152192 281448 152244
rect 281500 152232 281506 152244
rect 283208 152232 283236 152272
rect 292758 152260 292764 152272
rect 292816 152260 292822 152312
rect 341334 152300 341340 152312
rect 292868 152272 341340 152300
rect 281500 152204 283236 152232
rect 281500 152192 281506 152204
rect 284386 152192 284392 152244
rect 284444 152232 284450 152244
rect 288158 152232 288164 152244
rect 284444 152204 288164 152232
rect 284444 152192 284450 152204
rect 288158 152192 288164 152204
rect 288216 152192 288222 152244
rect 290918 152192 290924 152244
rect 290976 152232 290982 152244
rect 292868 152232 292896 152272
rect 341334 152260 341340 152272
rect 341392 152260 341398 152312
rect 342162 152260 342168 152312
rect 342220 152300 342226 152312
rect 344554 152300 344560 152312
rect 342220 152272 344560 152300
rect 342220 152260 342226 152272
rect 344554 152260 344560 152272
rect 344612 152260 344618 152312
rect 344646 152260 344652 152312
rect 344704 152300 344710 152312
rect 379882 152300 379888 152312
rect 344704 152272 379888 152300
rect 344704 152260 344710 152272
rect 379882 152260 379888 152272
rect 379940 152260 379946 152312
rect 380986 152260 380992 152312
rect 381044 152300 381050 152312
rect 392118 152300 392124 152312
rect 381044 152272 392124 152300
rect 381044 152260 381050 152272
rect 392118 152260 392124 152272
rect 392176 152260 392182 152312
rect 392302 152260 392308 152312
rect 392360 152300 392366 152312
rect 417786 152300 417792 152312
rect 392360 152272 417792 152300
rect 392360 152260 392366 152272
rect 417786 152260 417792 152272
rect 417844 152260 417850 152312
rect 431218 152300 431224 152312
rect 422266 152272 431224 152300
rect 290976 152204 292896 152232
rect 290976 152192 290982 152204
rect 293126 152192 293132 152244
rect 293184 152232 293190 152244
rect 295058 152232 295064 152244
rect 293184 152204 295064 152232
rect 293184 152192 293190 152204
rect 295058 152192 295064 152204
rect 295116 152192 295122 152244
rect 295168 152204 295472 152232
rect 279694 152164 279700 152176
rect 211212 152136 216260 152164
rect 216324 152136 279700 152164
rect 211212 152124 211218 152136
rect 216324 152096 216352 152136
rect 279694 152124 279700 152136
rect 279752 152124 279758 152176
rect 282454 152124 282460 152176
rect 282512 152164 282518 152176
rect 295168 152164 295196 152204
rect 282512 152136 295196 152164
rect 295444 152164 295472 152204
rect 295518 152192 295524 152244
rect 295576 152232 295582 152244
rect 340690 152232 340696 152244
rect 295576 152204 340696 152232
rect 295576 152192 295582 152204
rect 340690 152192 340696 152204
rect 340748 152192 340754 152244
rect 340782 152192 340788 152244
rect 340840 152232 340846 152244
rect 377306 152232 377312 152244
rect 340840 152204 377312 152232
rect 340840 152192 340846 152204
rect 377306 152192 377312 152204
rect 377364 152192 377370 152244
rect 380894 152192 380900 152244
rect 380952 152232 380958 152244
rect 389542 152232 389548 152244
rect 380952 152204 389548 152232
rect 380952 152192 380958 152204
rect 389542 152192 389548 152204
rect 389600 152192 389606 152244
rect 390922 152192 390928 152244
rect 390980 152232 390986 152244
rect 415210 152232 415216 152244
rect 390980 152204 415216 152232
rect 390980 152192 390986 152204
rect 415210 152192 415216 152204
rect 415268 152192 415274 152244
rect 331122 152164 331128 152176
rect 295444 152136 331128 152164
rect 282512 152124 282518 152136
rect 331122 152124 331128 152136
rect 331180 152124 331186 152176
rect 333974 152124 333980 152176
rect 334032 152164 334038 152176
rect 372798 152164 372804 152176
rect 334032 152136 372804 152164
rect 334032 152124 334038 152136
rect 372798 152124 372804 152136
rect 372856 152124 372862 152176
rect 388530 152124 388536 152176
rect 388588 152164 388594 152176
rect 410058 152164 410064 152176
rect 388588 152136 410064 152164
rect 388588 152124 388594 152136
rect 410058 152124 410064 152136
rect 410116 152124 410122 152176
rect 411714 152124 411720 152176
rect 411772 152164 411778 152176
rect 422266 152164 422294 152272
rect 431218 152260 431224 152272
rect 431276 152260 431282 152312
rect 444098 152300 444104 152312
rect 431788 152272 444104 152300
rect 423214 152192 423220 152244
rect 423272 152232 423278 152244
rect 423272 152204 423720 152232
rect 423272 152192 423278 152204
rect 411772 152136 422294 152164
rect 411772 152124 411778 152136
rect 211080 152068 216352 152096
rect 217042 152056 217048 152108
rect 217100 152096 217106 152108
rect 284846 152096 284852 152108
rect 217100 152068 284852 152096
rect 217100 152056 217106 152068
rect 284846 152056 284852 152068
rect 284904 152056 284910 152108
rect 287330 152056 287336 152108
rect 287388 152096 287394 152108
rect 289998 152096 290004 152108
rect 287388 152068 290004 152096
rect 287388 152056 287394 152068
rect 289998 152056 290004 152068
rect 290056 152056 290062 152108
rect 290090 152056 290096 152108
rect 290148 152096 290154 152108
rect 295334 152096 295340 152108
rect 290148 152068 295340 152096
rect 290148 152056 290154 152068
rect 295334 152056 295340 152068
rect 295392 152056 295398 152108
rect 341978 152096 341984 152108
rect 295444 152068 341984 152096
rect 47302 151988 47308 152040
rect 47360 152028 47366 152040
rect 110046 152028 110052 152040
rect 47360 152000 110052 152028
rect 47360 151988 47366 152000
rect 110046 151988 110052 152000
rect 110104 151988 110110 152040
rect 123386 151988 123392 152040
rect 123444 152028 123450 152040
rect 128170 152028 128176 152040
rect 123444 152000 128176 152028
rect 123444 151988 123450 152000
rect 128170 151988 128176 152000
rect 128228 151988 128234 152040
rect 128446 151988 128452 152040
rect 128504 152028 128510 152040
rect 213546 152028 213552 152040
rect 128504 152000 213552 152028
rect 128504 151988 128510 152000
rect 213546 151988 213552 152000
rect 213604 151988 213610 152040
rect 214374 151988 214380 152040
rect 214432 152028 214438 152040
rect 221274 152028 221280 152040
rect 214432 152000 221280 152028
rect 214432 151988 214438 152000
rect 221274 151988 221280 152000
rect 221332 151988 221338 152040
rect 223574 151988 223580 152040
rect 223632 152028 223638 152040
rect 226426 152028 226432 152040
rect 223632 152000 226432 152028
rect 223632 151988 223638 152000
rect 226426 151988 226432 152000
rect 226484 151988 226490 152040
rect 290642 152028 290648 152040
rect 226812 152000 290648 152028
rect 54202 151920 54208 151972
rect 54260 151960 54266 151972
rect 116670 151960 116676 151972
rect 54260 151932 116676 151960
rect 54260 151920 54266 151932
rect 116670 151920 116676 151932
rect 116728 151920 116734 151972
rect 125686 151920 125692 151972
rect 125744 151960 125750 151972
rect 139762 151960 139768 151972
rect 125744 151932 128354 151960
rect 125744 151920 125750 151932
rect 40494 151852 40500 151904
rect 40552 151892 40558 151904
rect 109954 151892 109960 151904
rect 40552 151864 109960 151892
rect 40552 151852 40558 151864
rect 109954 151852 109960 151864
rect 110012 151852 110018 151904
rect 110138 151852 110144 151904
rect 110196 151892 110202 151904
rect 126882 151892 126888 151904
rect 110196 151864 126888 151892
rect 110196 151852 110202 151864
rect 126882 151852 126888 151864
rect 126940 151852 126946 151904
rect 128326 151892 128354 151932
rect 128464 151932 139768 151960
rect 128464 151892 128492 151932
rect 139762 151920 139768 151932
rect 139820 151920 139826 151972
rect 142614 151920 142620 151972
rect 142672 151960 142678 151972
rect 223850 151960 223856 151972
rect 142672 151932 223856 151960
rect 142672 151920 142678 151932
rect 223850 151920 223856 151932
rect 223908 151920 223914 151972
rect 224586 151920 224592 151972
rect 224644 151960 224650 151972
rect 226812 151960 226840 152000
rect 290642 151988 290648 152000
rect 290700 151988 290706 152040
rect 292758 151988 292764 152040
rect 292816 152028 292822 152040
rect 295150 152028 295156 152040
rect 292816 152000 295156 152028
rect 292816 151988 292822 152000
rect 295150 151988 295156 152000
rect 295208 151988 295214 152040
rect 295242 151988 295248 152040
rect 295300 152028 295306 152040
rect 295444 152028 295472 152068
rect 341978 152056 341984 152068
rect 342036 152056 342042 152108
rect 342070 152056 342076 152108
rect 342128 152096 342134 152108
rect 344646 152096 344652 152108
rect 342128 152068 344652 152096
rect 342128 152056 342134 152068
rect 344646 152056 344652 152068
rect 344704 152056 344710 152108
rect 345474 152056 345480 152108
rect 345532 152096 345538 152108
rect 345532 152068 345980 152096
rect 345532 152056 345538 152068
rect 295300 152000 295472 152028
rect 295300 151988 295306 152000
rect 296806 151988 296812 152040
rect 296864 152028 296870 152040
rect 345842 152028 345848 152040
rect 296864 152000 345848 152028
rect 296864 151988 296870 152000
rect 345842 151988 345848 152000
rect 345900 151988 345906 152040
rect 345952 152028 345980 152068
rect 347130 152056 347136 152108
rect 347188 152096 347194 152108
rect 355226 152096 355232 152108
rect 347188 152068 355232 152096
rect 347188 152056 347194 152068
rect 355226 152056 355232 152068
rect 355284 152056 355290 152108
rect 355318 152056 355324 152108
rect 355376 152096 355382 152108
rect 383102 152096 383108 152108
rect 355376 152068 383108 152096
rect 355376 152056 355382 152068
rect 383102 152056 383108 152068
rect 383160 152056 383166 152108
rect 388438 152056 388444 152108
rect 388496 152096 388502 152108
rect 404906 152096 404912 152108
rect 388496 152068 404912 152096
rect 388496 152056 388502 152068
rect 404906 152056 404912 152068
rect 404964 152056 404970 152108
rect 404998 152056 405004 152108
rect 405056 152096 405062 152108
rect 423582 152096 423588 152108
rect 405056 152068 423588 152096
rect 405056 152056 405062 152068
rect 423582 152056 423588 152068
rect 423640 152056 423646 152108
rect 423692 152096 423720 152204
rect 425238 152192 425244 152244
rect 425296 152232 425302 152244
rect 431788 152232 431816 152272
rect 444098 152260 444104 152272
rect 444156 152260 444162 152312
rect 425296 152204 431816 152232
rect 425296 152192 425302 152204
rect 508406 152192 508412 152244
rect 508464 152232 508470 152244
rect 509142 152232 509148 152244
rect 508464 152204 509148 152232
rect 508464 152192 508470 152204
rect 509142 152192 509148 152204
rect 509200 152192 509206 152244
rect 439590 152164 439596 152176
rect 431328 152136 439596 152164
rect 431328 152096 431356 152136
rect 439590 152124 439596 152136
rect 439648 152124 439654 152176
rect 423692 152068 431356 152096
rect 347222 152028 347228 152040
rect 345952 152000 347228 152028
rect 347222 151988 347228 152000
rect 347280 151988 347286 152040
rect 348050 151988 348056 152040
rect 348108 152028 348114 152040
rect 385034 152028 385040 152040
rect 348108 152000 385040 152028
rect 348108 151988 348114 152000
rect 385034 151988 385040 152000
rect 385092 151988 385098 152040
rect 385678 151988 385684 152040
rect 385736 152028 385742 152040
rect 399754 152028 399760 152040
rect 385736 152000 399760 152028
rect 385736 151988 385742 152000
rect 399754 151988 399760 152000
rect 399812 151988 399818 152040
rect 407298 151988 407304 152040
rect 407356 152028 407362 152040
rect 426158 152028 426164 152040
rect 407356 152000 426164 152028
rect 407356 151988 407362 152000
rect 426158 151988 426164 152000
rect 426216 151988 426222 152040
rect 430574 151988 430580 152040
rect 430632 152028 430638 152040
rect 431770 152028 431776 152040
rect 430632 152000 431776 152028
rect 430632 151988 430638 152000
rect 431770 151988 431776 152000
rect 431828 151988 431834 152040
rect 488534 151988 488540 152040
rect 488592 152028 488598 152040
rect 490926 152028 490932 152040
rect 488592 152000 490932 152028
rect 488592 151988 488598 152000
rect 490926 151988 490932 152000
rect 490984 151988 490990 152040
rect 224644 151932 226840 151960
rect 224644 151920 224650 151932
rect 226978 151920 226984 151972
rect 227036 151960 227042 151972
rect 227036 151932 233924 151960
rect 227036 151920 227042 151932
rect 128326 151864 128492 151892
rect 128538 151852 128544 151904
rect 128596 151892 128602 151904
rect 208486 151892 208492 151904
rect 128596 151864 208492 151892
rect 128596 151852 128602 151864
rect 208486 151852 208492 151864
rect 208544 151852 208550 151904
rect 208670 151852 208676 151904
rect 208728 151892 208734 151904
rect 211062 151892 211068 151904
rect 208728 151864 211068 151892
rect 208728 151852 208734 151864
rect 211062 151852 211068 151864
rect 211120 151852 211126 151904
rect 227806 151852 227812 151904
rect 227864 151892 227870 151904
rect 231578 151892 231584 151904
rect 227864 151864 231584 151892
rect 227864 151852 227870 151864
rect 231578 151852 231584 151864
rect 231636 151852 231642 151904
rect 233896 151892 233924 151932
rect 233970 151920 233976 151972
rect 234028 151960 234034 151972
rect 262674 151960 262680 151972
rect 234028 151932 262680 151960
rect 234028 151920 234034 151932
rect 262674 151920 262680 151932
rect 262732 151920 262738 151972
rect 262766 151920 262772 151972
rect 262824 151960 262830 151972
rect 267550 151960 267556 151972
rect 262824 151932 267556 151960
rect 262824 151920 262830 151932
rect 267550 151920 267556 151932
rect 267608 151920 267614 151972
rect 269022 151920 269028 151972
rect 269080 151960 269086 151972
rect 277118 151960 277124 151972
rect 269080 151932 277124 151960
rect 269080 151920 269086 151932
rect 277118 151920 277124 151932
rect 277176 151920 277182 151972
rect 277210 151920 277216 151972
rect 277268 151960 277274 151972
rect 316586 151960 316592 151972
rect 277268 151932 316592 151960
rect 277268 151920 277274 151932
rect 316586 151920 316592 151932
rect 316644 151920 316650 151972
rect 316696 151932 321554 151960
rect 289998 151892 290004 151904
rect 233896 151864 258074 151892
rect 77110 151784 77116 151836
rect 77168 151824 77174 151836
rect 128078 151824 128084 151836
rect 77168 151796 128084 151824
rect 77168 151784 77174 151796
rect 128078 151784 128084 151796
rect 128136 151784 128142 151836
rect 128262 151784 128268 151836
rect 128320 151824 128326 151836
rect 167546 151824 167552 151836
rect 128320 151796 167552 151824
rect 128320 151784 128326 151796
rect 167546 151784 167552 151796
rect 167604 151784 167610 151836
rect 167638 151784 167644 151836
rect 167696 151824 167702 151836
rect 172514 151824 172520 151836
rect 167696 151796 172520 151824
rect 167696 151784 167702 151796
rect 172514 151784 172520 151796
rect 172572 151784 172578 151836
rect 190840 151796 191880 151824
rect 96522 151716 96528 151768
rect 96580 151756 96586 151768
rect 190730 151756 190736 151768
rect 96580 151728 190736 151756
rect 96580 151716 96586 151728
rect 190730 151716 190736 151728
rect 190788 151716 190794 151768
rect 97718 151648 97724 151700
rect 97776 151688 97782 151700
rect 190840 151688 190868 151796
rect 190914 151716 190920 151768
rect 190972 151756 190978 151768
rect 191742 151756 191748 151768
rect 190972 151728 191748 151756
rect 190972 151716 190978 151728
rect 191742 151716 191748 151728
rect 191800 151716 191806 151768
rect 191852 151756 191880 151796
rect 194594 151784 194600 151836
rect 194652 151824 194658 151836
rect 254670 151824 254676 151836
rect 194652 151796 254676 151824
rect 194652 151784 194658 151796
rect 254670 151784 254676 151796
rect 254728 151784 254734 151836
rect 258046 151824 258074 151864
rect 262784 151864 290004 151892
rect 262784 151824 262812 151864
rect 289998 151852 290004 151864
rect 290056 151852 290062 151904
rect 290090 151852 290096 151904
rect 290148 151892 290154 151904
rect 297726 151892 297732 151904
rect 290148 151864 297732 151892
rect 290148 151852 290154 151864
rect 297726 151852 297732 151864
rect 297784 151852 297790 151904
rect 297818 151852 297824 151904
rect 297876 151892 297882 151904
rect 302510 151892 302516 151904
rect 297876 151864 302516 151892
rect 297876 151852 297882 151864
rect 302510 151852 302516 151864
rect 302568 151852 302574 151904
rect 316696 151892 316724 151932
rect 302620 151864 316724 151892
rect 321526 151892 321554 151932
rect 323670 151920 323676 151972
rect 323728 151960 323734 151972
rect 326798 151960 326804 151972
rect 323728 151932 326804 151960
rect 323728 151920 323734 151932
rect 326798 151920 326804 151932
rect 326856 151920 326862 151972
rect 328426 151932 332732 151960
rect 328426 151892 328454 151932
rect 321526 151864 328454 151892
rect 332704 151892 332732 151932
rect 332778 151920 332784 151972
rect 332836 151960 332842 151972
rect 367002 151960 367008 151972
rect 332836 151932 367008 151960
rect 332836 151920 332842 151932
rect 367002 151920 367008 151932
rect 367060 151920 367066 151972
rect 386230 151920 386236 151972
rect 386288 151960 386294 151972
rect 397178 151960 397184 151972
rect 386288 151932 397184 151960
rect 386288 151920 386294 151932
rect 397178 151920 397184 151932
rect 397236 151920 397242 151972
rect 398098 151920 398104 151972
rect 398156 151960 398162 151972
rect 405550 151960 405556 151972
rect 398156 151932 405556 151960
rect 398156 151920 398162 151932
rect 405550 151920 405556 151932
rect 405608 151920 405614 151972
rect 405642 151920 405648 151972
rect 405700 151960 405706 151972
rect 421006 151960 421012 151972
rect 405700 151932 421012 151960
rect 405700 151920 405706 151932
rect 421006 151920 421012 151932
rect 421064 151920 421070 151972
rect 422570 151920 422576 151972
rect 422628 151960 422634 151972
rect 437014 151960 437020 151972
rect 422628 151932 437020 151960
rect 422628 151920 422634 151932
rect 437014 151920 437020 151932
rect 437072 151920 437078 151972
rect 479518 151920 479524 151972
rect 479576 151960 479582 151972
rect 481358 151960 481364 151972
rect 479576 151932 481364 151960
rect 479576 151920 479582 151932
rect 481358 151920 481364 151932
rect 481416 151920 481422 151972
rect 507026 151920 507032 151972
rect 507084 151960 507090 151972
rect 507578 151960 507584 151972
rect 507084 151932 507584 151960
rect 507084 151920 507090 151932
rect 507578 151920 507584 151932
rect 507636 151920 507642 151972
rect 332704 151864 340874 151892
rect 258046 151796 262812 151824
rect 262858 151784 262864 151836
rect 262916 151824 262922 151836
rect 270126 151824 270132 151836
rect 262916 151796 270132 151824
rect 262916 151784 262922 151796
rect 270126 151784 270132 151796
rect 270184 151784 270190 151836
rect 271506 151784 271512 151836
rect 271564 151824 271570 151836
rect 274634 151824 274640 151836
rect 271564 151796 274640 151824
rect 271564 151784 271570 151796
rect 274634 151784 274640 151796
rect 274692 151784 274698 151836
rect 274726 151784 274732 151836
rect 274784 151824 274790 151836
rect 292574 151824 292580 151836
rect 274784 151796 292580 151824
rect 274784 151784 274790 151796
rect 292574 151784 292580 151796
rect 292632 151784 292638 151836
rect 293954 151784 293960 151836
rect 294012 151824 294018 151836
rect 298370 151824 298376 151836
rect 294012 151796 298376 151824
rect 294012 151784 294018 151796
rect 298370 151784 298376 151796
rect 298428 151784 298434 151836
rect 298462 151784 298468 151836
rect 298520 151824 298526 151836
rect 302620 151824 302648 151864
rect 298520 151796 302648 151824
rect 298520 151784 298526 151796
rect 306374 151784 306380 151836
rect 306432 151824 306438 151836
rect 316678 151824 316684 151836
rect 306432 151796 316684 151824
rect 306432 151784 306438 151796
rect 316678 151784 316684 151796
rect 316736 151784 316742 151836
rect 325970 151824 325976 151836
rect 316788 151796 325976 151824
rect 193674 151756 193680 151768
rect 191852 151728 193680 151756
rect 193674 151716 193680 151728
rect 193732 151716 193738 151768
rect 265618 151756 265624 151768
rect 195946 151728 265624 151756
rect 97776 151660 190868 151688
rect 97776 151648 97782 151660
rect 191006 151648 191012 151700
rect 191064 151688 191070 151700
rect 195054 151688 195060 151700
rect 191064 151660 195060 151688
rect 191064 151648 191070 151660
rect 195054 151648 195060 151660
rect 195112 151648 195118 151700
rect 85390 151580 85396 151632
rect 85448 151620 85454 151632
rect 183370 151620 183376 151632
rect 85448 151592 183376 151620
rect 85448 151580 85454 151592
rect 183370 151580 183376 151592
rect 183428 151580 183434 151632
rect 186222 151580 186228 151632
rect 186280 151620 186286 151632
rect 191098 151620 191104 151632
rect 186280 151592 191104 151620
rect 186280 151580 186286 151592
rect 191098 151580 191104 151592
rect 191156 151580 191162 151632
rect 191926 151580 191932 151632
rect 191984 151620 191990 151632
rect 195946 151620 195974 151728
rect 265618 151716 265624 151728
rect 265676 151716 265682 151768
rect 316586 151716 316592 151768
rect 316644 151756 316650 151768
rect 316788 151756 316816 151796
rect 325970 151784 325976 151796
rect 326028 151784 326034 151836
rect 326062 151784 326068 151836
rect 326120 151824 326126 151836
rect 328546 151824 328552 151836
rect 326120 151796 328552 151824
rect 326120 151784 326126 151796
rect 328546 151784 328552 151796
rect 328604 151784 328610 151836
rect 332686 151784 332692 151836
rect 332744 151824 332750 151836
rect 334342 151824 334348 151836
rect 332744 151796 334348 151824
rect 332744 151784 332750 151796
rect 334342 151784 334348 151796
rect 334400 151784 334406 151836
rect 337838 151784 337844 151836
rect 337896 151824 337902 151836
rect 338758 151824 338764 151836
rect 337896 151796 338764 151824
rect 337896 151784 337902 151796
rect 338758 151784 338764 151796
rect 338816 151784 338822 151836
rect 340846 151824 340874 151864
rect 344922 151852 344928 151904
rect 344980 151892 344986 151904
rect 349706 151892 349712 151904
rect 344980 151864 349712 151892
rect 344980 151852 344986 151864
rect 349706 151852 349712 151864
rect 349764 151852 349770 151904
rect 393406 151892 393412 151904
rect 373966 151864 393412 151892
rect 347130 151824 347136 151836
rect 340846 151796 347136 151824
rect 347130 151784 347136 151796
rect 347188 151784 347194 151836
rect 347222 151784 347228 151836
rect 347280 151824 347286 151836
rect 355318 151824 355324 151836
rect 347280 151796 355324 151824
rect 347280 151784 347286 151796
rect 355318 151784 355324 151796
rect 355376 151784 355382 151836
rect 358906 151784 358912 151836
rect 358964 151824 358970 151836
rect 373966 151824 373994 151864
rect 393406 151852 393412 151864
rect 393464 151852 393470 151904
rect 396442 151852 396448 151904
rect 396500 151892 396506 151904
rect 402974 151892 402980 151904
rect 396500 151864 402980 151892
rect 396500 151852 396506 151864
rect 402974 151852 402980 151864
rect 403032 151852 403038 151904
rect 415854 151892 415860 151904
rect 403084 151864 415860 151892
rect 358964 151796 373994 151824
rect 358964 151784 358970 151796
rect 398834 151784 398840 151836
rect 398892 151824 398898 151836
rect 398892 151796 402192 151824
rect 398892 151784 398898 151796
rect 316644 151728 316816 151756
rect 402164 151756 402192 151796
rect 402238 151784 402244 151836
rect 402296 151824 402302 151836
rect 403084 151824 403112 151864
rect 415854 151852 415860 151864
rect 415912 151852 415918 151904
rect 420178 151852 420184 151904
rect 420236 151892 420242 151904
rect 434438 151892 434444 151904
rect 420236 151864 434444 151892
rect 420236 151852 420242 151864
rect 434438 151852 434444 151864
rect 434496 151852 434502 151904
rect 449986 151852 449992 151904
rect 450044 151892 450050 151904
rect 451826 151892 451832 151904
rect 450044 151864 451832 151892
rect 450044 151852 450050 151864
rect 451826 151852 451832 151864
rect 451884 151852 451890 151904
rect 459554 151852 459560 151904
rect 459612 151892 459618 151904
rect 462038 151892 462044 151904
rect 459612 151864 462044 151892
rect 459612 151852 459618 151864
rect 462038 151852 462044 151864
rect 462096 151852 462102 151904
rect 477678 151852 477684 151904
rect 477736 151892 477742 151904
rect 480714 151892 480720 151904
rect 477736 151864 480720 151892
rect 477736 151852 477742 151864
rect 480714 151852 480720 151864
rect 480772 151852 480778 151904
rect 488902 151852 488908 151904
rect 488960 151892 488966 151904
rect 490282 151892 490288 151904
rect 488960 151864 490288 151892
rect 488960 151852 488966 151864
rect 490282 151852 490288 151864
rect 490340 151852 490346 151904
rect 410702 151824 410708 151836
rect 402296 151796 403112 151824
rect 403176 151796 410708 151824
rect 402296 151784 402302 151796
rect 403176 151756 403204 151796
rect 410702 151784 410708 151796
rect 410760 151784 410766 151836
rect 416682 151784 416688 151836
rect 416740 151824 416746 151836
rect 424226 151824 424232 151836
rect 416740 151796 424232 151824
rect 416740 151784 416746 151796
rect 424226 151784 424232 151796
rect 424284 151784 424290 151836
rect 402164 151728 403204 151756
rect 316644 151716 316650 151728
rect 196066 151648 196072 151700
rect 196124 151688 196130 151700
rect 268838 151688 268844 151700
rect 196124 151660 268844 151688
rect 196124 151648 196130 151660
rect 268838 151648 268844 151660
rect 268896 151648 268902 151700
rect 191984 151592 195974 151620
rect 191984 151580 191990 151592
rect 198550 151580 198556 151632
rect 198608 151620 198614 151632
rect 270770 151620 270776 151632
rect 198608 151592 270776 151620
rect 198608 151580 198614 151592
rect 270770 151580 270776 151592
rect 270828 151580 270834 151632
rect 91002 151512 91008 151564
rect 91060 151552 91066 151564
rect 188522 151552 188528 151564
rect 91060 151524 188528 151552
rect 91060 151512 91066 151524
rect 188522 151512 188528 151524
rect 188580 151512 188586 151564
rect 188614 151512 188620 151564
rect 188672 151552 188678 151564
rect 263042 151552 263048 151564
rect 188672 151524 263048 151552
rect 188672 151512 188678 151524
rect 263042 151512 263048 151524
rect 263100 151512 263106 151564
rect 82722 151444 82728 151496
rect 82780 151484 82786 151496
rect 181438 151484 181444 151496
rect 82780 151456 181444 151484
rect 82780 151444 82786 151456
rect 181438 151444 181444 151456
rect 181496 151444 181502 151496
rect 181990 151444 181996 151496
rect 182048 151484 182054 151496
rect 257890 151484 257896 151496
rect 182048 151456 257896 151484
rect 182048 151444 182054 151456
rect 257890 151444 257896 151456
rect 257948 151444 257954 151496
rect 74258 151376 74264 151428
rect 74316 151416 74322 151428
rect 175550 151416 175556 151428
rect 74316 151388 175556 151416
rect 74316 151376 74322 151388
rect 175550 151376 175556 151388
rect 175608 151376 175614 151428
rect 175642 151376 175648 151428
rect 175700 151416 175706 151428
rect 191006 151416 191012 151428
rect 175700 151388 191012 151416
rect 175700 151376 175706 151388
rect 191006 151376 191012 151388
rect 191064 151376 191070 151428
rect 191098 151376 191104 151428
rect 191156 151416 191162 151428
rect 261110 151416 261116 151428
rect 191156 151388 261116 151416
rect 191156 151376 191162 151388
rect 261110 151376 261116 151388
rect 261168 151376 261174 151428
rect 71682 151308 71688 151360
rect 71740 151348 71746 151360
rect 173802 151348 173808 151360
rect 71740 151320 173808 151348
rect 71740 151308 71746 151320
rect 173802 151308 173808 151320
rect 173860 151308 173866 151360
rect 175182 151308 175188 151360
rect 175240 151348 175246 151360
rect 252738 151348 252744 151360
rect 175240 151320 252744 151348
rect 175240 151308 175246 151320
rect 252738 151308 252744 151320
rect 252796 151308 252802 151360
rect 24670 151240 24676 151292
rect 24728 151280 24734 151292
rect 137830 151280 137836 151292
rect 24728 151252 137836 151280
rect 24728 151240 24734 151252
rect 137830 151240 137836 151252
rect 137888 151240 137894 151292
rect 155678 151240 155684 151292
rect 155736 151280 155742 151292
rect 237374 151280 237380 151292
rect 155736 151252 237380 151280
rect 155736 151240 155742 151252
rect 237374 151240 237380 151252
rect 237432 151240 237438 151292
rect 263502 151240 263508 151292
rect 263560 151280 263566 151292
rect 320174 151280 320180 151292
rect 263560 151252 320180 151280
rect 263560 151240 263566 151252
rect 320174 151240 320180 151252
rect 320232 151240 320238 151292
rect 19242 151172 19248 151224
rect 19300 151212 19306 151224
rect 132678 151212 132684 151224
rect 19300 151184 132684 151212
rect 19300 151172 19306 151184
rect 132678 151172 132684 151184
rect 132736 151172 132742 151224
rect 137278 151172 137284 151224
rect 137336 151212 137342 151224
rect 220630 151212 220636 151224
rect 137336 151184 220636 151212
rect 137336 151172 137342 151184
rect 220630 151172 220636 151184
rect 220688 151172 220694 151224
rect 256418 151172 256424 151224
rect 256476 151212 256482 151224
rect 315022 151212 315028 151224
rect 256476 151184 315028 151212
rect 256476 151172 256482 151184
rect 315022 151172 315028 151184
rect 315080 151172 315086 151224
rect 12342 151104 12348 151156
rect 12400 151144 12406 151156
rect 127526 151144 127532 151156
rect 12400 151116 127532 151144
rect 12400 151104 12406 151116
rect 127526 151104 127532 151116
rect 127584 151104 127590 151156
rect 135162 151104 135168 151156
rect 135220 151144 135226 151156
rect 221918 151144 221924 151156
rect 135220 151116 221924 151144
rect 135220 151104 135226 151116
rect 221918 151104 221924 151116
rect 221976 151104 221982 151156
rect 246390 151104 246396 151156
rect 246448 151144 246454 151156
rect 307294 151144 307300 151156
rect 246448 151116 307300 151144
rect 246448 151104 246454 151116
rect 307294 151104 307300 151116
rect 307352 151104 307358 151156
rect 5350 151036 5356 151088
rect 5408 151076 5414 151088
rect 123018 151076 123024 151088
rect 5408 151048 123024 151076
rect 5408 151036 5414 151048
rect 123018 151036 123024 151048
rect 123076 151036 123082 151088
rect 127986 151036 127992 151088
rect 128044 151076 128050 151088
rect 216766 151076 216772 151088
rect 128044 151048 216772 151076
rect 128044 151036 128050 151048
rect 216766 151036 216772 151048
rect 216824 151036 216830 151088
rect 223482 151036 223488 151088
rect 223540 151076 223546 151088
rect 289354 151076 289360 151088
rect 223540 151048 289360 151076
rect 223540 151036 223546 151048
rect 289354 151036 289360 151048
rect 289412 151036 289418 151088
rect 102042 150968 102048 151020
rect 102100 151008 102106 151020
rect 196250 151008 196256 151020
rect 102100 150980 196256 151008
rect 102100 150968 102106 150980
rect 196250 150968 196256 150980
rect 196308 150968 196314 151020
rect 199378 150968 199384 151020
rect 199436 151008 199442 151020
rect 271414 151008 271420 151020
rect 199436 150980 271420 151008
rect 199436 150968 199442 150980
rect 271414 150968 271420 150980
rect 271472 150968 271478 151020
rect 108942 150900 108948 150952
rect 109000 150940 109006 150952
rect 201402 150940 201408 150952
rect 109000 150912 201408 150940
rect 109000 150900 109006 150912
rect 201402 150900 201408 150912
rect 201460 150900 201466 150952
rect 202690 150900 202696 150952
rect 202748 150940 202754 150952
rect 273898 150940 273904 150952
rect 202748 150912 273904 150940
rect 202748 150900 202754 150912
rect 273898 150900 273904 150912
rect 273956 150900 273962 150952
rect 43898 150832 43904 150884
rect 43956 150872 43962 150884
rect 116854 150872 116860 150884
rect 43956 150844 116860 150872
rect 43956 150832 43962 150844
rect 116854 150832 116860 150844
rect 116912 150832 116918 150884
rect 206554 150872 206560 150884
rect 117056 150844 206560 150872
rect 95510 150764 95516 150816
rect 95568 150804 95574 150816
rect 110322 150804 110328 150816
rect 95568 150776 110328 150804
rect 95568 150764 95574 150776
rect 110322 150764 110328 150776
rect 110380 150764 110386 150816
rect 115750 150764 115756 150816
rect 115808 150804 115814 150816
rect 117056 150804 117084 150844
rect 206554 150832 206560 150844
rect 206612 150832 206618 150884
rect 209406 150832 209412 150884
rect 209464 150872 209470 150884
rect 279050 150872 279056 150884
rect 209464 150844 279056 150872
rect 209464 150832 209470 150844
rect 279050 150832 279056 150844
rect 279108 150832 279114 150884
rect 115808 150776 117084 150804
rect 115808 150764 115814 150776
rect 118602 150764 118608 150816
rect 118660 150804 118666 150816
rect 209130 150804 209136 150816
rect 118660 150776 209136 150804
rect 118660 150764 118666 150776
rect 209130 150764 209136 150776
rect 209188 150764 209194 150816
rect 92014 150696 92020 150748
rect 92072 150736 92078 150748
rect 111518 150736 111524 150748
rect 92072 150708 111524 150736
rect 92072 150696 92078 150708
rect 111518 150696 111524 150708
rect 111576 150696 111582 150748
rect 121362 150696 121368 150748
rect 121420 150736 121426 150748
rect 211614 150736 211620 150748
rect 121420 150708 211620 150736
rect 121420 150696 121426 150708
rect 211614 150696 211620 150708
rect 211672 150696 211678 150748
rect 88610 150628 88616 150680
rect 88668 150668 88674 150680
rect 111426 150668 111432 150680
rect 88668 150640 111432 150668
rect 88668 150628 88674 150640
rect 111426 150628 111432 150640
rect 111484 150628 111490 150680
rect 116762 150628 116768 150680
rect 116820 150668 116826 150680
rect 116820 150640 118694 150668
rect 116820 150628 116826 150640
rect 85206 150560 85212 150612
rect 85264 150600 85270 150612
rect 117222 150600 117228 150612
rect 85264 150572 117228 150600
rect 85264 150560 85270 150572
rect 117222 150560 117228 150572
rect 117280 150560 117286 150612
rect 50798 150492 50804 150544
rect 50856 150532 50862 150544
rect 116946 150532 116952 150544
rect 50856 150504 116952 150532
rect 50856 150492 50862 150504
rect 116946 150492 116952 150504
rect 117004 150492 117010 150544
rect 118666 150532 118694 150640
rect 168282 150628 168288 150680
rect 168340 150668 168346 150680
rect 247586 150668 247592 150680
rect 168340 150640 247592 150668
rect 168340 150628 168346 150640
rect 247586 150628 247592 150640
rect 247644 150628 247650 150680
rect 164970 150560 164976 150612
rect 165028 150600 165034 150612
rect 245010 150600 245016 150612
rect 165028 150572 245016 150600
rect 165028 150560 165034 150572
rect 245010 150560 245016 150572
rect 245068 150560 245074 150612
rect 194962 150532 194968 150544
rect 118666 150504 194968 150532
rect 194962 150492 194968 150504
rect 195020 150492 195026 150544
rect 195054 150492 195060 150544
rect 195112 150532 195118 150544
rect 238662 150532 238668 150544
rect 195112 150504 238668 150532
rect 195112 150492 195118 150504
rect 238662 150492 238668 150504
rect 238720 150492 238726 150544
rect 98914 150424 98920 150476
rect 98972 150464 98978 150476
rect 111242 150464 111248 150476
rect 98972 150436 111248 150464
rect 98972 150424 98978 150436
rect 111242 150424 111248 150436
rect 111300 150424 111306 150476
rect 117130 150424 117136 150476
rect 117188 150464 117194 150476
rect 179598 150464 179604 150476
rect 117188 150436 179604 150464
rect 117188 150424 117194 150436
rect 179598 150424 179604 150436
rect 179656 150424 179662 150476
rect 180058 150424 180064 150476
rect 180116 150464 180122 150476
rect 251450 150464 251456 150476
rect 180116 150436 251456 150464
rect 180116 150424 180122 150436
rect 251450 150424 251456 150436
rect 251508 150424 251514 150476
rect 78306 150356 78312 150408
rect 78364 150396 78370 150408
rect 114094 150396 114100 150408
rect 78364 150368 114100 150396
rect 78364 150356 78370 150368
rect 114094 150356 114100 150368
rect 114152 150356 114158 150408
rect 74810 150288 74816 150340
rect 74868 150328 74874 150340
rect 114002 150328 114008 150340
rect 74868 150300 114008 150328
rect 74868 150288 74874 150300
rect 114002 150288 114008 150300
rect 114060 150288 114066 150340
rect 71406 150220 71412 150272
rect 71464 150260 71470 150272
rect 115198 150260 115204 150272
rect 71464 150232 115204 150260
rect 71464 150220 71470 150232
rect 115198 150220 115204 150232
rect 115256 150220 115262 150272
rect 102594 150152 102600 150204
rect 102652 150192 102658 150204
rect 116026 150192 116032 150204
rect 102652 150164 116032 150192
rect 102652 150152 102658 150164
rect 116026 150152 116032 150164
rect 116084 150152 116090 150204
rect 147674 150152 147680 150204
rect 147732 150192 147738 150204
rect 148824 150192 148830 150204
rect 147732 150164 148830 150192
rect 147732 150152 147738 150164
rect 148824 150152 148830 150164
rect 148882 150152 148888 150204
rect 218238 150152 218244 150204
rect 218296 150192 218302 150204
rect 219388 150192 219394 150204
rect 218296 150164 219394 150192
rect 218296 150152 218302 150164
rect 219388 150152 219394 150164
rect 219446 150152 219452 150204
rect 265158 150152 265164 150204
rect 265216 150192 265222 150204
rect 266308 150192 266314 150204
rect 265216 150164 266314 150192
rect 265216 150152 265222 150164
rect 266308 150152 266314 150164
rect 266366 150152 266372 150204
rect 292482 150152 292488 150204
rect 292540 150192 292546 150204
rect 293908 150192 293914 150204
rect 292540 150164 293914 150192
rect 292540 150152 292546 150164
rect 293908 150152 293914 150164
rect 293966 150152 293972 150204
rect 394878 150152 394884 150204
rect 394936 150192 394942 150204
rect 396028 150192 396034 150204
rect 394936 150164 396034 150192
rect 394936 150152 394942 150164
rect 396028 150152 396034 150164
rect 396086 150152 396092 150204
rect 451366 150152 451372 150204
rect 451424 150192 451430 150204
rect 452516 150192 452522 150204
rect 451424 150164 452522 150192
rect 451424 150152 451430 150164
rect 452516 150152 452522 150164
rect 452574 150152 452580 150204
rect 455414 150152 455420 150204
rect 455472 150192 455478 150204
rect 456380 150192 456386 150204
rect 455472 150164 456386 150192
rect 455472 150152 455478 150164
rect 456380 150152 456386 150164
rect 456438 150152 456444 150204
rect 456794 150152 456800 150204
rect 456852 150192 456858 150204
rect 457668 150192 457674 150204
rect 456852 150164 457674 150192
rect 456852 150152 456858 150164
rect 457668 150152 457674 150164
rect 457726 150152 457732 150204
rect 462314 150152 462320 150204
rect 462372 150192 462378 150204
rect 463372 150192 463378 150204
rect 462372 150164 463378 150192
rect 462372 150152 462378 150164
rect 463372 150152 463378 150164
rect 463430 150152 463436 150204
rect 468018 150152 468024 150204
rect 468076 150192 468082 150204
rect 469168 150192 469174 150204
rect 468076 150164 469174 150192
rect 468076 150152 468082 150164
rect 469168 150152 469174 150164
rect 469226 150152 469232 150204
rect 471974 150152 471980 150204
rect 472032 150192 472038 150204
rect 473032 150192 473038 150204
rect 472032 150164 473038 150192
rect 472032 150152 472038 150164
rect 473032 150152 473038 150164
rect 473090 150152 473096 150204
rect 496906 150152 496912 150204
rect 496964 150192 496970 150204
rect 498056 150192 498062 150204
rect 496964 150164 498062 150192
rect 496964 150152 496970 150164
rect 498056 150152 498062 150164
rect 498114 150152 498120 150204
rect 500954 150152 500960 150204
rect 501012 150192 501018 150204
rect 501920 150192 501926 150204
rect 501012 150164 501926 150192
rect 501012 150152 501018 150164
rect 501920 150152 501926 150164
rect 501978 150152 501984 150204
rect 68002 150084 68008 150136
rect 68060 150084 68066 150136
rect 92474 150084 92480 150136
rect 92532 150124 92538 150136
rect 117130 150124 117136 150136
rect 92532 150096 117136 150124
rect 92532 150084 92538 150096
rect 117130 150084 117136 150096
rect 117188 150084 117194 150136
rect 202736 150084 202742 150136
rect 202794 150084 202800 150136
rect 292390 150084 292396 150136
rect 292448 150124 292454 150136
rect 299060 150124 299066 150136
rect 292448 150096 299066 150124
rect 292448 150084 292454 150096
rect 299060 150084 299066 150096
rect 299118 150084 299124 150136
rect 68020 150056 68048 150084
rect 111058 150056 111064 150068
rect 68020 150028 111064 150056
rect 111058 150016 111064 150028
rect 111116 150016 111122 150068
rect 111610 150016 111616 150068
rect 111668 150056 111674 150068
rect 202754 150056 202782 150084
rect 111668 150028 202782 150056
rect 111668 150016 111674 150028
rect 111150 148996 111156 149048
rect 111208 149036 111214 149048
rect 116118 149036 116124 149048
rect 111208 149008 116124 149036
rect 111208 148996 111214 149008
rect 116118 148996 116124 149008
rect 116176 148996 116182 149048
rect 116670 146956 116676 147008
rect 116728 146996 116734 147008
rect 117038 146996 117044 147008
rect 116728 146968 117044 146996
rect 116728 146956 116734 146968
rect 117038 146956 117044 146968
rect 117096 146956 117102 147008
rect 111242 143488 111248 143540
rect 111300 143528 111306 143540
rect 116118 143528 116124 143540
rect 111300 143500 116124 143528
rect 111300 143488 111306 143500
rect 116118 143488 116124 143500
rect 116176 143488 116182 143540
rect 111058 143148 111064 143200
rect 111116 143188 111122 143200
rect 111426 143188 111432 143200
rect 111116 143160 111432 143188
rect 111116 143148 111122 143160
rect 111426 143148 111432 143160
rect 111484 143148 111490 143200
rect 111518 140700 111524 140752
rect 111576 140740 111582 140752
rect 116118 140740 116124 140752
rect 111576 140712 116124 140740
rect 111576 140700 111582 140712
rect 116118 140700 116124 140712
rect 116176 140700 116182 140752
rect 111334 137912 111340 137964
rect 111392 137952 111398 137964
rect 116118 137952 116124 137964
rect 111392 137924 116124 137952
rect 111392 137912 111398 137924
rect 116118 137912 116124 137924
rect 116176 137912 116182 137964
rect 114094 132132 114100 132184
rect 114152 132172 114158 132184
rect 115934 132172 115940 132184
rect 114152 132144 115940 132172
rect 114152 132132 114158 132144
rect 115934 132132 115940 132144
rect 115992 132132 115998 132184
rect 114002 131044 114008 131096
rect 114060 131084 114066 131096
rect 115934 131084 115940 131096
rect 114060 131056 115940 131084
rect 114060 131044 114066 131056
rect 115934 131044 115940 131056
rect 115992 131044 115998 131096
rect 111150 126896 111156 126948
rect 111208 126936 111214 126948
rect 116118 126936 116124 126948
rect 111208 126908 116124 126936
rect 111208 126896 111214 126908
rect 116118 126896 116124 126908
rect 116176 126896 116182 126948
rect 112898 124108 112904 124160
rect 112956 124148 112962 124160
rect 116118 124148 116124 124160
rect 112956 124120 116124 124148
rect 112956 124108 112962 124120
rect 116118 124108 116124 124120
rect 116176 124108 116182 124160
rect 112714 122748 112720 122800
rect 112772 122788 112778 122800
rect 116118 122788 116124 122800
rect 112772 122760 116124 122788
rect 112772 122748 112778 122760
rect 116118 122748 116124 122760
rect 116176 122748 116182 122800
rect 112530 121388 112536 121440
rect 112588 121428 112594 121440
rect 116118 121428 116124 121440
rect 112588 121400 116124 121428
rect 112588 121388 112594 121400
rect 116118 121388 116124 121400
rect 116176 121388 116182 121440
rect 112438 107584 112444 107636
rect 112496 107624 112502 107636
rect 116118 107624 116124 107636
rect 112496 107596 116124 107624
rect 112496 107584 112502 107596
rect 116118 107584 116124 107596
rect 116176 107584 116182 107636
rect 111610 104796 111616 104848
rect 111668 104836 111674 104848
rect 116118 104836 116124 104848
rect 111668 104808 116124 104836
rect 111668 104796 111674 104808
rect 116118 104796 116124 104808
rect 116176 104796 116182 104848
rect 111426 102076 111432 102128
rect 111484 102116 111490 102128
rect 115934 102116 115940 102128
rect 111484 102088 115940 102116
rect 111484 102076 111490 102088
rect 115934 102076 115940 102088
rect 115992 102076 115998 102128
rect 111242 96568 111248 96620
rect 111300 96608 111306 96620
rect 116118 96608 116124 96620
rect 111300 96580 116124 96608
rect 111300 96568 111306 96580
rect 116118 96568 116124 96580
rect 116176 96568 116182 96620
rect 111058 93780 111064 93832
rect 111116 93820 111122 93832
rect 116118 93820 116124 93832
rect 111116 93792 116124 93820
rect 111116 93780 111122 93792
rect 116118 93780 116124 93792
rect 116176 93780 116182 93832
rect 113818 88272 113824 88324
rect 113876 88312 113882 88324
rect 115934 88312 115940 88324
rect 113876 88284 115940 88312
rect 113876 88272 113882 88284
rect 115934 88272 115940 88284
rect 115992 88272 115998 88324
rect 113910 86912 113916 86964
rect 113968 86952 113974 86964
rect 116394 86952 116400 86964
rect 113968 86924 116400 86952
rect 113968 86912 113974 86924
rect 116394 86912 116400 86924
rect 116452 86912 116458 86964
rect 114002 83920 114008 83972
rect 114060 83960 114066 83972
rect 116578 83960 116584 83972
rect 114060 83932 116584 83960
rect 114060 83920 114066 83932
rect 116578 83920 116584 83932
rect 116636 83920 116642 83972
rect 114094 82764 114100 82816
rect 114152 82804 114158 82816
rect 116302 82804 116308 82816
rect 114152 82776 116308 82804
rect 114152 82764 114158 82776
rect 116302 82764 116308 82776
rect 116360 82764 116366 82816
rect 114186 79976 114192 80028
rect 114244 80016 114250 80028
rect 115934 80016 115940 80028
rect 114244 79988 115940 80016
rect 114244 79976 114250 79988
rect 115934 79976 115940 79988
rect 115992 79976 115998 80028
rect 114278 78616 114284 78668
rect 114336 78656 114342 78668
rect 116210 78656 116216 78668
rect 114336 78628 116216 78656
rect 114336 78616 114342 78628
rect 116210 78616 116216 78628
rect 116268 78616 116274 78668
rect 114186 71748 114192 71800
rect 114244 71788 114250 71800
rect 116578 71788 116584 71800
rect 114244 71760 116584 71788
rect 114244 71748 114250 71760
rect 116578 71748 116584 71760
rect 116636 71748 116642 71800
rect 114094 69028 114100 69080
rect 114152 69068 114158 69080
rect 116302 69068 116308 69080
rect 114152 69040 116308 69068
rect 114152 69028 114158 69040
rect 116302 69028 116308 69040
rect 116360 69028 116366 69080
rect 114002 67600 114008 67652
rect 114060 67640 114066 67652
rect 116118 67640 116124 67652
rect 114060 67612 116124 67640
rect 114060 67600 114066 67612
rect 116118 67600 116124 67612
rect 116176 67600 116182 67652
rect 113910 66240 113916 66292
rect 113968 66280 113974 66292
rect 116578 66280 116584 66292
rect 113968 66252 116584 66280
rect 113968 66240 113974 66252
rect 116578 66240 116584 66252
rect 116636 66240 116642 66292
rect 113358 64676 113364 64728
rect 113416 64716 113422 64728
rect 116578 64716 116584 64728
rect 113416 64688 116584 64716
rect 113416 64676 113422 64688
rect 116578 64676 116584 64688
rect 116636 64676 116642 64728
rect 113818 63520 113824 63572
rect 113876 63560 113882 63572
rect 116210 63560 116216 63572
rect 113876 63532 116216 63560
rect 113876 63520 113882 63532
rect 116210 63520 116216 63532
rect 116268 63520 116274 63572
rect 112438 62092 112444 62144
rect 112496 62132 112502 62144
rect 116118 62132 116124 62144
rect 112496 62104 116124 62132
rect 112496 62092 112502 62104
rect 116118 62092 116124 62104
rect 116176 62092 116182 62144
rect 112530 44140 112536 44192
rect 112588 44180 112594 44192
rect 116118 44180 116124 44192
rect 112588 44152 116124 44180
rect 112588 44140 112594 44152
rect 116118 44140 116124 44152
rect 116176 44140 116182 44192
rect 112622 34484 112628 34536
rect 112680 34524 112686 34536
rect 115934 34524 115940 34536
rect 112680 34496 115940 34524
rect 112680 34484 112686 34496
rect 115934 34484 115940 34496
rect 115992 34484 115998 34536
rect 114094 33124 114100 33176
rect 114152 33164 114158 33176
rect 115934 33164 115940 33176
rect 114152 33136 115940 33164
rect 114152 33124 114158 33136
rect 115934 33124 115940 33136
rect 115992 33124 115998 33176
rect 112714 28976 112720 29028
rect 112772 29016 112778 29028
rect 116118 29016 116124 29028
rect 112772 28988 116124 29016
rect 112772 28976 112778 28988
rect 116118 28976 116124 28988
rect 116176 28976 116182 29028
rect 112806 24828 112812 24880
rect 112864 24868 112870 24880
rect 116118 24868 116124 24880
rect 112864 24840 116124 24868
rect 112864 24828 112870 24840
rect 116118 24828 116124 24840
rect 116176 24828 116182 24880
rect 114002 23468 114008 23520
rect 114060 23508 114066 23520
rect 115934 23508 115940 23520
rect 114060 23480 115940 23508
rect 114060 23468 114066 23480
rect 115934 23468 115940 23480
rect 115992 23468 115998 23520
rect 112898 22108 112904 22160
rect 112956 22148 112962 22160
rect 116118 22148 116124 22160
rect 112956 22120 116124 22148
rect 112956 22108 112962 22120
rect 116118 22108 116124 22120
rect 116176 22108 116182 22160
rect 116394 11704 116400 11756
rect 116452 11744 116458 11756
rect 116854 11744 116860 11756
rect 116452 11716 116860 11744
rect 116452 11704 116458 11716
rect 116854 11704 116860 11716
rect 116912 11704 116918 11756
rect 116026 11636 116032 11688
rect 116084 11676 116090 11688
rect 117038 11676 117044 11688
rect 116084 11648 117044 11676
rect 116084 11636 116090 11648
rect 117038 11636 117044 11648
rect 117096 11636 117102 11688
rect 111150 5516 111156 5568
rect 111208 5556 111214 5568
rect 115934 5556 115940 5568
rect 111208 5528 115940 5556
rect 111208 5516 111214 5528
rect 115934 5516 115940 5528
rect 115992 5516 115998 5568
rect 111794 4156 111800 4208
rect 111852 4196 111858 4208
rect 116118 4196 116124 4208
rect 111852 4168 116124 4196
rect 111852 4156 111858 4168
rect 116118 4156 116124 4168
rect 116176 4156 116182 4208
rect 111058 2796 111064 2848
rect 111116 2836 111122 2848
rect 111116 2808 143672 2836
rect 111116 2796 111122 2808
rect 143644 2508 143672 2808
rect 425808 2808 443684 2836
rect 425808 2508 425836 2808
rect 443656 2508 443684 2808
rect 143626 2456 143632 2508
rect 143684 2456 143690 2508
rect 425790 2456 425796 2508
rect 425848 2456 425854 2508
rect 443638 2456 443644 2508
rect 443696 2456 443702 2508
rect 102686 1912 102692 1964
rect 102744 1952 102750 1964
rect 116578 1952 116584 1964
rect 102744 1924 116584 1952
rect 102744 1912 102750 1924
rect 116578 1912 116584 1924
rect 116636 1912 116642 1964
rect 92658 1844 92664 1896
rect 92716 1884 92722 1896
rect 94406 1884 94412 1896
rect 92716 1856 94412 1884
rect 92716 1844 92722 1856
rect 94406 1844 94412 1856
rect 94464 1844 94470 1896
rect 95970 1844 95976 1896
rect 96028 1884 96034 1896
rect 96028 1856 105952 1884
rect 96028 1844 96034 1856
rect 89346 1776 89352 1828
rect 89404 1816 89410 1828
rect 105814 1816 105820 1828
rect 89404 1788 105820 1816
rect 89404 1776 89410 1788
rect 105814 1776 105820 1788
rect 105872 1776 105878 1828
rect 105924 1816 105952 1856
rect 105998 1844 106004 1896
rect 106056 1884 106062 1896
rect 109678 1884 109684 1896
rect 106056 1856 109684 1884
rect 106056 1844 106062 1856
rect 109678 1844 109684 1856
rect 109736 1844 109742 1896
rect 109034 1816 109040 1828
rect 105924 1788 109040 1816
rect 109034 1776 109040 1788
rect 109092 1776 109098 1828
rect 109310 1776 109316 1828
rect 109368 1816 109374 1828
rect 112438 1816 112444 1828
rect 109368 1788 112444 1816
rect 109368 1776 109374 1788
rect 112438 1776 112444 1788
rect 112496 1776 112502 1828
rect 65978 1708 65984 1760
rect 66036 1748 66042 1760
rect 88886 1748 88892 1760
rect 66036 1720 88892 1748
rect 66036 1708 66042 1720
rect 88886 1708 88892 1720
rect 88944 1708 88950 1760
rect 99374 1708 99380 1760
rect 99432 1748 99438 1760
rect 116670 1748 116676 1760
rect 99432 1720 116676 1748
rect 99432 1708 99438 1720
rect 116670 1708 116676 1720
rect 116728 1708 116734 1760
rect 86034 1640 86040 1692
rect 86092 1680 86098 1692
rect 86092 1652 105768 1680
rect 86092 1640 86098 1652
rect 82630 1572 82636 1624
rect 82688 1612 82694 1624
rect 105630 1612 105636 1624
rect 82688 1584 105636 1612
rect 82688 1572 82694 1584
rect 105630 1572 105636 1584
rect 105688 1572 105694 1624
rect 72694 1504 72700 1556
rect 72752 1544 72758 1556
rect 100294 1544 100300 1556
rect 72752 1516 100300 1544
rect 72752 1504 72758 1516
rect 100294 1504 100300 1516
rect 100352 1504 100358 1556
rect 105740 1544 105768 1652
rect 105814 1640 105820 1692
rect 105872 1640 105878 1692
rect 105906 1640 105912 1692
rect 105964 1680 105970 1692
rect 108942 1680 108948 1692
rect 105964 1652 108948 1680
rect 105964 1640 105970 1652
rect 108942 1640 108948 1652
rect 109000 1640 109006 1692
rect 109034 1640 109040 1692
rect 109092 1680 109098 1692
rect 109770 1680 109776 1692
rect 109092 1652 109776 1680
rect 109092 1640 109098 1652
rect 109770 1640 109776 1652
rect 109828 1640 109834 1692
rect 105832 1612 105860 1640
rect 109862 1612 109868 1624
rect 105832 1584 109868 1612
rect 109862 1572 109868 1584
rect 109920 1572 109926 1624
rect 109954 1544 109960 1556
rect 105740 1516 109960 1544
rect 109954 1504 109960 1516
rect 110012 1504 110018 1556
rect 110138 1504 110144 1556
rect 110196 1544 110202 1556
rect 193582 1544 193588 1556
rect 110196 1516 193588 1544
rect 110196 1504 110202 1516
rect 193582 1504 193588 1516
rect 193640 1504 193646 1556
rect 32674 1436 32680 1488
rect 32732 1476 32738 1488
rect 116394 1476 116400 1488
rect 32732 1448 116400 1476
rect 32732 1436 32738 1448
rect 116394 1436 116400 1448
rect 116452 1436 116458 1488
rect 29270 1368 29276 1420
rect 29328 1408 29334 1420
rect 115934 1408 115940 1420
rect 29328 1380 115940 1408
rect 29328 1368 29334 1380
rect 115934 1368 115940 1380
rect 115992 1368 115998 1420
rect 294782 1368 294788 1420
rect 294840 1408 294846 1420
rect 343634 1408 343640 1420
rect 294840 1380 343640 1408
rect 294840 1368 294846 1380
rect 343634 1368 343640 1380
rect 343692 1368 343698 1420
rect 491294 1368 491300 1420
rect 491352 1408 491358 1420
rect 493594 1408 493600 1420
rect 491352 1380 493600 1408
rect 491352 1368 491358 1380
rect 493594 1368 493600 1380
rect 493652 1368 493658 1420
rect 2682 1300 2688 1352
rect 2740 1340 2746 1352
rect 116118 1340 116124 1352
rect 2740 1312 116124 1340
rect 2740 1300 2746 1312
rect 116118 1300 116124 1312
rect 116176 1300 116182 1352
rect 5994 1232 6000 1284
rect 6052 1272 6058 1284
rect 111794 1272 111800 1284
rect 6052 1244 111800 1272
rect 6052 1232 6058 1244
rect 111794 1232 111800 1244
rect 111852 1232 111858 1284
rect 9306 1164 9312 1216
rect 9364 1204 9370 1216
rect 111150 1204 111156 1216
rect 9364 1176 111156 1204
rect 9364 1164 9370 1176
rect 111150 1164 111156 1176
rect 111208 1164 111214 1216
rect 35986 1096 35992 1148
rect 36044 1136 36050 1148
rect 112898 1136 112904 1148
rect 36044 1108 112904 1136
rect 36044 1096 36050 1108
rect 112898 1096 112904 1108
rect 112956 1096 112962 1148
rect 39298 1028 39304 1080
rect 39356 1068 39362 1080
rect 114002 1068 114008 1080
rect 39356 1040 114008 1068
rect 39356 1028 39362 1040
rect 114002 1028 114008 1040
rect 114060 1028 114066 1080
rect 42610 960 42616 1012
rect 42668 1000 42674 1012
rect 112806 1000 112812 1012
rect 42668 972 112812 1000
rect 42668 960 42674 972
rect 112806 960 112812 972
rect 112864 960 112870 1012
rect 46014 892 46020 944
rect 46072 932 46078 944
rect 46072 904 113174 932
rect 46072 892 46078 904
rect 49326 824 49332 876
rect 49384 864 49390 876
rect 112714 864 112720 876
rect 49384 836 112720 864
rect 49384 824 49390 836
rect 112714 824 112720 836
rect 112772 824 112778 876
rect 52638 756 52644 808
rect 52696 796 52702 808
rect 113146 796 113174 904
rect 115382 796 115388 808
rect 52696 768 108344 796
rect 113146 768 115388 796
rect 52696 756 52702 768
rect 59354 688 59360 740
rect 59412 728 59418 740
rect 108206 728 108212 740
rect 59412 700 108212 728
rect 59412 688 59418 700
rect 108206 688 108212 700
rect 108264 688 108270 740
rect 62666 620 62672 672
rect 62724 660 62730 672
rect 108316 660 108344 768
rect 115382 756 115388 768
rect 115440 756 115446 808
rect 108390 688 108396 740
rect 108448 728 108454 740
rect 114094 728 114100 740
rect 108448 700 114100 728
rect 108448 688 108454 700
rect 114094 688 114100 700
rect 114152 688 114158 740
rect 62724 632 108068 660
rect 108316 632 113174 660
rect 62724 620 62730 632
rect 69290 552 69296 604
rect 69348 592 69354 604
rect 108040 592 108068 632
rect 112622 592 112628 604
rect 69348 564 103652 592
rect 108040 564 112628 592
rect 69348 552 69354 564
rect 79318 484 79324 536
rect 79376 524 79382 536
rect 79376 496 103514 524
rect 79376 484 79382 496
rect 103486 388 103514 496
rect 103624 456 103652 564
rect 112622 552 112628 564
rect 112680 552 112686 604
rect 113146 592 113174 632
rect 115290 592 115296 604
rect 113146 564 115296 592
rect 115290 552 115296 564
rect 115348 552 115354 604
rect 115198 456 115204 468
rect 103624 428 115204 456
rect 115198 416 115204 428
rect 115256 416 115262 468
rect 112530 388 112536 400
rect 103486 360 112536 388
rect 112530 348 112536 360
rect 112588 348 112594 400
<< via1 >>
rect 31392 158516 31444 158568
rect 142712 158516 142764 158568
rect 96068 158448 96120 158500
rect 192392 158448 192444 158500
rect 89352 158380 89404 158432
rect 186688 158380 186740 158432
rect 82636 158312 82688 158364
rect 182088 158312 182140 158364
rect 75920 158244 75972 158296
rect 177028 158244 177080 158296
rect 69204 158176 69256 158228
rect 171876 158176 171928 158228
rect 72608 158108 72660 158160
rect 174452 158108 174504 158160
rect 65892 158040 65944 158092
rect 169300 158040 169352 158092
rect 62488 157972 62540 158024
rect 165988 157972 166040 158024
rect 59084 157904 59136 157956
rect 163872 157904 163924 157956
rect 55772 157836 55824 157888
rect 161664 157836 161716 157888
rect 52368 157768 52420 157820
rect 158996 157768 159048 157820
rect 45652 157700 45704 157752
rect 153752 157700 153804 157752
rect 49056 157632 49108 157684
rect 156328 157632 156380 157684
rect 42340 157564 42392 157616
rect 151268 157564 151320 157616
rect 38936 157496 38988 157548
rect 147680 157496 147732 157548
rect 35624 157428 35676 157480
rect 146208 157428 146260 157480
rect 102784 157360 102836 157412
rect 197544 157360 197596 157412
rect 47400 157292 47452 157344
rect 155132 157292 155184 157344
rect 156052 157292 156104 157344
rect 160284 157292 160336 157344
rect 161940 157292 161992 157344
rect 165436 157292 165488 157344
rect 172520 157292 172572 157344
rect 250812 157292 250864 157344
rect 43996 157224 44048 157276
rect 152556 157224 152608 157276
rect 155868 157224 155920 157276
rect 162584 157224 162636 157276
rect 171692 157224 171744 157276
rect 250168 157224 250220 157276
rect 37280 157156 37332 157208
rect 146852 157156 146904 157208
rect 40684 157088 40736 157140
rect 149980 157156 150032 157208
rect 152924 157156 152976 157208
rect 157708 157156 157760 157208
rect 161572 157156 161624 157208
rect 242440 157156 242492 157208
rect 148140 157088 148192 157140
rect 28080 157020 28132 157072
rect 140412 157020 140464 157072
rect 144828 157020 144880 157072
rect 23848 156952 23900 157004
rect 137100 156952 137152 157004
rect 143448 156952 143500 157004
rect 148140 156952 148192 157004
rect 21364 156884 21416 156936
rect 135352 156884 135404 156936
rect 138112 156884 138164 156936
rect 148324 157020 148376 157072
rect 151544 157020 151596 157072
rect 158260 157088 158312 157140
rect 239956 157088 240008 157140
rect 156420 156952 156472 157004
rect 232228 157020 232280 157072
rect 249800 157020 249852 157072
rect 309876 157020 309928 157072
rect 234804 156952 234856 157004
rect 243084 156952 243136 157004
rect 304724 156952 304776 157004
rect 14648 156816 14700 156868
rect 130108 156816 130160 156868
rect 141424 156816 141476 156868
rect 229560 156884 229612 156936
rect 239680 156884 239732 156936
rect 302240 156884 302292 156936
rect 7104 156748 7156 156800
rect 3700 156680 3752 156732
rect 121736 156680 121788 156732
rect 122748 156748 122800 156800
rect 143448 156748 143500 156800
rect 224132 156816 224184 156868
rect 226248 156816 226300 156868
rect 291936 156816 291988 156868
rect 226892 156748 226944 156800
rect 232964 156748 233016 156800
rect 297088 156748 297140 156800
rect 124312 156680 124364 156732
rect 131396 156680 131448 156732
rect 218244 156680 218296 156732
rect 219532 156680 219584 156732
rect 286784 156680 286836 156732
rect 388 156612 440 156664
rect 118976 156612 119028 156664
rect 124588 156612 124640 156664
rect 214196 156612 214248 156664
rect 216128 156612 216180 156664
rect 284116 156612 284168 156664
rect 50712 156544 50764 156596
rect 152924 156544 152976 156596
rect 153016 156544 153068 156596
rect 207848 156544 207900 156596
rect 54116 156476 54168 156528
rect 156052 156476 156104 156528
rect 156420 156476 156472 156528
rect 162124 156476 162176 156528
rect 60832 156408 60884 156460
rect 161940 156408 161992 156460
rect 70860 156340 70912 156392
rect 173072 156476 173124 156528
rect 174544 156476 174596 156528
rect 178040 156476 178092 156528
rect 179236 156476 179288 156528
rect 255964 156476 256016 156528
rect 162584 156408 162636 156460
rect 176200 156408 176252 156460
rect 176292 156408 176344 156460
rect 178960 156408 179012 156460
rect 183376 156408 183428 156460
rect 259184 156408 259236 156460
rect 321100 156408 321152 156460
rect 327264 156408 327316 156460
rect 162492 156340 162544 156392
rect 175832 156340 175884 156392
rect 78404 156272 78456 156324
rect 175924 156272 175976 156324
rect 181168 156340 181220 156392
rect 185124 156340 185176 156392
rect 260012 156340 260064 156392
rect 80980 156204 81032 156256
rect 178408 156272 178460 156324
rect 176200 156204 176252 156256
rect 121276 156136 121328 156188
rect 185308 156136 185360 156188
rect 87696 156068 87748 156120
rect 185400 156068 185452 156120
rect 185768 156272 185820 156324
rect 189816 156272 189868 156324
rect 195152 156272 195204 156324
rect 268108 156272 268160 156324
rect 185676 156204 185728 156256
rect 191288 156204 191340 156256
rect 192668 156204 192720 156256
rect 265164 156204 265216 156256
rect 255412 156136 255464 156188
rect 223212 156068 223264 156120
rect 94412 156000 94464 156052
rect 185676 156000 185728 156052
rect 77576 155932 77628 155984
rect 174544 155932 174596 155984
rect 175832 155932 175884 155984
rect 205180 155932 205232 155984
rect 15476 155864 15528 155916
rect 84200 155864 84252 155916
rect 84292 155864 84344 155916
rect 85396 155864 85448 155916
rect 95240 155864 95292 155916
rect 96528 155864 96580 155916
rect 101128 155864 101180 155916
rect 102048 155864 102100 155916
rect 106188 155864 106240 155916
rect 109408 155864 109460 155916
rect 109500 155864 109552 155916
rect 111616 155864 111668 155916
rect 111800 155864 111852 155916
rect 195704 155864 195756 155916
rect 12072 155660 12124 155712
rect 76748 155796 76800 155848
rect 66720 155728 66772 155780
rect 82820 155728 82872 155780
rect 77116 155660 77168 155712
rect 81808 155660 81860 155712
rect 82728 155660 82780 155712
rect 83464 155796 83516 155848
rect 173440 155796 173492 155848
rect 83004 155728 83056 155780
rect 152924 155728 152976 155780
rect 153660 155728 153712 155780
rect 156696 155728 156748 155780
rect 158812 155728 158864 155780
rect 175648 155796 175700 155848
rect 175832 155796 175884 155848
rect 177764 155796 177816 155848
rect 180064 155796 180116 155848
rect 185492 155796 185544 155848
rect 174176 155728 174228 155780
rect 49884 155592 49936 155644
rect 134616 155592 134668 155644
rect 134708 155592 134760 155644
rect 135168 155592 135220 155644
rect 136364 155592 136416 155644
rect 146944 155592 146996 155644
rect 164240 155660 164292 155712
rect 153292 155592 153344 155644
rect 167460 155660 167512 155712
rect 171048 155660 171100 155712
rect 171140 155660 171192 155712
rect 176016 155660 176068 155712
rect 177580 155728 177632 155780
rect 187516 155796 187568 155848
rect 187608 155796 187660 155848
rect 185676 155728 185728 155780
rect 191104 155728 191156 155780
rect 194324 155796 194376 155848
rect 200672 155864 200724 155916
rect 200764 155864 200816 155916
rect 205916 155864 205968 155916
rect 206928 155864 206980 155916
rect 209780 155932 209832 155984
rect 244556 155932 244608 155984
rect 246304 155932 246356 155984
rect 200304 155796 200356 155848
rect 201040 155796 201092 155848
rect 270224 155864 270276 155916
rect 270776 155864 270828 155916
rect 277216 155864 277268 155916
rect 283012 155932 283064 155984
rect 292212 155932 292264 155984
rect 295800 155932 295852 155984
rect 321376 155932 321428 155984
rect 321560 155932 321612 155984
rect 324504 155932 324556 155984
rect 326620 155932 326672 155984
rect 209688 155796 209740 155848
rect 200396 155728 200448 155780
rect 200580 155728 200632 155780
rect 240416 155728 240468 155780
rect 240508 155728 240560 155780
rect 196900 155660 196952 155712
rect 200212 155660 200264 155712
rect 200304 155660 200356 155712
rect 244556 155660 244608 155712
rect 222752 155592 222804 155644
rect 222844 155592 222896 155644
rect 223488 155592 223540 155644
rect 223580 155592 223632 155644
rect 228456 155592 228508 155644
rect 230388 155592 230440 155644
rect 233976 155592 234028 155644
rect 234620 155592 234672 155644
rect 243544 155592 243596 155644
rect 244832 155728 244884 155780
rect 248144 155728 248196 155780
rect 249064 155728 249116 155780
rect 257252 155728 257304 155780
rect 259828 155796 259880 155848
rect 281632 155864 281684 155916
rect 299434 155864 299486 155916
rect 299572 155864 299624 155916
rect 326160 155864 326212 155916
rect 333612 156000 333664 156052
rect 336004 156000 336056 156052
rect 277492 155796 277544 155848
rect 282460 155796 282512 155848
rect 283288 155796 283340 155848
rect 287336 155796 287388 155848
rect 287520 155796 287572 155848
rect 295708 155796 295760 155848
rect 295800 155796 295852 155848
rect 326436 155796 326488 155848
rect 335268 155864 335320 155916
rect 348884 155932 348936 155984
rect 356520 155932 356572 155984
rect 261392 155728 261444 155780
rect 261484 155728 261536 155780
rect 299480 155728 299532 155780
rect 299572 155728 299624 155780
rect 311624 155728 311676 155780
rect 246304 155660 246356 155712
rect 262128 155660 262180 155712
rect 264060 155660 264112 155712
rect 266728 155660 266780 155712
rect 268200 155660 268252 155712
rect 321376 155728 321428 155780
rect 321468 155728 321520 155780
rect 331772 155728 331824 155780
rect 312084 155660 312136 155712
rect 315948 155660 316000 155712
rect 316592 155660 316644 155712
rect 320180 155660 320232 155712
rect 320272 155660 320324 155712
rect 326344 155660 326396 155712
rect 326528 155660 326580 155712
rect 333796 155796 333848 155848
rect 336188 155796 336240 155848
rect 343916 155864 343968 155916
rect 344652 155864 344704 155916
rect 382372 155864 382424 155916
rect 337844 155796 337896 155848
rect 337936 155796 337988 155848
rect 340788 155796 340840 155848
rect 342168 155796 342220 155848
rect 380532 155796 380584 155848
rect 381636 155796 381688 155848
rect 398840 155796 398892 155848
rect 331956 155728 332008 155780
rect 351276 155728 351328 155780
rect 355232 155728 355284 155780
rect 357992 155728 358044 155780
rect 358084 155728 358136 155780
rect 364708 155728 364760 155780
rect 364800 155728 364852 155780
rect 384580 155728 384632 155780
rect 388352 155728 388404 155780
rect 402244 155864 402296 155916
rect 411812 155864 411864 155916
rect 413928 155864 413980 155916
rect 443736 155864 443788 155916
rect 458272 155864 458324 155916
rect 460572 155864 460624 155916
rect 470508 155864 470560 155916
rect 471428 155864 471480 155916
rect 476120 155864 476172 155916
rect 476488 155864 476540 155916
rect 482928 155864 482980 155916
rect 488264 155864 488316 155916
rect 490380 155864 490432 155916
rect 499212 155864 499264 155916
rect 500592 155864 500644 155916
rect 509056 155864 509108 155916
rect 510068 155864 510120 155916
rect 516048 155864 516100 155916
rect 519360 155864 519412 155916
rect 401784 155796 401836 155848
rect 407304 155796 407356 155848
rect 419356 155796 419408 155848
rect 423220 155796 423272 155848
rect 442080 155796 442132 155848
rect 456984 155796 457036 155848
rect 458916 155796 458968 155848
rect 399208 155728 399260 155780
rect 416688 155728 416740 155780
rect 424416 155728 424468 155780
rect 437480 155728 437532 155780
rect 439596 155728 439648 155780
rect 455052 155728 455104 155780
rect 456340 155728 456392 155780
rect 464344 155728 464396 155780
rect 332048 155660 332100 155712
rect 333980 155660 334032 155712
rect 335452 155660 335504 155712
rect 292580 155592 292632 155644
rect 295892 155592 295944 155644
rect 299664 155592 299716 155644
rect 300124 155592 300176 155644
rect 302792 155592 302844 155644
rect 302884 155592 302936 155644
rect 340972 155592 341024 155644
rect 341064 155592 341116 155644
rect 349896 155592 349948 155644
rect 365352 155660 365404 155712
rect 382464 155660 382516 155712
rect 356520 155592 356572 155644
rect 365076 155592 365128 155644
rect 365260 155592 365312 155644
rect 385592 155592 385644 155644
rect 398380 155592 398432 155644
rect 404912 155592 404964 155644
rect 405096 155660 405148 155712
rect 408868 155660 408920 155712
rect 433708 155660 433760 155712
rect 448612 155660 448664 155712
rect 411352 155592 411404 155644
rect 412640 155592 412692 155644
rect 420184 155592 420236 155644
rect 435364 155592 435416 155644
rect 60004 155524 60056 155576
rect 153660 155524 153712 155576
rect 154856 155524 154908 155576
rect 155684 155524 155736 155576
rect 156512 155524 156564 155576
rect 158812 155524 158864 155576
rect 159916 155524 159968 155576
rect 164332 155524 164384 155576
rect 164424 155524 164476 155576
rect 169760 155524 169812 155576
rect 170864 155524 170916 155576
rect 173256 155524 173308 155576
rect 173348 155524 173400 155576
rect 180064 155524 180116 155576
rect 180892 155524 180944 155576
rect 185676 155524 185728 155576
rect 70032 155456 70084 155508
rect 162124 155456 162176 155508
rect 164148 155456 164200 155508
rect 165620 155456 165672 155508
rect 166632 155456 166684 155508
rect 232320 155524 232372 155576
rect 232504 155524 232556 155576
rect 233148 155524 233200 155576
rect 233884 155524 233936 155576
rect 272524 155524 272576 155576
rect 272708 155524 272760 155576
rect 299572 155524 299624 155576
rect 306840 155524 306892 155576
rect 325424 155524 325476 155576
rect 326620 155524 326672 155576
rect 328644 155524 328696 155576
rect 328736 155524 328788 155576
rect 336096 155524 336148 155576
rect 336188 155524 336240 155576
rect 364984 155524 365036 155576
rect 365352 155524 365404 155576
rect 375472 155524 375524 155576
rect 379060 155524 379112 155576
rect 408776 155524 408828 155576
rect 410156 155524 410208 155576
rect 417424 155524 417476 155576
rect 421104 155524 421156 155576
rect 430580 155524 430632 155576
rect 431960 155524 432012 155576
rect 445208 155524 445260 155576
rect 446404 155592 446456 155644
rect 452844 155660 452896 155712
rect 453856 155660 453908 155712
rect 465540 155660 465592 155712
rect 466460 155796 466512 155848
rect 473084 155796 473136 155848
rect 480720 155796 480772 155848
rect 486332 155796 486384 155848
rect 498384 155796 498436 155848
rect 499580 155796 499632 155848
rect 469312 155728 469364 155780
rect 469772 155728 469824 155780
rect 474740 155728 474792 155780
rect 479064 155728 479116 155780
rect 484952 155728 485004 155780
rect 517336 155728 517388 155780
rect 521016 155728 521068 155780
rect 468116 155660 468168 155712
rect 473636 155660 473688 155712
rect 475660 155660 475712 155712
rect 480720 155660 480772 155712
rect 492496 155660 492548 155712
rect 495348 155660 495400 155712
rect 515496 155660 515548 155712
rect 518532 155660 518584 155712
rect 452108 155592 452160 155644
rect 186780 155456 186832 155508
rect 191012 155456 191064 155508
rect 191104 155456 191156 155508
rect 249064 155456 249116 155508
rect 249156 155456 249208 155508
rect 254124 155456 254176 155508
rect 257344 155456 257396 155508
rect 260564 155456 260616 155508
rect 260656 155456 260708 155508
rect 311716 155456 311768 155508
rect 311808 155456 311860 155508
rect 314568 155456 314620 155508
rect 315304 155456 315356 155508
rect 321376 155456 321428 155508
rect 321468 155456 321520 155508
rect 10416 155388 10468 155440
rect 107752 155388 107804 155440
rect 107844 155388 107896 155440
rect 108948 155388 109000 155440
rect 109040 155388 109092 155440
rect 110144 155388 110196 155440
rect 111156 155388 111208 155440
rect 111708 155388 111760 155440
rect 115388 155388 115440 155440
rect 115848 155388 115900 155440
rect 116216 155388 116268 155440
rect 117228 155388 117280 155440
rect 117872 155388 117924 155440
rect 118608 155388 118660 155440
rect 120540 155388 120592 155440
rect 122748 155388 122800 155440
rect 123484 155388 123536 155440
rect 200764 155388 200816 155440
rect 200856 155388 200908 155440
rect 209688 155388 209740 155440
rect 209780 155388 209832 155440
rect 262864 155388 262916 155440
rect 264888 155388 264940 155440
rect 266452 155388 266504 155440
rect 267372 155388 267424 155440
rect 272524 155388 272576 155440
rect 272800 155388 272852 155440
rect 273996 155388 274048 155440
rect 274088 155388 274140 155440
rect 299664 155388 299716 155440
rect 299756 155388 299808 155440
rect 316684 155388 316736 155440
rect 316776 155388 316828 155440
rect 320272 155388 320324 155440
rect 327264 155456 327316 155508
rect 351644 155456 351696 155508
rect 351736 155456 351788 155508
rect 355232 155456 355284 155508
rect 355324 155456 355376 155508
rect 362684 155456 362736 155508
rect 369032 155456 369084 155508
rect 401048 155456 401100 155508
rect 405924 155456 405976 155508
rect 419172 155456 419224 155508
rect 426992 155456 427044 155508
rect 445116 155456 445168 155508
rect 325240 155388 325292 155440
rect 325424 155388 325476 155440
rect 331220 155388 331272 155440
rect 331312 155388 331364 155440
rect 335912 155388 335964 155440
rect 336096 155388 336148 155440
rect 370228 155388 370280 155440
rect 375748 155388 375800 155440
rect 406200 155388 406252 155440
rect 413560 155388 413612 155440
rect 435088 155388 435140 155440
rect 438676 155388 438728 155440
rect 446404 155388 446456 155440
rect 449624 155524 449676 155576
rect 462688 155524 462740 155576
rect 463884 155592 463936 155644
rect 473360 155592 473412 155644
rect 474832 155592 474884 155644
rect 480812 155592 480864 155644
rect 481548 155592 481600 155644
rect 487068 155592 487120 155644
rect 491668 155592 491720 155644
rect 494612 155592 494664 155644
rect 513564 155592 513616 155644
rect 515956 155592 516008 155644
rect 464620 155524 464672 155576
rect 464712 155524 464764 155576
rect 473912 155524 473964 155576
rect 483204 155524 483256 155576
rect 485872 155524 485924 155576
rect 490748 155524 490800 155576
rect 493968 155524 494020 155576
rect 494152 155524 494204 155576
rect 496728 155524 496780 155576
rect 497464 155524 497516 155576
rect 499304 155524 499356 155576
rect 501696 155524 501748 155576
rect 502432 155524 502484 155576
rect 507768 155524 507820 155576
rect 508412 155524 508464 155576
rect 510528 155524 510580 155576
rect 511816 155524 511868 155576
rect 512276 155524 512328 155576
rect 514300 155524 514352 155576
rect 514852 155524 514904 155576
rect 517612 155524 517664 155576
rect 447968 155456 448020 155508
rect 461400 155456 461452 155508
rect 464344 155456 464396 155508
rect 467748 155456 467800 155508
rect 472348 155456 472400 155508
rect 477592 155456 477644 155508
rect 482376 155456 482428 155508
rect 487712 155456 487764 155508
rect 500040 155456 500092 155508
rect 501236 155456 501288 155508
rect 514208 155456 514260 155508
rect 516784 155456 516836 155508
rect 449992 155388 450044 155440
rect 450452 155388 450504 155440
rect 454592 155388 454644 155440
rect 454684 155388 454736 155440
rect 466368 155388 466420 155440
rect 468944 155388 468996 155440
rect 477500 155388 477552 155440
rect 478144 155388 478196 155440
rect 484308 155388 484360 155440
rect 11244 155320 11296 155372
rect 12348 155320 12400 155372
rect 36452 155320 36504 155372
rect 50344 155320 50396 155372
rect 53288 155320 53340 155372
rect 153936 155320 153988 155372
rect 154028 155320 154080 155372
rect 160652 155320 160704 155372
rect 160744 155320 160796 155372
rect 175924 155320 175976 155372
rect 176016 155320 176068 155372
rect 242900 155320 242952 155372
rect 242992 155320 243044 155372
rect 244648 155320 244700 155372
rect 244740 155320 244792 155372
rect 252560 155320 252612 155372
rect 253940 155320 253992 155372
rect 299572 155320 299624 155372
rect 299848 155320 299900 155372
rect 311900 155320 311952 155372
rect 311992 155320 312044 155372
rect 313188 155320 313240 155372
rect 314384 155320 314436 155372
rect 39856 155252 39908 155304
rect 132960 155252 133012 155304
rect 133052 155252 133104 155304
rect 137008 155252 137060 155304
rect 137376 155252 137428 155304
rect 140780 155252 140832 155304
rect 143080 155252 143132 155304
rect 17960 155184 18012 155236
rect 19248 155184 19300 155236
rect 22192 155184 22244 155236
rect 135904 155184 135956 155236
rect 137192 155184 137244 155236
rect 142620 155184 142672 155236
rect 143908 155184 143960 155236
rect 147588 155184 147640 155236
rect 149796 155184 149848 155236
rect 156604 155184 156656 155236
rect 191012 155252 191064 155304
rect 191104 155252 191156 155304
rect 230388 155252 230440 155304
rect 230480 155252 230532 155304
rect 238668 155252 238720 155304
rect 238760 155252 238812 155304
rect 245476 155252 245528 155304
rect 248052 155252 248104 155304
rect 294052 155252 294104 155304
rect 160836 155184 160888 155236
rect 234620 155184 234672 155236
rect 237196 155184 237248 155236
rect 240508 155184 240560 155236
rect 241336 155184 241388 155236
rect 299480 155252 299532 155304
rect 302792 155252 302844 155304
rect 307116 155252 307168 155304
rect 294236 155184 294288 155236
rect 300860 155184 300912 155236
rect 300952 155184 301004 155236
rect 302884 155184 302936 155236
rect 304356 155184 304408 155236
rect 306380 155184 306432 155236
rect 306932 155184 306984 155236
rect 308496 155252 308548 155304
rect 308588 155252 308640 155304
rect 341064 155252 341116 155304
rect 307668 155184 307720 155236
rect 348792 155252 348844 155304
rect 351276 155252 351328 155304
rect 355416 155252 355468 155304
rect 362316 155320 362368 155372
rect 394884 155320 394936 155372
rect 406844 155320 406896 155372
rect 422668 155320 422720 155372
rect 422760 155320 422812 155372
rect 424968 155320 425020 155372
rect 437020 155320 437072 155372
rect 451280 155320 451332 155372
rect 358452 155252 358504 155304
rect 364708 155252 364760 155304
rect 392400 155252 392452 155304
rect 395068 155252 395120 155304
rect 405648 155252 405700 155304
rect 420276 155252 420328 155304
rect 440240 155252 440292 155304
rect 442908 155252 442960 155304
rect 453120 155320 453172 155372
rect 465080 155320 465132 155372
rect 465632 155320 465684 155372
rect 474924 155320 474976 155372
rect 489920 155320 489972 155372
rect 493232 155320 493284 155372
rect 495808 155320 495860 155372
rect 496912 155320 496964 155372
rect 518072 155320 518124 155372
rect 521844 155320 521896 155372
rect 456800 155252 456852 155304
rect 462228 155252 462280 155304
rect 472348 155252 472400 155304
rect 473176 155252 473228 155304
rect 477684 155252 477736 155304
rect 479892 155252 479944 155304
rect 485688 155252 485740 155304
rect 487436 155252 487488 155304
rect 491208 155252 491260 155304
rect 494980 155252 495032 155304
rect 497372 155252 497424 155304
rect 512920 155252 512972 155304
rect 515128 155252 515180 155304
rect 518808 155252 518860 155304
rect 522672 155252 522724 155304
rect 341248 155184 341300 155236
rect 344928 155184 344980 155236
rect 355600 155184 355652 155236
rect 390744 155184 390796 155236
rect 404268 155184 404320 155236
rect 427728 155184 427780 155236
rect 434536 155184 434588 155236
rect 448520 155184 448572 155236
rect 454592 155184 454644 155236
rect 462320 155184 462372 155236
rect 467288 155184 467340 155236
rect 476212 155184 476264 155236
rect 493324 155184 493376 155236
rect 495808 155184 495860 155236
rect 503352 155184 503404 155236
rect 503812 155184 503864 155236
rect 510988 155184 511040 155236
rect 512644 155184 512696 155236
rect 516784 155184 516836 155236
rect 520188 155184 520240 155236
rect 521844 155184 521896 155236
rect 523500 155184 523552 155236
rect 90180 155116 90232 155168
rect 175832 155116 175884 155168
rect 175924 155116 175976 155168
rect 191104 155116 191156 155168
rect 191196 155116 191248 155168
rect 249156 155116 249208 155168
rect 253112 155116 253164 155168
rect 272616 155116 272668 155168
rect 273260 155116 273312 155168
rect 282092 155116 282144 155168
rect 282184 155116 282236 155168
rect 283288 155116 283340 155168
rect 283380 155116 283432 155168
rect 284300 155116 284352 155168
rect 286692 155116 286744 155168
rect 292304 155116 292356 155168
rect 292580 155116 292632 155168
rect 295616 155116 295668 155168
rect 295708 155116 295760 155168
rect 326436 155116 326488 155168
rect 326988 155116 327040 155168
rect 351276 155116 351328 155168
rect 351828 155116 351880 155168
rect 387616 155116 387668 155168
rect 391664 155116 391716 155168
rect 404176 155116 404228 155168
rect 416044 155116 416096 155168
rect 422576 155116 422628 155168
rect 422668 155116 422720 155168
rect 429936 155116 429988 155168
rect 437848 155116 437900 155168
rect 453212 155116 453264 155168
rect 457996 155116 458048 155168
rect 468024 155116 468076 155168
rect 484860 155116 484912 155168
rect 488448 155116 488500 155168
rect 489092 155116 489144 155168
rect 492588 155116 492640 155168
rect 84200 155048 84252 155100
rect 91100 155048 91152 155100
rect 96896 155048 96948 155100
rect 184204 155048 184256 155100
rect 184296 155048 184348 155100
rect 186136 155048 186188 155100
rect 187516 155048 187568 155100
rect 190828 155048 190880 155100
rect 191012 155048 191064 155100
rect 200488 155048 200540 155100
rect 200764 155048 200816 155100
rect 260196 155048 260248 155100
rect 261392 155048 261444 155100
rect 262772 155048 262824 155100
rect 262864 155048 262916 155100
rect 269028 155048 269080 155100
rect 269948 155048 270000 155100
rect 299388 155048 299440 155100
rect 300860 155048 300912 155100
rect 336004 155048 336056 155100
rect 336096 155048 336148 155100
rect 341156 155048 341208 155100
rect 341340 155048 341392 155100
rect 342076 155048 342128 155100
rect 343824 155048 343876 155100
rect 377220 155048 377272 155100
rect 380808 155048 380860 155100
rect 384488 155048 384540 155100
rect 384580 155048 384632 155100
rect 395436 155048 395488 155100
rect 408500 155048 408552 155100
rect 411720 155048 411772 155100
rect 436192 155048 436244 155100
rect 451372 155048 451424 155100
rect 451464 155048 451516 155100
rect 463700 155048 463752 155100
rect 470692 155048 470744 155100
rect 477408 155048 477460 155100
rect 64144 154980 64196 155032
rect 57428 154912 57480 154964
rect 103520 154912 103572 154964
rect 103612 154912 103664 154964
rect 111800 154912 111852 154964
rect 114560 154980 114612 155032
rect 115756 154980 115808 155032
rect 115940 154980 115992 155032
rect 117136 154980 117188 155032
rect 117228 154980 117280 155032
rect 120632 154980 120684 155032
rect 123392 154980 123444 155032
rect 123760 154980 123812 155032
rect 128268 154980 128320 155032
rect 130476 154980 130528 155032
rect 133236 154980 133288 155032
rect 133880 154980 133932 155032
rect 79324 154844 79376 154896
rect 113180 154844 113232 154896
rect 86040 154776 86092 154828
rect 116584 154844 116636 154896
rect 117044 154844 117096 154896
rect 128544 154912 128596 154964
rect 134616 154912 134668 154964
rect 136916 154912 136968 154964
rect 137652 154980 137704 155032
rect 213092 154980 213144 155032
rect 213644 154980 213696 155032
rect 216496 154980 216548 155032
rect 221188 154980 221240 155032
rect 279884 154980 279936 155032
rect 279976 154980 280028 155032
rect 287704 154980 287756 155032
rect 288348 154980 288400 155032
rect 321928 154980 321980 155032
rect 322112 154980 322164 155032
rect 325976 154980 326028 155032
rect 326344 154980 326396 155032
rect 211896 154912 211948 154964
rect 211988 154912 212040 154964
rect 212448 154912 212500 154964
rect 212540 154912 212592 154964
rect 214380 154912 214432 154964
rect 214564 154912 214616 154964
rect 232044 154912 232096 154964
rect 232320 154912 232372 154964
rect 241428 154912 241480 154964
rect 243544 154912 243596 154964
rect 292396 154912 292448 154964
rect 294052 154912 294104 154964
rect 306932 154912 306984 154964
rect 307208 154912 307260 154964
rect 321836 154912 321888 154964
rect 322204 154912 322256 154964
rect 340512 154912 340564 154964
rect 355232 154980 355284 155032
rect 355416 154980 355468 155032
rect 357440 154980 357492 155032
rect 371516 154980 371568 155032
rect 341064 154912 341116 154964
rect 348792 154912 348844 154964
rect 127164 154844 127216 154896
rect 137376 154844 137428 154896
rect 137560 154844 137612 154896
rect 144828 154844 144880 154896
rect 146944 154844 146996 154896
rect 155868 154844 155920 154896
rect 113456 154776 113508 154828
rect 120540 154776 120592 154828
rect 120632 154776 120684 154828
rect 153016 154776 153068 154828
rect 153108 154776 153160 154828
rect 161204 154844 161256 154896
rect 161296 154844 161348 154896
rect 164240 154844 164292 154896
rect 164332 154844 164384 154896
rect 233700 154844 233752 154896
rect 233792 154844 233844 154896
rect 156604 154776 156656 154828
rect 103520 154708 103572 154760
rect 109132 154708 109184 154760
rect 109408 154708 109460 154760
rect 161296 154708 161348 154760
rect 220728 154776 220780 154828
rect 223764 154776 223816 154828
rect 226984 154776 227036 154828
rect 227076 154776 227128 154828
rect 233884 154776 233936 154828
rect 233976 154776 234028 154828
rect 237380 154776 237432 154828
rect 238024 154844 238076 154896
rect 238760 154844 238812 154896
rect 238852 154844 238904 154896
rect 247132 154844 247184 154896
rect 247224 154844 247276 154896
rect 238576 154776 238628 154828
rect 238668 154776 238720 154828
rect 162124 154708 162176 154760
rect 167644 154708 167696 154760
rect 175832 154708 175884 154760
rect 183284 154708 183336 154760
rect 184204 154708 184256 154760
rect 99472 154640 99524 154692
rect 116768 154640 116820 154692
rect 116860 154640 116912 154692
rect 121276 154640 121328 154692
rect 122932 154640 122984 154692
rect 92756 154572 92808 154624
rect 113640 154572 113692 154624
rect 113732 154572 113784 154624
rect 123484 154572 123536 154624
rect 128820 154640 128872 154692
rect 129556 154640 129608 154692
rect 129648 154640 129700 154692
rect 184940 154640 184992 154692
rect 184848 154572 184900 154624
rect 185492 154708 185544 154760
rect 238760 154708 238812 154760
rect 239036 154776 239088 154828
rect 282184 154776 282236 154828
rect 285036 154776 285088 154828
rect 287060 154776 287112 154828
rect 287520 154776 287572 154828
rect 291200 154776 291252 154828
rect 292120 154776 292172 154828
rect 293132 154776 293184 154828
rect 293408 154844 293460 154896
rect 321376 154844 321428 154896
rect 321928 154844 321980 154896
rect 326528 154844 326580 154896
rect 326620 154844 326672 154896
rect 355324 154912 355376 154964
rect 357256 154912 357308 154964
rect 380992 154912 381044 154964
rect 396448 154980 396500 155032
rect 441252 154980 441304 155032
rect 455420 154980 455472 155032
rect 455512 154980 455564 155032
rect 384672 154912 384724 154964
rect 388536 154912 388588 154964
rect 392492 154912 392544 154964
rect 415492 154912 415544 154964
rect 440424 154912 440476 154964
rect 455696 154912 455748 154964
rect 457168 154980 457220 155032
rect 468484 154980 468536 155032
rect 474004 154980 474056 155032
rect 479524 154980 479576 155032
rect 511632 154980 511684 155032
rect 513472 154980 513524 155032
rect 467012 154912 467064 154964
rect 351644 154844 351696 154896
rect 364248 154844 364300 154896
rect 364984 154844 365036 154896
rect 374000 154844 374052 154896
rect 374920 154844 374972 154896
rect 398104 154844 398156 154896
rect 446312 154844 446364 154896
rect 459652 154844 459704 154896
rect 294328 154776 294380 154828
rect 281448 154708 281500 154760
rect 282092 154708 282144 154760
rect 306932 154776 306984 154828
rect 310244 154776 310296 154828
rect 340328 154776 340380 154828
rect 294696 154708 294748 154760
rect 301044 154708 301096 154760
rect 301872 154708 301924 154760
rect 307024 154708 307076 154760
rect 307116 154708 307168 154760
rect 185124 154640 185176 154692
rect 193220 154640 193272 154692
rect 193496 154640 193548 154692
rect 200764 154640 200816 154692
rect 200948 154640 201000 154692
rect 209596 154640 209648 154692
rect 209688 154640 209740 154692
rect 263600 154640 263652 154692
rect 263692 154640 263744 154692
rect 264520 154640 264572 154692
rect 266544 154640 266596 154692
rect 188988 154572 189040 154624
rect 190920 154572 190972 154624
rect 191840 154572 191892 154624
rect 192024 154572 192076 154624
rect 194600 154572 194652 154624
rect 197728 154572 197780 154624
rect 214564 154572 214616 154624
rect 216496 154572 216548 154624
rect 271512 154572 271564 154624
rect 272616 154640 272668 154692
rect 278688 154640 278740 154692
rect 280804 154640 280856 154692
rect 287520 154572 287572 154624
rect 287704 154640 287756 154692
rect 311440 154640 311492 154692
rect 311808 154708 311860 154760
rect 313464 154708 313516 154760
rect 313556 154708 313608 154760
rect 340236 154708 340288 154760
rect 292212 154572 292264 154624
rect 292488 154572 292540 154624
rect 316592 154572 316644 154624
rect 316684 154572 316736 154624
rect 321836 154572 321888 154624
rect 322020 154640 322072 154692
rect 326620 154640 326672 154692
rect 327908 154640 327960 154692
rect 363880 154776 363932 154828
rect 363972 154776 364024 154828
rect 386236 154776 386288 154828
rect 444564 154776 444616 154828
rect 458364 154776 458416 154828
rect 463056 154776 463108 154828
rect 471980 154776 472032 154828
rect 484032 154776 484084 154828
rect 489000 154776 489052 154828
rect 509700 154776 509752 154828
rect 510896 154776 510948 154828
rect 340880 154708 340932 154760
rect 351828 154708 351880 154760
rect 353852 154708 353904 154760
rect 380900 154708 380952 154760
rect 341156 154640 341208 154692
rect 367100 154640 367152 154692
rect 367376 154640 367428 154692
rect 385684 154708 385736 154760
rect 385776 154708 385828 154760
rect 413192 154708 413244 154760
rect 445392 154708 445444 154760
rect 458732 154708 458784 154760
rect 461492 154708 461544 154760
rect 471704 154708 471756 154760
rect 485780 154708 485832 154760
rect 488908 154708 488960 154760
rect 496636 154708 496688 154760
rect 498200 154708 498252 154760
rect 387524 154640 387576 154692
rect 390928 154640 390980 154692
rect 445208 154640 445260 154692
rect 447232 154640 447284 154692
rect 448796 154640 448848 154692
rect 459560 154640 459612 154692
rect 477316 154640 477368 154692
rect 481732 154640 481784 154692
rect 326068 154572 326120 154624
rect 326160 154572 326212 154624
rect 332508 154572 332560 154624
rect 334624 154572 334676 154624
rect 368480 154572 368532 154624
rect 374092 154572 374144 154624
rect 388444 154572 388496 154624
rect 390836 154572 390888 154624
rect 392308 154572 392360 154624
rect 447140 154572 447192 154624
rect 458180 154572 458232 154624
rect 459744 154572 459796 154624
rect 470416 154572 470468 154624
rect 486608 154572 486660 154624
rect 488540 154572 488592 154624
rect 51540 154504 51592 154556
rect 158352 154504 158404 154556
rect 159088 154504 159140 154556
rect 238024 154504 238076 154556
rect 54944 154436 54996 154488
rect 160928 154436 160980 154488
rect 162032 154436 162084 154488
rect 243084 154504 243136 154556
rect 245568 154504 245620 154556
rect 248788 154504 248840 154556
rect 248880 154504 248932 154556
rect 238944 154436 238996 154488
rect 249064 154436 249116 154488
rect 249156 154436 249208 154488
rect 48228 154368 48280 154420
rect 155592 154368 155644 154420
rect 155776 154368 155828 154420
rect 41512 154300 41564 154352
rect 150624 154300 150676 154352
rect 152372 154300 152424 154352
rect 34796 154232 34848 154284
rect 145564 154232 145616 154284
rect 145656 154232 145708 154284
rect 230296 154232 230348 154284
rect 232964 154300 233016 154352
rect 235264 154368 235316 154420
rect 235356 154368 235408 154420
rect 238116 154368 238168 154420
rect 238208 154368 238260 154420
rect 240600 154368 240652 154420
rect 242164 154368 242216 154420
rect 299480 154436 299532 154488
rect 306932 154504 306984 154556
rect 316408 154504 316460 154556
rect 316500 154504 316552 154556
rect 360660 154504 360712 154556
rect 363880 154504 363932 154556
rect 369584 154504 369636 154556
rect 369860 154504 369912 154556
rect 401692 154504 401744 154556
rect 233700 154300 233752 154352
rect 236184 154300 236236 154352
rect 236368 154300 236420 154352
rect 292672 154300 292724 154352
rect 306656 154368 306708 154420
rect 306932 154368 306984 154420
rect 307116 154436 307168 154488
rect 311440 154436 311492 154488
rect 312728 154436 312780 154488
rect 358084 154436 358136 154488
rect 363144 154436 363196 154488
rect 396540 154436 396592 154488
rect 403440 154436 403492 154488
rect 427360 154436 427412 154488
rect 309232 154368 309284 154420
rect 309416 154368 309468 154420
rect 355508 154368 355560 154420
rect 358452 154368 358504 154420
rect 359372 154368 359424 154420
rect 366456 154368 366508 154420
rect 399116 154368 399168 154420
rect 400956 154368 401008 154420
rect 425520 154368 425572 154420
rect 304080 154300 304132 154352
rect 306012 154300 306064 154352
rect 352840 154300 352892 154352
rect 233148 154232 233200 154284
rect 292304 154232 292356 154284
rect 295984 154232 296036 154284
rect 336096 154232 336148 154284
rect 336188 154232 336240 154284
rect 340144 154232 340196 154284
rect 340420 154232 340472 154284
rect 345664 154232 345716 154284
rect 345756 154232 345808 154284
rect 350356 154232 350408 154284
rect 38108 154164 38160 154216
rect 148140 154164 148192 154216
rect 148968 154164 149020 154216
rect 232872 154164 232924 154216
rect 232964 154164 233016 154216
rect 235356 154164 235408 154216
rect 235448 154164 235500 154216
rect 287152 154164 287204 154216
rect 287796 154164 287848 154216
rect 292488 154164 292540 154216
rect 292948 154164 293000 154216
rect 30564 154096 30616 154148
rect 142344 154096 142396 154148
rect 142436 154096 142488 154148
rect 227720 154096 227772 154148
rect 228732 154096 228784 154148
rect 287612 154096 287664 154148
rect 291200 154096 291252 154148
rect 297364 154096 297416 154148
rect 13820 154028 13872 154080
rect 129464 154028 129516 154080
rect 129556 154028 129608 154080
rect 217416 154028 217468 154080
rect 217508 154028 217560 154080
rect 221924 154028 221976 154080
rect 222016 154028 222068 154080
rect 225328 154028 225380 154080
rect 225420 154028 225472 154080
rect 286968 154028 287020 154080
rect 287152 154028 287204 154080
rect 292396 154028 292448 154080
rect 292672 154028 292724 154080
rect 296444 154028 296496 154080
rect 297272 154028 297324 154080
rect 301596 154096 301648 154148
rect 302700 154164 302752 154216
rect 342720 154164 342772 154216
rect 342812 154164 342864 154216
rect 348516 154164 348568 154216
rect 351828 154164 351880 154216
rect 358728 154300 358780 154352
rect 359740 154300 359792 154352
rect 394056 154300 394108 154352
rect 400128 154300 400180 154352
rect 424876 154300 424928 154352
rect 355324 154232 355376 154284
rect 365720 154232 365772 154284
rect 393412 154232 393464 154284
rect 419724 154232 419776 154284
rect 353116 154164 353168 154216
rect 388904 154164 388956 154216
rect 396724 154164 396776 154216
rect 422300 154164 422352 154216
rect 336004 154096 336056 154148
rect 336096 154096 336148 154148
rect 345204 154096 345256 154148
rect 346308 154096 346360 154148
rect 383752 154096 383804 154148
rect 386604 154096 386656 154148
rect 414572 154096 414624 154148
rect 417424 154096 417476 154148
rect 432512 154096 432564 154148
rect 299296 154028 299348 154080
rect 347780 154028 347832 154080
rect 349712 154028 349764 154080
rect 386328 154028 386380 154080
rect 390008 154028 390060 154080
rect 417148 154028 417200 154080
rect 427820 154028 427872 154080
rect 446036 154028 446088 154080
rect 17132 153960 17184 154012
rect 132040 153960 132092 154012
rect 132224 153960 132276 154012
rect 219992 153960 220044 154012
rect 220728 153960 220780 154012
rect 228272 153960 228324 154012
rect 228364 153960 228416 154012
rect 288716 153960 288768 154012
rect 289268 153960 289320 154012
rect 335912 153960 335964 154012
rect 336004 153960 336056 154012
rect 342628 153960 342680 154012
rect 342996 153960 343048 154012
rect 381176 153960 381228 154012
rect 383292 153960 383344 154012
rect 411996 153960 412048 154012
rect 423588 153960 423640 154012
rect 442816 153960 442868 154012
rect 4528 153892 4580 153944
rect 122380 153892 122432 153944
rect 1216 153824 1268 153876
rect 119804 153824 119856 153876
rect 122104 153824 122156 153876
rect 212264 153892 212316 153944
rect 212816 153892 212868 153944
rect 217508 153892 217560 153944
rect 217600 153892 217652 153944
rect 280988 153892 281040 153944
rect 282552 153892 282604 153944
rect 125508 153824 125560 153876
rect 214840 153824 214892 153876
rect 215300 153824 215352 153876
rect 217692 153824 217744 153876
rect 218704 153824 218756 153876
rect 286140 153824 286192 153876
rect 286232 153824 286284 153876
rect 326068 153824 326120 153876
rect 58256 153756 58308 153808
rect 163504 153756 163556 153808
rect 165804 153756 165856 153808
rect 245660 153756 245712 153808
rect 68376 153688 68428 153740
rect 171232 153688 171284 153740
rect 175740 153688 175792 153740
rect 64972 153620 65024 153672
rect 168656 153620 168708 153672
rect 169116 153620 169168 153672
rect 248236 153688 248288 153740
rect 252284 153756 252336 153808
rect 306932 153756 306984 153808
rect 307024 153756 307076 153808
rect 325332 153756 325384 153808
rect 326252 153892 326304 153944
rect 326436 153824 326488 153876
rect 335544 153824 335596 153876
rect 336280 153892 336332 153944
rect 376024 153892 376076 153944
rect 376576 153892 376628 153944
rect 406844 153892 406896 153944
rect 407672 153892 407724 153944
rect 430488 153892 430540 153944
rect 430580 153892 430632 153944
rect 440884 153892 440936 153944
rect 337476 153824 337528 153876
rect 339592 153824 339644 153876
rect 378600 153824 378652 153876
rect 379888 153824 379940 153876
rect 409420 153824 409472 153876
rect 416872 153824 416924 153876
rect 437664 153824 437716 153876
rect 326528 153756 326580 153808
rect 326620 153756 326672 153808
rect 350724 153756 350776 153808
rect 253388 153688 253440 153740
rect 255596 153688 255648 153740
rect 311716 153688 311768 153740
rect 311808 153688 311860 153740
rect 312360 153688 312412 153740
rect 312728 153688 312780 153740
rect 324688 153688 324740 153740
rect 326344 153688 326396 153740
rect 363236 153756 363288 153808
rect 367100 153756 367152 153808
rect 372160 153756 372212 153808
rect 373172 153756 373224 153808
rect 404268 153756 404320 153808
rect 350908 153688 350960 153740
rect 355324 153688 355376 153740
rect 357440 153688 357492 153740
rect 368940 153688 368992 153740
rect 247132 153620 247184 153672
rect 256516 153620 256568 153672
rect 259000 153620 259052 153672
rect 316316 153620 316368 153672
rect 316408 153620 316460 153672
rect 327908 153620 327960 153672
rect 329564 153620 329616 153672
rect 370872 153620 370924 153672
rect 8760 153552 8812 153604
rect 109040 153552 109092 153604
rect 112076 153552 112128 153604
rect 204628 153552 204680 153604
rect 208584 153552 208636 153604
rect 278412 153552 278464 153604
rect 279148 153552 279200 153604
rect 75092 153484 75144 153536
rect 176384 153484 176436 153536
rect 182548 153484 182600 153536
rect 258540 153484 258592 153536
rect 269120 153484 269172 153536
rect 312360 153484 312412 153536
rect 332416 153552 332468 153604
rect 332876 153552 332928 153604
rect 373448 153552 373500 153604
rect 27252 153416 27304 153468
rect 125692 153416 125744 153468
rect 135536 153416 135588 153468
rect 222568 153416 222620 153468
rect 225328 153416 225380 153468
rect 228364 153416 228416 153468
rect 228456 153416 228508 153468
rect 236092 153416 236144 153468
rect 236184 153416 236236 153468
rect 241244 153416 241296 153468
rect 241428 153416 241480 153468
rect 246304 153416 246356 153468
rect 249064 153416 249116 153468
rect 297272 153416 297324 153468
rect 297364 153416 297416 153468
rect 322756 153484 322808 153536
rect 322848 153484 322900 153536
rect 326620 153484 326672 153536
rect 85120 153348 85172 153400
rect 184020 153348 184072 153400
rect 184848 153348 184900 153400
rect 88524 153280 88576 153332
rect 186596 153280 186648 153332
rect 189264 153348 189316 153400
rect 263692 153348 263744 153400
rect 272432 153348 272484 153400
rect 327264 153416 327316 153468
rect 312912 153348 312964 153400
rect 317604 153348 317656 153400
rect 317788 153348 317840 153400
rect 319352 153348 319404 153400
rect 319444 153348 319496 153400
rect 326344 153348 326396 153400
rect 326712 153348 326764 153400
rect 364892 153484 364944 153536
rect 327632 153416 327684 153468
rect 327540 153348 327592 153400
rect 331404 153348 331456 153400
rect 212908 153280 212960 153332
rect 213000 153280 213052 153332
rect 217600 153280 217652 153332
rect 217692 153280 217744 153332
rect 105360 153212 105412 153264
rect 199476 153212 199528 153264
rect 200488 153212 200540 153264
rect 220728 153212 220780 153264
rect 221924 153280 221976 153332
rect 281632 153280 281684 153332
rect 283012 153280 283064 153332
rect 286876 153280 286928 153332
rect 286968 153280 287020 153332
rect 291292 153280 291344 153332
rect 283564 153212 283616 153264
rect 284300 153212 284352 153264
rect 326436 153280 326488 153332
rect 326528 153280 326580 153332
rect 334900 153348 334952 153400
rect 335268 153348 335320 153400
rect 337016 153348 337068 153400
rect 337108 153348 337160 153400
rect 342904 153348 342956 153400
rect 331588 153280 331640 153332
rect 343272 153280 343324 153332
rect 345664 153416 345716 153468
rect 364984 153416 365036 153468
rect 345388 153348 345440 153400
rect 376668 153484 376720 153536
rect 365168 153416 365220 153468
rect 379244 153416 379296 153468
rect 368480 153348 368532 153400
rect 374736 153348 374788 153400
rect 348424 153280 348476 153332
rect 348516 153280 348568 153332
rect 356152 153280 356204 153332
rect 291476 153212 291528 153264
rect 311808 153212 311860 153264
rect 311900 153212 311952 153264
rect 314384 153212 314436 153264
rect 314568 153212 314620 153264
rect 316224 153212 316276 153264
rect 316316 153212 316368 153264
rect 316960 153212 317012 153264
rect 317144 153212 317196 153264
rect 333060 153212 333112 153264
rect 335912 153212 335964 153264
rect 340052 153212 340104 153264
rect 340144 153212 340196 153264
rect 353576 153212 353628 153264
rect 355232 153212 355284 153264
rect 363880 153280 363932 153332
rect 364892 153280 364944 153332
rect 368296 153280 368348 153332
rect 356428 153212 356480 153264
rect 391480 153212 391532 153264
rect 437480 153212 437532 153264
rect 443460 153212 443512 153264
rect 80152 153144 80204 153196
rect 180248 153144 180300 153196
rect 183284 153144 183336 153196
rect 187884 153144 187936 153196
rect 190092 153144 190144 153196
rect 264428 153144 264480 153196
rect 264520 153144 264572 153196
rect 315672 153144 315724 153196
rect 315948 153144 316000 153196
rect 318248 153144 318300 153196
rect 318616 153144 318668 153196
rect 362592 153144 362644 153196
rect 365628 153144 365680 153196
rect 398472 153144 398524 153196
rect 404176 153144 404228 153196
rect 418436 153144 418488 153196
rect 418528 153144 418580 153196
rect 438952 153144 439004 153196
rect 448520 153144 448572 153196
rect 451188 153144 451240 153196
rect 451280 153144 451332 153196
rect 453120 153144 453172 153196
rect 458180 153144 458232 153196
rect 460756 153144 460808 153196
rect 473084 153144 473136 153196
rect 475568 153144 475620 153196
rect 477408 153144 477460 153196
rect 478788 153144 478840 153196
rect 480812 153144 480864 153196
rect 482008 153144 482060 153196
rect 490380 153144 490432 153196
rect 492220 153144 492272 153196
rect 73436 153076 73488 153128
rect 175096 153076 175148 153128
rect 176660 153076 176712 153128
rect 63316 153008 63368 153060
rect 167368 153008 167420 153060
rect 169760 153008 169812 153060
rect 177672 153008 177724 153060
rect 177764 153008 177816 153060
rect 182732 153008 182784 153060
rect 186136 153076 186188 153128
rect 259828 153076 259880 153128
rect 260196 153076 260248 153128
rect 266912 153076 266964 153128
rect 271880 153076 271932 153128
rect 254032 153008 254084 153060
rect 254124 153008 254176 153060
rect 261760 153008 261812 153060
rect 263600 153008 263652 153060
rect 272064 153008 272116 153060
rect 276664 153076 276716 153128
rect 330484 153076 330536 153128
rect 330760 153076 330812 153128
rect 371516 153076 371568 153128
rect 377404 153076 377456 153128
rect 407488 153076 407540 153128
rect 414388 153076 414440 153128
rect 435732 153076 435784 153128
rect 447232 153076 447284 153128
rect 449256 153076 449308 153128
rect 452844 153076 452896 153128
rect 454408 153076 454460 153128
rect 473636 153076 473688 153128
rect 476948 153076 477000 153128
rect 481732 153076 481784 153128
rect 483940 153076 483992 153128
rect 326620 153008 326672 153060
rect 56600 152940 56652 152992
rect 162216 152940 162268 152992
rect 169944 152940 169996 152992
rect 248880 152940 248932 152992
rect 250628 152940 250680 152992
rect 254308 152940 254360 152992
rect 266728 152940 266780 152992
rect 320824 152940 320876 152992
rect 321560 152940 321612 152992
rect 324044 152940 324096 152992
rect 325700 152940 325752 152992
rect 367652 153008 367704 153060
rect 370688 153008 370740 153060
rect 402336 153008 402388 153060
rect 413928 153008 413980 153060
rect 433800 153008 433852 153060
rect 448612 153008 448664 153060
rect 450636 153008 450688 153060
rect 474740 153008 474792 153060
rect 478144 153008 478196 153060
rect 480720 153008 480772 153060
rect 482652 153008 482704 153060
rect 326804 152940 326856 152992
rect 366364 152940 366416 152992
rect 372344 152940 372396 152992
rect 403624 152940 403676 152992
rect 410984 152940 411036 152992
rect 433156 152940 433208 152992
rect 46572 152872 46624 152924
rect 154488 152872 154540 152924
rect 156696 152872 156748 152924
rect 164792 152872 164844 152924
rect 165620 152872 165672 152924
rect 244372 152872 244424 152924
rect 245476 152872 245528 152924
rect 300952 152872 301004 152924
rect 301044 152872 301096 152924
rect 307944 152872 307996 152924
rect 309140 152872 309192 152924
rect 313096 152872 313148 152924
rect 313188 152872 313240 152924
rect 313832 152872 313884 152924
rect 316684 152872 316736 152924
rect 351644 152872 351696 152924
rect 354772 152872 354824 152924
rect 390192 152872 390244 152924
rect 394240 152872 394292 152924
rect 420368 152872 420420 152924
rect 421932 152872 421984 152924
rect 441528 152872 441580 152924
rect 502524 152872 502576 152924
rect 503168 152872 503220 152924
rect 43168 152804 43220 152856
rect 151912 152804 151964 152856
rect 153936 152804 153988 152856
rect 159640 152804 159692 152856
rect 163228 152804 163280 152856
rect 243728 152804 243780 152856
rect 251456 152804 251508 152856
rect 33140 152736 33192 152788
rect 144276 152736 144328 152788
rect 144828 152736 144880 152788
rect 157064 152736 157116 152788
rect 157340 152736 157392 152788
rect 239312 152736 239364 152788
rect 242900 152736 242952 152788
rect 246948 152736 247000 152788
rect 258172 152804 258224 152856
rect 316316 152804 316368 152856
rect 317052 152804 317104 152856
rect 361304 152804 361356 152856
rect 368204 152804 368256 152856
rect 400404 152804 400456 152856
rect 409328 152804 409380 152856
rect 430580 152804 430632 152856
rect 431132 152804 431184 152856
rect 448612 152804 448664 152856
rect 488448 152804 488500 152856
rect 489644 152804 489696 152856
rect 311164 152736 311216 152788
rect 311532 152736 311584 152788
rect 356796 152736 356848 152788
rect 356888 152736 356940 152788
rect 26332 152668 26384 152720
rect 139124 152668 139176 152720
rect 139768 152668 139820 152720
rect 141792 152668 141844 152720
rect 147588 152668 147640 152720
rect 229008 152668 229060 152720
rect 233240 152668 233292 152720
rect 233976 152668 234028 152720
rect 234620 152668 234672 152720
rect 236736 152668 236788 152720
rect 240508 152668 240560 152720
rect 300308 152668 300360 152720
rect 32220 152600 32272 152652
rect 143632 152600 143684 152652
rect 146484 152600 146536 152652
rect 25504 152532 25556 152584
rect 138480 152532 138532 152584
rect 140780 152532 140832 152584
rect 149428 152532 149480 152584
rect 150716 152600 150768 152652
rect 234160 152600 234212 152652
rect 244280 152600 244332 152652
rect 230940 152532 230992 152584
rect 237380 152532 237432 152584
rect 241888 152532 241940 152584
rect 243544 152532 243596 152584
rect 249524 152532 249576 152584
rect 254308 152600 254360 152652
rect 310520 152668 310572 152720
rect 305000 152600 305052 152652
rect 351000 152668 351052 152720
rect 352196 152668 352248 152720
rect 360752 152736 360804 152788
rect 394700 152736 394752 152788
rect 397552 152736 397604 152788
rect 422944 152736 422996 152788
rect 424968 152736 425020 152788
rect 442172 152736 442224 152788
rect 476120 152736 476172 152788
rect 479432 152736 479484 152788
rect 302516 152532 302568 152584
rect 12900 152464 12952 152516
rect 128820 152464 128872 152516
rect 137008 152464 137060 152516
rect 137284 152464 137336 152516
rect 138020 152464 138072 152516
rect 141700 152464 141752 152516
rect 141792 152464 141844 152516
rect 225788 152464 225840 152516
rect 231308 152464 231360 152516
rect 295800 152464 295852 152516
rect 299572 152464 299624 152516
rect 302884 152464 302936 152516
rect 303436 152532 303488 152584
rect 313464 152600 313516 152652
rect 318892 152600 318944 152652
rect 318984 152600 319036 152652
rect 357440 152600 357492 152652
rect 305184 152532 305236 152584
rect 352288 152532 352340 152584
rect 346492 152464 346544 152516
rect 350540 152464 350592 152516
rect 356888 152532 356940 152584
rect 386972 152668 387024 152720
rect 389180 152668 389232 152720
rect 416504 152668 416556 152720
rect 417700 152668 417752 152720
rect 438308 152668 438360 152720
rect 485872 152668 485924 152720
rect 488448 152668 488500 152720
rect 357992 152600 358044 152652
rect 360016 152600 360068 152652
rect 361488 152600 361540 152652
rect 395344 152600 395396 152652
rect 395436 152600 395488 152652
rect 397828 152600 397880 152652
rect 402612 152600 402664 152652
rect 426808 152600 426860 152652
rect 430304 152600 430356 152652
rect 447968 152600 448020 152652
rect 388260 152532 388312 152584
rect 395896 152532 395948 152584
rect 421656 152532 421708 152584
rect 426164 152532 426216 152584
rect 444748 152532 444800 152584
rect 355232 152464 355284 152516
rect 384396 152464 384448 152516
rect 384948 152464 385000 152516
rect 413100 152464 413152 152516
rect 415216 152464 415268 152516
rect 436376 152464 436428 152516
rect 477592 152464 477644 152516
rect 480076 152464 480128 152516
rect 86868 152396 86920 152448
rect 185308 152396 185360 152448
rect 188988 152396 189040 152448
rect 193036 152396 193088 152448
rect 195980 152396 196032 152448
rect 198188 152396 198240 152448
rect 203616 152396 203668 152448
rect 274548 152396 274600 152448
rect 274640 152396 274692 152448
rect 282276 152396 282328 152448
rect 282920 152396 282972 152448
rect 288072 152396 288124 152448
rect 288164 152396 288216 152448
rect 336188 152396 336240 152448
rect 338764 152396 338816 152448
rect 377956 152396 378008 152448
rect 378232 152396 378284 152448
rect 408132 152396 408184 152448
rect 408868 152396 408920 152448
rect 428648 152396 428700 152448
rect 428740 152396 428792 152448
rect 446680 152396 446732 152448
rect 50344 152328 50396 152380
rect 146760 152328 146812 152380
rect 161204 152328 161256 152380
rect 169944 152328 169996 152380
rect 173256 152328 173308 152380
rect 243544 152328 243596 152380
rect 248144 152328 248196 152380
rect 252100 152328 252152 152380
rect 252560 152328 252612 152380
rect 306012 152328 306064 152380
rect 310612 152328 310664 152380
rect 313740 152328 313792 152380
rect 313832 152328 313884 152380
rect 318984 152328 319036 152380
rect 319352 152328 319404 152380
rect 361948 152328 362000 152380
rect 362684 152328 362736 152380
rect 365168 152328 365220 152380
rect 377220 152328 377272 152380
rect 381820 152328 381872 152380
rect 384120 152328 384172 152380
rect 412640 152328 412692 152380
rect 415492 152328 415544 152380
rect 419080 152328 419132 152380
rect 419172 152328 419224 152380
rect 429292 152328 429344 152380
rect 429476 152328 429528 152380
rect 447324 152328 447376 152380
rect 100300 152260 100352 152312
rect 195612 152260 195664 152312
rect 204444 152260 204496 152312
rect 275192 152260 275244 152312
rect 279516 152260 279568 152312
rect 282920 152260 282972 152312
rect 107016 152192 107068 152244
rect 200764 152192 200816 152244
rect 213092 152192 213144 152244
rect 216128 152192 216180 152244
rect 110328 152124 110380 152176
rect 203340 152124 203392 152176
rect 210332 152124 210384 152176
rect 6092 152056 6144 152108
rect 80612 152056 80664 152108
rect 81716 152056 81768 152108
rect 92480 152056 92532 152108
rect 105820 152056 105872 152108
rect 116492 152056 116544 152108
rect 119620 152056 119672 152108
rect 210424 152056 210476 152108
rect 211160 152124 211212 152176
rect 280344 152192 280396 152244
rect 281448 152192 281500 152244
rect 292764 152260 292816 152312
rect 284392 152192 284444 152244
rect 288164 152192 288216 152244
rect 290924 152192 290976 152244
rect 341340 152260 341392 152312
rect 342168 152260 342220 152312
rect 344560 152260 344612 152312
rect 344652 152260 344704 152312
rect 379888 152260 379940 152312
rect 380992 152260 381044 152312
rect 392124 152260 392176 152312
rect 392308 152260 392360 152312
rect 417792 152260 417844 152312
rect 293132 152192 293184 152244
rect 295064 152192 295116 152244
rect 279700 152124 279752 152176
rect 282460 152124 282512 152176
rect 295524 152192 295576 152244
rect 340696 152192 340748 152244
rect 340788 152192 340840 152244
rect 377312 152192 377364 152244
rect 380900 152192 380952 152244
rect 389548 152192 389600 152244
rect 390928 152192 390980 152244
rect 415216 152192 415268 152244
rect 331128 152124 331180 152176
rect 333980 152124 334032 152176
rect 372804 152124 372856 152176
rect 388536 152124 388588 152176
rect 410064 152124 410116 152176
rect 411720 152124 411772 152176
rect 431224 152260 431276 152312
rect 423220 152192 423272 152244
rect 217048 152056 217100 152108
rect 284852 152056 284904 152108
rect 287336 152056 287388 152108
rect 290004 152056 290056 152108
rect 290096 152056 290148 152108
rect 295340 152056 295392 152108
rect 47308 151988 47360 152040
rect 110052 151988 110104 152040
rect 123392 151988 123444 152040
rect 128176 151988 128228 152040
rect 128452 151988 128504 152040
rect 213552 151988 213604 152040
rect 214380 151988 214432 152040
rect 221280 151988 221332 152040
rect 223580 151988 223632 152040
rect 226432 151988 226484 152040
rect 54208 151920 54260 151972
rect 116676 151920 116728 151972
rect 125692 151920 125744 151972
rect 40500 151852 40552 151904
rect 109960 151852 110012 151904
rect 110144 151852 110196 151904
rect 126888 151852 126940 151904
rect 139768 151920 139820 151972
rect 142620 151920 142672 151972
rect 223856 151920 223908 151972
rect 224592 151920 224644 151972
rect 290648 151988 290700 152040
rect 292764 151988 292816 152040
rect 295156 151988 295208 152040
rect 295248 151988 295300 152040
rect 341984 152056 342036 152108
rect 342076 152056 342128 152108
rect 344652 152056 344704 152108
rect 345480 152056 345532 152108
rect 296812 151988 296864 152040
rect 345848 151988 345900 152040
rect 347136 152056 347188 152108
rect 355232 152056 355284 152108
rect 355324 152056 355376 152108
rect 383108 152056 383160 152108
rect 388444 152056 388496 152108
rect 404912 152056 404964 152108
rect 405004 152056 405056 152108
rect 423588 152056 423640 152108
rect 425244 152192 425296 152244
rect 444104 152260 444156 152312
rect 508412 152192 508464 152244
rect 509148 152192 509200 152244
rect 439596 152124 439648 152176
rect 347228 151988 347280 152040
rect 348056 151988 348108 152040
rect 385040 151988 385092 152040
rect 385684 151988 385736 152040
rect 399760 151988 399812 152040
rect 407304 151988 407356 152040
rect 426164 151988 426216 152040
rect 430580 151988 430632 152040
rect 431776 151988 431828 152040
rect 488540 151988 488592 152040
rect 490932 151988 490984 152040
rect 226984 151920 227036 151972
rect 128544 151852 128596 151904
rect 208492 151852 208544 151904
rect 208676 151852 208728 151904
rect 211068 151852 211120 151904
rect 227812 151852 227864 151904
rect 231584 151852 231636 151904
rect 233976 151920 234028 151972
rect 262680 151920 262732 151972
rect 262772 151920 262824 151972
rect 267556 151920 267608 151972
rect 269028 151920 269080 151972
rect 277124 151920 277176 151972
rect 277216 151920 277268 151972
rect 316592 151920 316644 151972
rect 77116 151784 77168 151836
rect 128084 151784 128136 151836
rect 128268 151784 128320 151836
rect 167552 151784 167604 151836
rect 167644 151784 167696 151836
rect 172520 151784 172572 151836
rect 96528 151716 96580 151768
rect 190736 151716 190788 151768
rect 97724 151648 97776 151700
rect 190920 151716 190972 151768
rect 191748 151716 191800 151768
rect 194600 151784 194652 151836
rect 254676 151784 254728 151836
rect 290004 151852 290056 151904
rect 290096 151852 290148 151904
rect 297732 151852 297784 151904
rect 297824 151852 297876 151904
rect 302516 151852 302568 151904
rect 323676 151920 323728 151972
rect 326804 151920 326856 151972
rect 332784 151920 332836 151972
rect 367008 151920 367060 151972
rect 386236 151920 386288 151972
rect 397184 151920 397236 151972
rect 398104 151920 398156 151972
rect 405556 151920 405608 151972
rect 405648 151920 405700 151972
rect 421012 151920 421064 151972
rect 422576 151920 422628 151972
rect 437020 151920 437072 151972
rect 479524 151920 479576 151972
rect 481364 151920 481416 151972
rect 507032 151920 507084 151972
rect 507584 151920 507636 151972
rect 262864 151784 262916 151836
rect 270132 151784 270184 151836
rect 271512 151784 271564 151836
rect 274640 151784 274692 151836
rect 274732 151784 274784 151836
rect 292580 151784 292632 151836
rect 293960 151784 294012 151836
rect 298376 151784 298428 151836
rect 298468 151784 298520 151836
rect 306380 151784 306432 151836
rect 316684 151784 316736 151836
rect 193680 151716 193732 151768
rect 191012 151648 191064 151700
rect 195060 151648 195112 151700
rect 85396 151580 85448 151632
rect 183376 151580 183428 151632
rect 186228 151580 186280 151632
rect 191104 151580 191156 151632
rect 191932 151580 191984 151632
rect 265624 151716 265676 151768
rect 316592 151716 316644 151768
rect 325976 151784 326028 151836
rect 326068 151784 326120 151836
rect 328552 151784 328604 151836
rect 332692 151784 332744 151836
rect 334348 151784 334400 151836
rect 337844 151784 337896 151836
rect 338764 151784 338816 151836
rect 344928 151852 344980 151904
rect 349712 151852 349764 151904
rect 347136 151784 347188 151836
rect 347228 151784 347280 151836
rect 355324 151784 355376 151836
rect 358912 151784 358964 151836
rect 393412 151852 393464 151904
rect 396448 151852 396500 151904
rect 402980 151852 403032 151904
rect 398840 151784 398892 151836
rect 402244 151784 402296 151836
rect 415860 151852 415912 151904
rect 420184 151852 420236 151904
rect 434444 151852 434496 151904
rect 449992 151852 450044 151904
rect 451832 151852 451884 151904
rect 459560 151852 459612 151904
rect 462044 151852 462096 151904
rect 477684 151852 477736 151904
rect 480720 151852 480772 151904
rect 488908 151852 488960 151904
rect 490288 151852 490340 151904
rect 410708 151784 410760 151836
rect 416688 151784 416740 151836
rect 424232 151784 424284 151836
rect 196072 151648 196124 151700
rect 268844 151648 268896 151700
rect 198556 151580 198608 151632
rect 270776 151580 270828 151632
rect 91008 151512 91060 151564
rect 188528 151512 188580 151564
rect 188620 151512 188672 151564
rect 263048 151512 263100 151564
rect 82728 151444 82780 151496
rect 181444 151444 181496 151496
rect 181996 151444 182048 151496
rect 257896 151444 257948 151496
rect 74264 151376 74316 151428
rect 175556 151376 175608 151428
rect 175648 151376 175700 151428
rect 191012 151376 191064 151428
rect 191104 151376 191156 151428
rect 261116 151376 261168 151428
rect 71688 151308 71740 151360
rect 173808 151308 173860 151360
rect 175188 151308 175240 151360
rect 252744 151308 252796 151360
rect 24676 151240 24728 151292
rect 137836 151240 137888 151292
rect 155684 151240 155736 151292
rect 237380 151240 237432 151292
rect 263508 151240 263560 151292
rect 320180 151240 320232 151292
rect 19248 151172 19300 151224
rect 132684 151172 132736 151224
rect 137284 151172 137336 151224
rect 220636 151172 220688 151224
rect 256424 151172 256476 151224
rect 315028 151172 315080 151224
rect 12348 151104 12400 151156
rect 127532 151104 127584 151156
rect 135168 151104 135220 151156
rect 221924 151104 221976 151156
rect 246396 151104 246448 151156
rect 307300 151104 307352 151156
rect 5356 151036 5408 151088
rect 123024 151036 123076 151088
rect 127992 151036 128044 151088
rect 216772 151036 216824 151088
rect 223488 151036 223540 151088
rect 289360 151036 289412 151088
rect 102048 150968 102100 151020
rect 196256 150968 196308 151020
rect 199384 150968 199436 151020
rect 271420 150968 271472 151020
rect 108948 150900 109000 150952
rect 201408 150900 201460 150952
rect 202696 150900 202748 150952
rect 273904 150900 273956 150952
rect 43904 150832 43956 150884
rect 116860 150832 116912 150884
rect 95516 150764 95568 150816
rect 110328 150764 110380 150816
rect 115756 150764 115808 150816
rect 206560 150832 206612 150884
rect 209412 150832 209464 150884
rect 279056 150832 279108 150884
rect 118608 150764 118660 150816
rect 209136 150764 209188 150816
rect 92020 150696 92072 150748
rect 111524 150696 111576 150748
rect 121368 150696 121420 150748
rect 211620 150696 211672 150748
rect 88616 150628 88668 150680
rect 111432 150628 111484 150680
rect 116768 150628 116820 150680
rect 85212 150560 85264 150612
rect 117228 150560 117280 150612
rect 50804 150492 50856 150544
rect 116952 150492 117004 150544
rect 168288 150628 168340 150680
rect 247592 150628 247644 150680
rect 164976 150560 165028 150612
rect 245016 150560 245068 150612
rect 194968 150492 195020 150544
rect 195060 150492 195112 150544
rect 238668 150492 238720 150544
rect 98920 150424 98972 150476
rect 111248 150424 111300 150476
rect 117136 150424 117188 150476
rect 179604 150424 179656 150476
rect 180064 150424 180116 150476
rect 251456 150424 251508 150476
rect 78312 150356 78364 150408
rect 114100 150356 114152 150408
rect 74816 150288 74868 150340
rect 114008 150288 114060 150340
rect 71412 150220 71464 150272
rect 115204 150220 115256 150272
rect 102600 150152 102652 150204
rect 116032 150152 116084 150204
rect 147680 150152 147732 150204
rect 148830 150152 148882 150204
rect 218244 150152 218296 150204
rect 219394 150152 219446 150204
rect 265164 150152 265216 150204
rect 266314 150152 266366 150204
rect 292488 150152 292540 150204
rect 293914 150152 293966 150204
rect 394884 150152 394936 150204
rect 396034 150152 396086 150204
rect 451372 150152 451424 150204
rect 452522 150152 452574 150204
rect 455420 150152 455472 150204
rect 456386 150152 456438 150204
rect 456800 150152 456852 150204
rect 457674 150152 457726 150204
rect 462320 150152 462372 150204
rect 463378 150152 463430 150204
rect 468024 150152 468076 150204
rect 469174 150152 469226 150204
rect 471980 150152 472032 150204
rect 473038 150152 473090 150204
rect 496912 150152 496964 150204
rect 498062 150152 498114 150204
rect 500960 150152 501012 150204
rect 501926 150152 501978 150204
rect 68008 150084 68060 150136
rect 92480 150084 92532 150136
rect 117136 150084 117188 150136
rect 202742 150084 202794 150136
rect 292396 150084 292448 150136
rect 299066 150084 299118 150136
rect 111064 150016 111116 150068
rect 111616 150016 111668 150068
rect 111156 148996 111208 149048
rect 116124 148996 116176 149048
rect 116676 146956 116728 147008
rect 117044 146956 117096 147008
rect 111248 143488 111300 143540
rect 116124 143488 116176 143540
rect 111064 143148 111116 143200
rect 111432 143148 111484 143200
rect 111524 140700 111576 140752
rect 116124 140700 116176 140752
rect 111340 137912 111392 137964
rect 116124 137912 116176 137964
rect 114100 132132 114152 132184
rect 115940 132132 115992 132184
rect 114008 131044 114060 131096
rect 115940 131044 115992 131096
rect 111156 126896 111208 126948
rect 116124 126896 116176 126948
rect 112904 124108 112956 124160
rect 116124 124108 116176 124160
rect 112720 122748 112772 122800
rect 116124 122748 116176 122800
rect 112536 121388 112588 121440
rect 116124 121388 116176 121440
rect 112444 107584 112496 107636
rect 116124 107584 116176 107636
rect 111616 104796 111668 104848
rect 116124 104796 116176 104848
rect 111432 102076 111484 102128
rect 115940 102076 115992 102128
rect 111248 96568 111300 96620
rect 116124 96568 116176 96620
rect 111064 93780 111116 93832
rect 116124 93780 116176 93832
rect 113824 88272 113876 88324
rect 115940 88272 115992 88324
rect 113916 86912 113968 86964
rect 116400 86912 116452 86964
rect 114008 83920 114060 83972
rect 116584 83920 116636 83972
rect 114100 82764 114152 82816
rect 116308 82764 116360 82816
rect 114192 79976 114244 80028
rect 115940 79976 115992 80028
rect 114284 78616 114336 78668
rect 116216 78616 116268 78668
rect 114192 71748 114244 71800
rect 116584 71748 116636 71800
rect 114100 69028 114152 69080
rect 116308 69028 116360 69080
rect 114008 67600 114060 67652
rect 116124 67600 116176 67652
rect 113916 66240 113968 66292
rect 116584 66240 116636 66292
rect 113364 64676 113416 64728
rect 116584 64676 116636 64728
rect 113824 63520 113876 63572
rect 116216 63520 116268 63572
rect 112444 62092 112496 62144
rect 116124 62092 116176 62144
rect 112536 44140 112588 44192
rect 116124 44140 116176 44192
rect 112628 34484 112680 34536
rect 115940 34484 115992 34536
rect 114100 33124 114152 33176
rect 115940 33124 115992 33176
rect 112720 28976 112772 29028
rect 116124 28976 116176 29028
rect 112812 24828 112864 24880
rect 116124 24828 116176 24880
rect 114008 23468 114060 23520
rect 115940 23468 115992 23520
rect 112904 22108 112956 22160
rect 116124 22108 116176 22160
rect 116400 11704 116452 11756
rect 116860 11704 116912 11756
rect 116032 11636 116084 11688
rect 117044 11636 117096 11688
rect 111156 5516 111208 5568
rect 115940 5516 115992 5568
rect 111800 4156 111852 4208
rect 116124 4156 116176 4208
rect 111064 2796 111116 2848
rect 143632 2456 143684 2508
rect 425796 2456 425848 2508
rect 443644 2456 443696 2508
rect 102692 1912 102744 1964
rect 116584 1912 116636 1964
rect 92664 1844 92716 1896
rect 94412 1844 94464 1896
rect 95976 1844 96028 1896
rect 89352 1776 89404 1828
rect 105820 1776 105872 1828
rect 106004 1844 106056 1896
rect 109684 1844 109736 1896
rect 109040 1776 109092 1828
rect 109316 1776 109368 1828
rect 112444 1776 112496 1828
rect 65984 1708 66036 1760
rect 88892 1708 88944 1760
rect 99380 1708 99432 1760
rect 116676 1708 116728 1760
rect 86040 1640 86092 1692
rect 82636 1572 82688 1624
rect 105636 1572 105688 1624
rect 72700 1504 72752 1556
rect 100300 1504 100352 1556
rect 105820 1640 105872 1692
rect 105912 1640 105964 1692
rect 108948 1640 109000 1692
rect 109040 1640 109092 1692
rect 109776 1640 109828 1692
rect 109868 1572 109920 1624
rect 109960 1504 110012 1556
rect 110144 1504 110196 1556
rect 193588 1504 193640 1556
rect 32680 1436 32732 1488
rect 116400 1436 116452 1488
rect 29276 1368 29328 1420
rect 115940 1368 115992 1420
rect 294788 1368 294840 1420
rect 343640 1368 343692 1420
rect 491300 1368 491352 1420
rect 493600 1368 493652 1420
rect 2688 1300 2740 1352
rect 116124 1300 116176 1352
rect 6000 1232 6052 1284
rect 111800 1232 111852 1284
rect 9312 1164 9364 1216
rect 111156 1164 111208 1216
rect 35992 1096 36044 1148
rect 112904 1096 112956 1148
rect 39304 1028 39356 1080
rect 114008 1028 114060 1080
rect 42616 960 42668 1012
rect 112812 960 112864 1012
rect 46020 892 46072 944
rect 49332 824 49384 876
rect 112720 824 112772 876
rect 52644 756 52696 808
rect 59360 688 59412 740
rect 108212 688 108264 740
rect 62672 620 62724 672
rect 115388 756 115440 808
rect 108396 688 108448 740
rect 114100 688 114152 740
rect 69296 552 69348 604
rect 79324 484 79376 536
rect 112628 552 112680 604
rect 115296 552 115348 604
rect 115204 416 115256 468
rect 112536 348 112588 400
<< metal2 >>
rect 386 159200 442 160400
rect 1214 159200 1270 160400
rect 2042 159200 2098 160400
rect 2870 159200 2926 160400
rect 3698 159200 3754 160400
rect 4526 159200 4582 160400
rect 5354 159200 5410 160400
rect 6182 159200 6238 160400
rect 7102 159200 7158 160400
rect 7930 159202 7986 160400
rect 8036 159310 8248 159338
rect 8036 159202 8064 159310
rect 7930 159200 8064 159202
rect 400 156670 428 159200
rect 388 156664 440 156670
rect 388 156606 440 156612
rect 1228 153882 1256 159200
rect 1216 153876 1268 153882
rect 1216 153818 1268 153824
rect 2056 153785 2084 159200
rect 2884 155145 2912 159200
rect 3712 156738 3740 159200
rect 3700 156732 3752 156738
rect 3700 156674 3752 156680
rect 2870 155136 2926 155145
rect 2870 155071 2926 155080
rect 4540 153950 4568 159200
rect 4528 153944 4580 153950
rect 4528 153886 4580 153892
rect 2042 153776 2098 153785
rect 2042 153711 2098 153720
rect 2686 151872 2742 151881
rect 2686 151807 2742 151816
rect 2700 149940 2728 151807
rect 5368 151094 5396 159200
rect 6196 152425 6224 159200
rect 7116 156806 7144 159200
rect 7944 159174 8064 159200
rect 7104 156800 7156 156806
rect 7104 156742 7156 156748
rect 8220 156074 8248 159310
rect 8758 159200 8814 160400
rect 9586 159200 9642 160400
rect 10414 159200 10470 160400
rect 11242 159200 11298 160400
rect 12070 159200 12126 160400
rect 12898 159200 12954 160400
rect 13818 159200 13874 160400
rect 14646 159200 14702 160400
rect 15474 159200 15530 160400
rect 16302 159200 16358 160400
rect 17130 159200 17186 160400
rect 17958 159200 18014 160400
rect 18786 159200 18842 160400
rect 19614 159200 19670 160400
rect 20534 159200 20590 160400
rect 21362 159200 21418 160400
rect 22190 159200 22246 160400
rect 23018 159200 23074 160400
rect 23846 159200 23902 160400
rect 24674 159200 24730 160400
rect 25502 159200 25558 160400
rect 26330 159200 26386 160400
rect 27250 159200 27306 160400
rect 28078 159200 28134 160400
rect 28906 159200 28962 160400
rect 29734 159200 29790 160400
rect 30562 159200 30618 160400
rect 31390 159200 31446 160400
rect 32218 159200 32274 160400
rect 33138 159200 33194 160400
rect 33966 159200 34022 160400
rect 34794 159200 34850 160400
rect 35622 159200 35678 160400
rect 36450 159200 36506 160400
rect 37278 159200 37334 160400
rect 38106 159200 38162 160400
rect 38934 159200 38990 160400
rect 39854 159200 39910 160400
rect 40682 159200 40738 160400
rect 41510 159200 41566 160400
rect 42338 159200 42394 160400
rect 43166 159200 43222 160400
rect 43994 159200 44050 160400
rect 44822 159200 44878 160400
rect 45650 159200 45706 160400
rect 46570 159200 46626 160400
rect 47398 159200 47454 160400
rect 48226 159200 48282 160400
rect 49054 159200 49110 160400
rect 49882 159200 49938 160400
rect 50710 159200 50766 160400
rect 51538 159200 51594 160400
rect 52366 159200 52422 160400
rect 53286 159200 53342 160400
rect 54114 159200 54170 160400
rect 54942 159200 54998 160400
rect 55770 159200 55826 160400
rect 56598 159200 56654 160400
rect 57426 159200 57482 160400
rect 58254 159200 58310 160400
rect 59082 159200 59138 160400
rect 60002 159200 60058 160400
rect 60830 159200 60886 160400
rect 61658 159200 61714 160400
rect 62486 159200 62542 160400
rect 63314 159200 63370 160400
rect 64142 159200 64198 160400
rect 64970 159200 65026 160400
rect 65890 159200 65946 160400
rect 66718 159200 66774 160400
rect 67546 159200 67602 160400
rect 68374 159200 68430 160400
rect 69202 159200 69258 160400
rect 70030 159200 70086 160400
rect 70858 159200 70914 160400
rect 71686 159200 71742 160400
rect 72606 159200 72662 160400
rect 73434 159200 73490 160400
rect 74262 159200 74318 160400
rect 75090 159200 75146 160400
rect 75918 159200 75974 160400
rect 76746 159200 76802 160400
rect 77574 159200 77630 160400
rect 78402 159200 78458 160400
rect 79322 159200 79378 160400
rect 80150 159200 80206 160400
rect 80978 159200 81034 160400
rect 81806 159200 81862 160400
rect 82634 159200 82690 160400
rect 83462 159200 83518 160400
rect 84290 159200 84346 160400
rect 85118 159200 85174 160400
rect 86038 159200 86094 160400
rect 86866 159200 86922 160400
rect 87694 159200 87750 160400
rect 88522 159200 88578 160400
rect 89350 159200 89406 160400
rect 90178 159200 90234 160400
rect 91006 159200 91062 160400
rect 91834 159200 91890 160400
rect 92754 159200 92810 160400
rect 93582 159200 93638 160400
rect 94410 159200 94466 160400
rect 95238 159200 95294 160400
rect 96066 159200 96122 160400
rect 96894 159200 96950 160400
rect 97722 159200 97778 160400
rect 98642 159200 98698 160400
rect 99470 159200 99526 160400
rect 100298 159200 100354 160400
rect 101126 159200 101182 160400
rect 101954 159200 102010 160400
rect 102782 159200 102838 160400
rect 103610 159200 103666 160400
rect 104438 159200 104494 160400
rect 105358 159200 105414 160400
rect 106186 159200 106242 160400
rect 107014 159200 107070 160400
rect 107842 159200 107898 160400
rect 108670 159200 108726 160400
rect 109498 159200 109554 160400
rect 110326 159200 110382 160400
rect 111154 159200 111210 160400
rect 112074 159200 112130 160400
rect 112902 159200 112958 160400
rect 113730 159200 113786 160400
rect 114558 159200 114614 160400
rect 115386 159200 115442 160400
rect 116214 159200 116270 160400
rect 117042 159200 117098 160400
rect 117870 159200 117926 160400
rect 118790 159200 118846 160400
rect 119618 159200 119674 160400
rect 120446 159200 120502 160400
rect 121274 159200 121330 160400
rect 122102 159200 122158 160400
rect 122930 159200 122986 160400
rect 123758 159200 123814 160400
rect 124586 159200 124642 160400
rect 125506 159200 125562 160400
rect 126334 159200 126390 160400
rect 127162 159200 127218 160400
rect 127990 159200 128046 160400
rect 128818 159200 128874 160400
rect 129646 159200 129702 160400
rect 130474 159200 130530 160400
rect 131394 159200 131450 160400
rect 132222 159200 132278 160400
rect 133050 159200 133106 160400
rect 133878 159200 133934 160400
rect 134706 159200 134762 160400
rect 135534 159200 135590 160400
rect 136362 159200 136418 160400
rect 137190 159200 137246 160400
rect 138110 159200 138166 160400
rect 138938 159200 138994 160400
rect 139766 159200 139822 160400
rect 140594 159200 140650 160400
rect 141422 159200 141478 160400
rect 142250 159200 142306 160400
rect 143078 159200 143134 160400
rect 143906 159200 143962 160400
rect 144826 159200 144882 160400
rect 145654 159200 145710 160400
rect 146482 159200 146538 160400
rect 147310 159200 147366 160400
rect 148138 159200 148194 160400
rect 148966 159200 149022 160400
rect 149794 159200 149850 160400
rect 150622 159200 150678 160400
rect 151542 159200 151598 160400
rect 152370 159200 152426 160400
rect 153198 159200 153254 160400
rect 154026 159200 154082 160400
rect 154854 159200 154910 160400
rect 155682 159200 155738 160400
rect 156510 159200 156566 160400
rect 157338 159200 157394 160400
rect 158258 159200 158314 160400
rect 159086 159200 159142 160400
rect 159914 159200 159970 160400
rect 160742 159200 160798 160400
rect 161570 159200 161626 160400
rect 162398 159200 162454 160400
rect 163226 159200 163282 160400
rect 164146 159200 164202 160400
rect 164974 159200 165030 160400
rect 165802 159200 165858 160400
rect 166630 159200 166686 160400
rect 167458 159200 167514 160400
rect 168286 159200 168342 160400
rect 169114 159200 169170 160400
rect 169942 159200 169998 160400
rect 170862 159200 170918 160400
rect 171690 159200 171746 160400
rect 172518 159200 172574 160400
rect 173346 159200 173402 160400
rect 174174 159200 174230 160400
rect 175002 159200 175058 160400
rect 175830 159200 175886 160400
rect 176658 159200 176714 160400
rect 177578 159200 177634 160400
rect 178406 159200 178462 160400
rect 179234 159200 179290 160400
rect 180062 159200 180118 160400
rect 180890 159200 180946 160400
rect 181718 159202 181774 160400
rect 181824 159310 182036 159338
rect 181824 159202 181852 159310
rect 181718 159200 181852 159202
rect 8298 156088 8354 156097
rect 8220 156046 8298 156074
rect 8298 156023 8354 156032
rect 8772 153610 8800 159200
rect 9600 155281 9628 159200
rect 10428 155446 10456 159200
rect 10416 155440 10468 155446
rect 10416 155382 10468 155388
rect 11256 155378 11284 159200
rect 12084 155718 12112 159200
rect 12072 155712 12124 155718
rect 12072 155654 12124 155660
rect 11244 155372 11296 155378
rect 11244 155314 11296 155320
rect 12348 155372 12400 155378
rect 12348 155314 12400 155320
rect 9586 155272 9642 155281
rect 9586 155207 9642 155216
rect 8760 153604 8812 153610
rect 8760 153546 8812 153552
rect 6182 152416 6238 152425
rect 6182 152351 6238 152360
rect 6092 152108 6144 152114
rect 6092 152050 6144 152056
rect 5356 151088 5408 151094
rect 5356 151030 5408 151036
rect 6104 149940 6132 152050
rect 9494 151464 9550 151473
rect 9494 151399 9550 151408
rect 9508 149940 9536 151399
rect 12360 151162 12388 155314
rect 12912 152522 12940 159200
rect 13832 154086 13860 159200
rect 14660 156874 14688 159200
rect 14648 156868 14700 156874
rect 14648 156810 14700 156816
rect 15488 155922 15516 159200
rect 15476 155916 15528 155922
rect 15476 155858 15528 155864
rect 16316 155553 16344 159200
rect 16302 155544 16358 155553
rect 16302 155479 16358 155488
rect 13820 154080 13872 154086
rect 13820 154022 13872 154028
rect 17144 154018 17172 159200
rect 17972 155242 18000 159200
rect 17960 155236 18012 155242
rect 17960 155178 18012 155184
rect 17132 154012 17184 154018
rect 17132 153954 17184 153960
rect 18800 152561 18828 159200
rect 19248 155236 19300 155242
rect 19248 155178 19300 155184
rect 18786 152552 18842 152561
rect 12900 152516 12952 152522
rect 18786 152487 18842 152496
rect 12900 152458 12952 152464
rect 16394 152008 16450 152017
rect 16394 151943 16450 151952
rect 12348 151156 12400 151162
rect 12348 151098 12400 151104
rect 12990 150648 13046 150657
rect 12990 150583 13046 150592
rect 13004 149940 13032 150583
rect 16408 149940 16436 151943
rect 19260 151230 19288 155178
rect 19628 152697 19656 159200
rect 20548 153921 20576 159200
rect 21376 156942 21404 159200
rect 21364 156936 21416 156942
rect 21364 156878 21416 156884
rect 22204 155242 22232 159200
rect 23032 155689 23060 159200
rect 23860 157010 23888 159200
rect 23848 157004 23900 157010
rect 23848 156946 23900 156952
rect 23018 155680 23074 155689
rect 23018 155615 23074 155624
rect 22192 155236 22244 155242
rect 22192 155178 22244 155184
rect 20534 153912 20590 153921
rect 20534 153847 20590 153856
rect 19614 152688 19670 152697
rect 19614 152623 19670 152632
rect 24688 151298 24716 159200
rect 25516 152590 25544 159200
rect 26344 152726 26372 159200
rect 27264 153474 27292 159200
rect 28092 157078 28120 159200
rect 28080 157072 28132 157078
rect 28080 157014 28132 157020
rect 28920 155961 28948 159200
rect 28906 155952 28962 155961
rect 28906 155887 28962 155896
rect 29748 155825 29776 159200
rect 29734 155816 29790 155825
rect 29734 155751 29790 155760
rect 30576 154154 30604 159200
rect 31404 158574 31432 159200
rect 31392 158568 31444 158574
rect 31392 158510 31444 158516
rect 30564 154148 30616 154154
rect 30564 154090 30616 154096
rect 27252 153468 27304 153474
rect 27252 153410 27304 153416
rect 26332 152720 26384 152726
rect 26332 152662 26384 152668
rect 32232 152658 32260 159200
rect 33152 152794 33180 159200
rect 33980 156641 34008 159200
rect 33966 156632 34022 156641
rect 33966 156567 34022 156576
rect 34808 154290 34836 159200
rect 35636 157486 35664 159200
rect 35624 157480 35676 157486
rect 35624 157422 35676 157428
rect 36464 155378 36492 159200
rect 37292 157214 37320 159200
rect 37280 157208 37332 157214
rect 37280 157150 37332 157156
rect 36452 155372 36504 155378
rect 36452 155314 36504 155320
rect 34796 154284 34848 154290
rect 34796 154226 34848 154232
rect 38120 154222 38148 159200
rect 38948 157554 38976 159200
rect 38936 157548 38988 157554
rect 38936 157490 38988 157496
rect 39868 155310 39896 159200
rect 40696 157146 40724 159200
rect 40684 157140 40736 157146
rect 40684 157082 40736 157088
rect 39856 155304 39908 155310
rect 39856 155246 39908 155252
rect 41524 154358 41552 159200
rect 42352 157622 42380 159200
rect 42340 157616 42392 157622
rect 42340 157558 42392 157564
rect 41512 154352 41564 154358
rect 41512 154294 41564 154300
rect 38108 154216 38160 154222
rect 38108 154158 38160 154164
rect 43180 152862 43208 159200
rect 44008 157282 44036 159200
rect 43996 157276 44048 157282
rect 43996 157218 44048 157224
rect 44836 154057 44864 159200
rect 45664 157758 45692 159200
rect 45652 157752 45704 157758
rect 45652 157694 45704 157700
rect 44822 154048 44878 154057
rect 44822 153983 44878 153992
rect 46584 152930 46612 159200
rect 47412 157350 47440 159200
rect 47400 157344 47452 157350
rect 47400 157286 47452 157292
rect 48240 154426 48268 159200
rect 49068 157690 49096 159200
rect 49056 157684 49108 157690
rect 49056 157626 49108 157632
rect 49896 155650 49924 159200
rect 50724 156602 50752 159200
rect 50712 156596 50764 156602
rect 50712 156538 50764 156544
rect 49884 155644 49936 155650
rect 49884 155586 49936 155592
rect 50344 155372 50396 155378
rect 50344 155314 50396 155320
rect 48228 154420 48280 154426
rect 48228 154362 48280 154368
rect 46572 152924 46624 152930
rect 46572 152866 46624 152872
rect 43168 152856 43220 152862
rect 43168 152798 43220 152804
rect 33140 152788 33192 152794
rect 33140 152730 33192 152736
rect 32220 152652 32272 152658
rect 32220 152594 32272 152600
rect 25504 152584 25556 152590
rect 25504 152526 25556 152532
rect 50356 152386 50384 155314
rect 51552 154562 51580 159200
rect 52380 157826 52408 159200
rect 52368 157820 52420 157826
rect 52368 157762 52420 157768
rect 53300 155378 53328 159200
rect 54128 156534 54156 159200
rect 54116 156528 54168 156534
rect 54116 156470 54168 156476
rect 53288 155372 53340 155378
rect 53288 155314 53340 155320
rect 51540 154556 51592 154562
rect 51540 154498 51592 154504
rect 54956 154494 54984 159200
rect 55784 157894 55812 159200
rect 55772 157888 55824 157894
rect 55772 157830 55824 157836
rect 54944 154488 54996 154494
rect 54944 154430 54996 154436
rect 56612 152998 56640 159200
rect 57440 154970 57468 159200
rect 57428 154964 57480 154970
rect 57428 154906 57480 154912
rect 58268 153814 58296 159200
rect 59096 157962 59124 159200
rect 59084 157956 59136 157962
rect 59084 157898 59136 157904
rect 60016 155582 60044 159200
rect 60844 156466 60872 159200
rect 60832 156460 60884 156466
rect 60832 156402 60884 156408
rect 60004 155576 60056 155582
rect 60004 155518 60056 155524
rect 61672 154193 61700 159200
rect 62500 158030 62528 159200
rect 62488 158024 62540 158030
rect 62488 157966 62540 157972
rect 61658 154184 61714 154193
rect 61658 154119 61714 154128
rect 58256 153808 58308 153814
rect 58256 153750 58308 153756
rect 63328 153066 63356 159200
rect 64156 155038 64184 159200
rect 64144 155032 64196 155038
rect 64144 154974 64196 154980
rect 64984 153678 65012 159200
rect 65904 158098 65932 159200
rect 65892 158092 65944 158098
rect 65892 158034 65944 158040
rect 66732 155786 66760 159200
rect 66720 155780 66772 155786
rect 66720 155722 66772 155728
rect 64972 153672 65024 153678
rect 64972 153614 65024 153620
rect 63316 153060 63368 153066
rect 63316 153002 63368 153008
rect 56600 152992 56652 152998
rect 56600 152934 56652 152940
rect 50344 152380 50396 152386
rect 50344 152322 50396 152328
rect 37002 152144 37058 152153
rect 37002 152079 37058 152088
rect 33598 151600 33654 151609
rect 33598 151535 33654 151544
rect 24676 151292 24728 151298
rect 24676 151234 24728 151240
rect 19248 151224 19300 151230
rect 19248 151166 19300 151172
rect 30194 151192 30250 151201
rect 30194 151127 30250 151136
rect 23294 150920 23350 150929
rect 23294 150855 23350 150864
rect 19798 150784 19854 150793
rect 19798 150719 19854 150728
rect 19812 149940 19840 150719
rect 23308 149940 23336 150855
rect 30208 149940 30236 151127
rect 33612 149940 33640 151535
rect 37016 149940 37044 152079
rect 47308 152040 47360 152046
rect 47308 151982 47360 151988
rect 40500 151904 40552 151910
rect 40500 151846 40552 151852
rect 40512 149940 40540 151846
rect 43904 150884 43956 150890
rect 43904 150826 43956 150832
rect 43916 149940 43944 150826
rect 47320 149940 47348 151982
rect 54208 151972 54260 151978
rect 54208 151914 54260 151920
rect 50804 150544 50856 150550
rect 50804 150486 50856 150492
rect 50816 149940 50844 150486
rect 54220 149940 54248 151914
rect 67560 151065 67588 159200
rect 68388 153746 68416 159200
rect 69216 158234 69244 159200
rect 69204 158228 69256 158234
rect 69204 158170 69256 158176
rect 70044 155514 70072 159200
rect 70872 156398 70900 159200
rect 70860 156392 70912 156398
rect 70860 156334 70912 156340
rect 70032 155508 70084 155514
rect 70032 155450 70084 155456
rect 68376 153740 68428 153746
rect 68376 153682 68428 153688
rect 71700 151366 71728 159200
rect 72620 158166 72648 159200
rect 72608 158160 72660 158166
rect 72608 158102 72660 158108
rect 73448 153134 73476 159200
rect 73436 153128 73488 153134
rect 73436 153070 73488 153076
rect 74276 151434 74304 159200
rect 75104 153542 75132 159200
rect 75932 158302 75960 159200
rect 75920 158296 75972 158302
rect 75920 158238 75972 158244
rect 76760 155854 76788 159200
rect 77588 155990 77616 159200
rect 78416 156330 78444 159200
rect 78404 156324 78456 156330
rect 78404 156266 78456 156272
rect 77576 155984 77628 155990
rect 77576 155926 77628 155932
rect 76748 155848 76800 155854
rect 76748 155790 76800 155796
rect 77116 155712 77168 155718
rect 77116 155654 77168 155660
rect 75092 153536 75144 153542
rect 75092 153478 75144 153484
rect 77128 151842 77156 155654
rect 79336 154902 79364 159200
rect 79324 154896 79376 154902
rect 79324 154838 79376 154844
rect 80164 153202 80192 159200
rect 80992 156262 81020 159200
rect 80980 156256 81032 156262
rect 80980 156198 81032 156204
rect 81820 155718 81848 159200
rect 82648 158370 82676 159200
rect 82636 158364 82688 158370
rect 82636 158306 82688 158312
rect 83476 155854 83504 159200
rect 84304 155922 84332 159200
rect 84200 155916 84252 155922
rect 84200 155858 84252 155864
rect 84292 155916 84344 155922
rect 84292 155858 84344 155864
rect 83464 155848 83516 155854
rect 82832 155786 83044 155802
rect 83464 155790 83516 155796
rect 82820 155780 83056 155786
rect 82872 155774 83004 155780
rect 82820 155722 82872 155728
rect 83004 155722 83056 155728
rect 81808 155712 81860 155718
rect 81808 155654 81860 155660
rect 82728 155712 82780 155718
rect 82728 155654 82780 155660
rect 80152 153196 80204 153202
rect 80152 153138 80204 153144
rect 80612 152108 80664 152114
rect 80612 152050 80664 152056
rect 81716 152108 81768 152114
rect 81716 152050 81768 152056
rect 77116 151836 77168 151842
rect 77116 151778 77168 151784
rect 74264 151428 74316 151434
rect 74264 151370 74316 151376
rect 71688 151360 71740 151366
rect 71688 151302 71740 151308
rect 67546 151056 67602 151065
rect 67546 150991 67602 151000
rect 78312 150408 78364 150414
rect 78312 150350 78364 150356
rect 74816 150340 74868 150346
rect 74816 150282 74868 150288
rect 71412 150272 71464 150278
rect 71412 150214 71464 150220
rect 68008 150136 68060 150142
rect 68008 150078 68060 150084
rect 68020 149940 68048 150078
rect 71424 149940 71452 150214
rect 74828 149940 74856 150282
rect 78324 149940 78352 150350
rect 80624 149705 80652 152050
rect 81728 149940 81756 152050
rect 82740 151502 82768 155654
rect 84212 155106 84240 155858
rect 84200 155100 84252 155106
rect 84200 155042 84252 155048
rect 85132 153406 85160 159200
rect 85396 155916 85448 155922
rect 85396 155858 85448 155864
rect 85120 153400 85172 153406
rect 85120 153342 85172 153348
rect 85408 151638 85436 155858
rect 86052 154834 86080 159200
rect 86040 154828 86092 154834
rect 86040 154770 86092 154776
rect 86880 152454 86908 159200
rect 87708 156126 87736 159200
rect 87696 156120 87748 156126
rect 87696 156062 87748 156068
rect 88536 153338 88564 159200
rect 89364 158438 89392 159200
rect 89352 158432 89404 158438
rect 89352 158374 89404 158380
rect 90192 155174 90220 159200
rect 90180 155168 90232 155174
rect 90180 155110 90232 155116
rect 88524 153332 88576 153338
rect 88524 153274 88576 153280
rect 86868 152448 86920 152454
rect 86868 152390 86920 152396
rect 85396 151632 85448 151638
rect 85396 151574 85448 151580
rect 91020 151570 91048 159200
rect 91848 156777 91876 159200
rect 91834 156768 91890 156777
rect 91834 156703 91890 156712
rect 91100 155100 91152 155106
rect 91100 155042 91152 155048
rect 91112 153105 91140 155042
rect 92768 154630 92796 159200
rect 92756 154624 92808 154630
rect 92756 154566 92808 154572
rect 91098 153096 91154 153105
rect 91098 153031 91154 153040
rect 93596 152833 93624 159200
rect 94424 156058 94452 159200
rect 94412 156052 94464 156058
rect 94412 155994 94464 156000
rect 95252 155922 95280 159200
rect 96080 158506 96108 159200
rect 96068 158500 96120 158506
rect 96068 158442 96120 158448
rect 95240 155916 95292 155922
rect 95240 155858 95292 155864
rect 96528 155916 96580 155922
rect 96528 155858 96580 155864
rect 93582 152824 93638 152833
rect 93582 152759 93638 152768
rect 92480 152108 92532 152114
rect 92480 152050 92532 152056
rect 91008 151564 91060 151570
rect 91008 151506 91060 151512
rect 82728 151496 82780 151502
rect 82728 151438 82780 151444
rect 92020 150748 92072 150754
rect 92020 150690 92072 150696
rect 88616 150680 88668 150686
rect 88616 150622 88668 150628
rect 85212 150612 85264 150618
rect 85212 150554 85264 150560
rect 85224 149940 85252 150554
rect 88628 149940 88656 150622
rect 92032 149940 92060 150690
rect 92492 150142 92520 152050
rect 96540 151774 96568 155858
rect 96908 155106 96936 159200
rect 96896 155100 96948 155106
rect 96896 155042 96948 155048
rect 96528 151768 96580 151774
rect 96528 151710 96580 151716
rect 97736 151706 97764 159200
rect 98656 154329 98684 159200
rect 99484 154698 99512 159200
rect 99472 154692 99524 154698
rect 99472 154634 99524 154640
rect 98642 154320 98698 154329
rect 98642 154255 98698 154264
rect 100312 152318 100340 159200
rect 101140 155922 101168 159200
rect 101968 156913 101996 159200
rect 102796 157418 102824 159200
rect 102784 157412 102836 157418
rect 102784 157354 102836 157360
rect 101954 156904 102010 156913
rect 101954 156839 102010 156848
rect 101128 155916 101180 155922
rect 101128 155858 101180 155864
rect 102048 155916 102100 155922
rect 102048 155858 102100 155864
rect 100300 152312 100352 152318
rect 100300 152254 100352 152260
rect 97724 151700 97776 151706
rect 97724 151642 97776 151648
rect 102060 151026 102088 155858
rect 103624 154970 103652 159200
rect 104452 157049 104480 159200
rect 104438 157040 104494 157049
rect 104438 156975 104494 156984
rect 103520 154964 103572 154970
rect 103520 154906 103572 154912
rect 103612 154964 103664 154970
rect 103612 154906 103664 154912
rect 103532 154766 103560 154906
rect 103520 154760 103572 154766
rect 103520 154702 103572 154708
rect 105372 153270 105400 159200
rect 106200 155922 106228 159200
rect 106188 155916 106240 155922
rect 106188 155858 106240 155864
rect 105360 153264 105412 153270
rect 105360 153206 105412 153212
rect 107028 152250 107056 159200
rect 107856 155446 107884 159200
rect 107752 155440 107804 155446
rect 107750 155408 107752 155417
rect 107844 155440 107896 155446
rect 107804 155408 107806 155417
rect 107844 155382 107896 155388
rect 107750 155343 107806 155352
rect 108684 154465 108712 159200
rect 109512 155922 109540 159200
rect 109408 155916 109460 155922
rect 109408 155858 109460 155864
rect 109500 155916 109552 155922
rect 109500 155858 109552 155864
rect 108948 155440 109000 155446
rect 109040 155440 109092 155446
rect 108948 155382 109000 155388
rect 109038 155408 109040 155417
rect 109092 155408 109094 155417
rect 108670 154456 108726 154465
rect 108670 154391 108726 154400
rect 107016 152244 107068 152250
rect 107016 152186 107068 152192
rect 105820 152108 105872 152114
rect 105820 152050 105872 152056
rect 102048 151020 102100 151026
rect 102048 150962 102100 150968
rect 95516 150816 95568 150822
rect 95516 150758 95568 150764
rect 92480 150136 92532 150142
rect 92480 150078 92532 150084
rect 95528 149940 95556 150758
rect 98920 150476 98972 150482
rect 98920 150418 98972 150424
rect 98932 149940 98960 150418
rect 102600 150204 102652 150210
rect 102600 150146 102652 150152
rect 102612 149954 102640 150146
rect 102350 149926 102640 149954
rect 105832 149940 105860 152050
rect 108960 150958 108988 155382
rect 109038 155343 109094 155352
rect 109420 154766 109448 155858
rect 110144 155440 110196 155446
rect 110144 155382 110196 155388
rect 109132 154760 109184 154766
rect 109132 154702 109184 154708
rect 109408 154760 109460 154766
rect 109408 154702 109460 154708
rect 109040 153604 109092 153610
rect 109040 153546 109092 153552
rect 109052 152289 109080 153546
rect 109144 152969 109172 154702
rect 109130 152960 109186 152969
rect 109130 152895 109186 152904
rect 109038 152280 109094 152289
rect 109038 152215 109094 152224
rect 109866 152144 109922 152153
rect 109866 152079 109922 152088
rect 109682 151872 109738 151881
rect 109682 151807 109738 151816
rect 108948 150952 109000 150958
rect 108948 150894 109000 150900
rect 109222 150512 109278 150521
rect 109222 150447 109278 150456
rect 109236 149940 109264 150447
rect 80610 149696 80666 149705
rect 80610 149631 80666 149640
rect 64694 149560 64750 149569
rect 64538 149518 64694 149546
rect 64694 149495 64750 149504
rect 26974 149424 27030 149433
rect 26726 149382 26974 149410
rect 57886 149424 57942 149433
rect 57730 149382 57886 149410
rect 26974 149359 27030 149368
rect 61474 149424 61530 149433
rect 61134 149382 61474 149410
rect 57886 149359 57942 149368
rect 61474 149359 61530 149368
rect 109696 93854 109724 151807
rect 109774 150784 109830 150793
rect 109774 150719 109830 150728
rect 109788 103514 109816 150719
rect 109880 107658 109908 152079
rect 110052 152040 110104 152046
rect 110052 151982 110104 151988
rect 109960 151904 110012 151910
rect 109960 151846 110012 151852
rect 109972 110650 110000 151846
rect 110064 132494 110092 151982
rect 110156 151910 110184 155382
rect 110340 152182 110368 159200
rect 111168 155446 111196 159200
rect 111616 155916 111668 155922
rect 111616 155858 111668 155864
rect 111800 155916 111852 155922
rect 111800 155858 111852 155864
rect 111156 155440 111208 155446
rect 111156 155382 111208 155388
rect 110328 152176 110380 152182
rect 110328 152118 110380 152124
rect 110144 151904 110196 151910
rect 110144 151846 110196 151852
rect 110878 151464 110934 151473
rect 110878 151399 110934 151408
rect 110328 150816 110380 150822
rect 110328 150758 110380 150764
rect 110340 140865 110368 150758
rect 110892 142154 110920 151399
rect 110970 150920 111026 150929
rect 110970 150855 111026 150864
rect 110984 146010 111012 150855
rect 111524 150748 111576 150754
rect 111524 150690 111576 150696
rect 111432 150680 111484 150686
rect 111338 150648 111394 150657
rect 111432 150622 111484 150628
rect 111338 150583 111394 150592
rect 111154 150512 111210 150521
rect 111154 150447 111210 150456
rect 111248 150476 111300 150482
rect 111064 150068 111116 150074
rect 111064 150010 111116 150016
rect 111076 146146 111104 150010
rect 111168 149054 111196 150447
rect 111248 150418 111300 150424
rect 111156 149048 111208 149054
rect 111156 148990 111208 148996
rect 111076 146118 111196 146146
rect 110984 145982 111104 146010
rect 111076 143206 111104 145982
rect 111064 143200 111116 143206
rect 111064 143142 111116 143148
rect 110892 142126 111104 142154
rect 110326 140856 110382 140865
rect 110326 140791 110382 140800
rect 110064 132466 110368 132494
rect 110340 113257 110368 132466
rect 110326 113248 110382 113257
rect 110326 113183 110382 113192
rect 110326 110664 110382 110673
rect 109972 110622 110326 110650
rect 110326 110599 110382 110608
rect 110326 107672 110382 107681
rect 109880 107630 110326 107658
rect 110326 107607 110382 107616
rect 109788 103486 110368 103514
rect 110340 98161 110368 103486
rect 110326 98152 110382 98161
rect 110326 98087 110382 98096
rect 109696 93826 110368 93854
rect 111076 93838 111104 142126
rect 111168 126954 111196 146118
rect 111260 143546 111288 150418
rect 111248 143540 111300 143546
rect 111248 143482 111300 143488
rect 111352 143426 111380 150583
rect 111260 143398 111380 143426
rect 111156 126948 111208 126954
rect 111156 126890 111208 126896
rect 111260 96626 111288 143398
rect 111444 143290 111472 150622
rect 111352 143262 111472 143290
rect 111352 137970 111380 143262
rect 111432 143200 111484 143206
rect 111432 143142 111484 143148
rect 111340 137964 111392 137970
rect 111340 137906 111392 137912
rect 111444 102134 111472 143142
rect 111536 140758 111564 150690
rect 111628 150074 111656 155858
rect 111708 155440 111760 155446
rect 111708 155382 111760 155388
rect 111720 151337 111748 155382
rect 111812 154970 111840 155858
rect 111800 154964 111852 154970
rect 111800 154906 111852 154912
rect 112088 153610 112116 159200
rect 112916 154737 112944 159200
rect 113180 154896 113232 154902
rect 113178 154864 113180 154873
rect 113232 154864 113234 154873
rect 113178 154799 113234 154808
rect 113456 154828 113508 154834
rect 113456 154770 113508 154776
rect 113468 154737 113496 154770
rect 112902 154728 112958 154737
rect 112902 154663 112958 154672
rect 113454 154728 113510 154737
rect 113454 154663 113510 154672
rect 113638 154728 113694 154737
rect 113638 154663 113694 154672
rect 113652 154630 113680 154663
rect 113744 154630 113772 159200
rect 114572 155038 114600 159200
rect 115400 155446 115428 159200
rect 116228 155446 116256 159200
rect 115388 155440 115440 155446
rect 115388 155382 115440 155388
rect 115848 155440 115900 155446
rect 115848 155382 115900 155388
rect 116216 155440 116268 155446
rect 116216 155382 116268 155388
rect 114560 155032 114612 155038
rect 114560 154974 114612 154980
rect 115756 155032 115808 155038
rect 115756 154974 115808 154980
rect 113640 154624 113692 154630
rect 113640 154566 113692 154572
rect 113732 154624 113784 154630
rect 113732 154566 113784 154572
rect 112076 153604 112128 153610
rect 112076 153546 112128 153552
rect 112442 151600 112498 151609
rect 112442 151535 112498 151544
rect 111706 151328 111762 151337
rect 111706 151263 111762 151272
rect 111706 151192 111762 151201
rect 111706 151127 111762 151136
rect 111616 150068 111668 150074
rect 111616 150010 111668 150016
rect 111720 142154 111748 151127
rect 111628 142126 111748 142154
rect 111524 140752 111576 140758
rect 111524 140694 111576 140700
rect 111628 104854 111656 142126
rect 112456 107642 112484 151535
rect 115768 150822 115796 154974
rect 115860 151201 115888 155382
rect 115940 155032 115992 155038
rect 115940 154974 115992 154980
rect 115952 154873 115980 154974
rect 117056 154902 117084 159200
rect 117884 155446 117912 159200
rect 117228 155440 117280 155446
rect 117228 155382 117280 155388
rect 117872 155440 117924 155446
rect 117872 155382 117924 155388
rect 118608 155440 118660 155446
rect 118608 155382 118660 155388
rect 117240 155038 117268 155382
rect 117136 155032 117188 155038
rect 117136 154974 117188 154980
rect 117228 155032 117280 155038
rect 117228 154974 117280 154980
rect 116584 154896 116636 154902
rect 115938 154864 115994 154873
rect 116584 154838 116636 154844
rect 117044 154896 117096 154902
rect 117044 154838 117096 154844
rect 115938 154799 115994 154808
rect 116492 152108 116544 152114
rect 116492 152050 116544 152056
rect 116214 152008 116270 152017
rect 116214 151943 116270 151952
rect 115846 151192 115902 151201
rect 115846 151127 115902 151136
rect 115756 150816 115808 150822
rect 115756 150758 115808 150764
rect 114100 150408 114152 150414
rect 114100 150350 114152 150356
rect 114008 150340 114060 150346
rect 114008 150282 114060 150288
rect 112902 149560 112958 149569
rect 112902 149495 112958 149504
rect 112718 149424 112774 149433
rect 112718 149359 112774 149368
rect 112534 149288 112590 149297
rect 112534 149223 112590 149232
rect 112548 121446 112576 149223
rect 112732 122806 112760 149359
rect 112916 124166 112944 149495
rect 113822 144256 113878 144265
rect 113822 144191 113878 144200
rect 112904 124160 112956 124166
rect 112904 124102 112956 124108
rect 112720 122800 112772 122806
rect 112720 122742 112772 122748
rect 112536 121440 112588 121446
rect 112536 121382 112588 121388
rect 112444 107636 112496 107642
rect 112444 107578 112496 107584
rect 111616 104848 111668 104854
rect 111616 104790 111668 104796
rect 111432 102128 111484 102134
rect 111432 102070 111484 102076
rect 111248 96620 111300 96626
rect 111248 96562 111300 96568
rect 110340 88369 110368 93826
rect 111064 93832 111116 93838
rect 111064 93774 111116 93780
rect 110326 88360 110382 88369
rect 113836 88330 113864 144191
rect 113914 132832 113970 132841
rect 113914 132767 113970 132776
rect 110326 88295 110382 88304
rect 113824 88324 113876 88330
rect 113824 88266 113876 88272
rect 113928 86970 113956 132767
rect 114020 131102 114048 150282
rect 114112 132190 114140 150350
rect 115204 150272 115256 150278
rect 115204 150214 115256 150220
rect 114100 132184 114152 132190
rect 114100 132126 114152 132132
rect 114008 131096 114060 131102
rect 114008 131038 114060 131044
rect 115216 127945 115244 150214
rect 116032 150204 116084 150210
rect 116032 150146 116084 150152
rect 116044 145217 116072 150146
rect 116124 149048 116176 149054
rect 116122 149016 116124 149025
rect 116176 149016 116178 149025
rect 116122 148951 116178 148960
rect 116030 145208 116086 145217
rect 116030 145143 116086 145152
rect 116124 143540 116176 143546
rect 116124 143482 116176 143488
rect 116136 143313 116164 143482
rect 116122 143304 116178 143313
rect 116122 143239 116178 143248
rect 116124 140752 116176 140758
rect 116124 140694 116176 140700
rect 116136 139505 116164 140694
rect 116122 139496 116178 139505
rect 116122 139431 116178 139440
rect 116124 137964 116176 137970
rect 116124 137906 116176 137912
rect 116136 137601 116164 137906
rect 116122 137592 116178 137601
rect 116122 137527 116178 137536
rect 115940 132184 115992 132190
rect 115940 132126 115992 132132
rect 115952 131753 115980 132126
rect 115938 131744 115994 131753
rect 115938 131679 115994 131688
rect 115940 131096 115992 131102
rect 115940 131038 115992 131044
rect 115952 129849 115980 131038
rect 115938 129840 115994 129849
rect 115938 129775 115994 129784
rect 115202 127936 115258 127945
rect 115202 127871 115258 127880
rect 116124 126948 116176 126954
rect 116124 126890 116176 126896
rect 116136 126041 116164 126890
rect 116122 126032 116178 126041
rect 116122 125967 116178 125976
rect 116124 124160 116176 124166
rect 116122 124128 116124 124137
rect 116176 124128 116178 124137
rect 116122 124063 116178 124072
rect 116124 122800 116176 122806
rect 116124 122742 116176 122748
rect 116136 122233 116164 122742
rect 116122 122224 116178 122233
rect 116122 122159 116178 122168
rect 116124 121440 116176 121446
rect 114006 121408 114062 121417
rect 116124 121382 116176 121388
rect 114006 121343 114062 121352
rect 113916 86964 113968 86970
rect 113916 86906 113968 86912
rect 114020 83978 114048 121343
rect 116136 120193 116164 121382
rect 116122 120184 116178 120193
rect 116122 120119 116178 120128
rect 114098 110120 114154 110129
rect 114098 110055 114154 110064
rect 114008 83972 114060 83978
rect 114008 83914 114060 83920
rect 114112 82822 114140 110055
rect 116124 107636 116176 107642
rect 116124 107578 116176 107584
rect 116136 106865 116164 107578
rect 116122 106856 116178 106865
rect 116122 106791 116178 106800
rect 116124 104848 116176 104854
rect 116122 104816 116124 104825
rect 116176 104816 116178 104825
rect 116122 104751 116178 104760
rect 115940 102128 115992 102134
rect 115940 102070 115992 102076
rect 115952 101017 115980 102070
rect 115938 101008 115994 101017
rect 115938 100943 115994 100952
rect 114190 98696 114246 98705
rect 114190 98631 114246 98640
rect 114100 82816 114152 82822
rect 114100 82758 114152 82764
rect 114204 80034 114232 98631
rect 116228 97209 116256 151943
rect 116398 149696 116454 149705
rect 116398 149631 116454 149640
rect 116412 142154 116440 149631
rect 116504 147121 116532 152050
rect 116596 151473 116624 154838
rect 116858 154728 116914 154737
rect 116768 154692 116820 154698
rect 116858 154663 116860 154672
rect 116768 154634 116820 154640
rect 116912 154663 116914 154672
rect 116860 154634 116912 154640
rect 116676 151972 116728 151978
rect 116676 151914 116728 151920
rect 116582 151464 116638 151473
rect 116582 151399 116638 151408
rect 116582 149152 116638 149161
rect 116582 149087 116638 149096
rect 116490 147112 116546 147121
rect 116490 147047 116546 147056
rect 116596 146826 116624 149087
rect 116688 147014 116716 151914
rect 116780 150686 116808 154634
rect 116860 150884 116912 150890
rect 116860 150826 116912 150832
rect 116768 150680 116820 150686
rect 116768 150622 116820 150628
rect 116676 147008 116728 147014
rect 116676 146950 116728 146956
rect 116596 146798 116716 146826
rect 116688 142154 116716 146798
rect 116412 142126 116624 142154
rect 116688 142126 116808 142154
rect 116214 97200 116270 97209
rect 116214 97135 116270 97144
rect 116124 96620 116176 96626
rect 116124 96562 116176 96568
rect 116136 95305 116164 96562
rect 116122 95296 116178 95305
rect 116122 95231 116178 95240
rect 116124 93832 116176 93838
rect 116124 93774 116176 93780
rect 116136 93401 116164 93774
rect 116122 93392 116178 93401
rect 116122 93327 116178 93336
rect 116596 91361 116624 142126
rect 116780 102921 116808 142126
rect 116872 112577 116900 150826
rect 116952 150544 117004 150550
rect 116952 150486 117004 150492
rect 116964 116385 116992 150486
rect 117148 150482 117176 154974
rect 118620 150822 118648 155382
rect 118804 153649 118832 159200
rect 118976 156664 119028 156670
rect 118976 156606 119028 156612
rect 118790 153640 118846 153649
rect 118790 153575 118846 153584
rect 118608 150816 118660 150822
rect 118608 150758 118660 150764
rect 117228 150612 117280 150618
rect 117228 150554 117280 150560
rect 117136 150476 117188 150482
rect 117136 150418 117188 150424
rect 117136 150136 117188 150142
rect 117136 150078 117188 150084
rect 117044 147008 117096 147014
rect 117044 146950 117096 146956
rect 117056 118289 117084 146950
rect 117148 133657 117176 150078
rect 117240 135561 117268 150554
rect 118988 149954 119016 156606
rect 119632 152114 119660 159200
rect 120460 155417 120488 159200
rect 121288 157334 121316 159200
rect 121288 157306 121408 157334
rect 121276 156188 121328 156194
rect 121276 156130 121328 156136
rect 120540 155440 120592 155446
rect 120446 155408 120502 155417
rect 120540 155382 120592 155388
rect 120446 155343 120502 155352
rect 120552 154834 120580 155382
rect 121090 155136 121146 155145
rect 121090 155071 121146 155080
rect 120632 155032 120684 155038
rect 120632 154974 120684 154980
rect 120644 154834 120672 154974
rect 120540 154828 120592 154834
rect 120540 154770 120592 154776
rect 120632 154828 120684 154834
rect 120632 154770 120684 154776
rect 119804 153876 119856 153882
rect 119804 153818 119856 153824
rect 119620 152108 119672 152114
rect 119620 152050 119672 152056
rect 119816 150090 119844 153818
rect 120446 153776 120502 153785
rect 120446 153711 120502 153720
rect 120460 150090 120488 153711
rect 121104 150090 121132 155071
rect 121288 154698 121316 156130
rect 121276 154692 121328 154698
rect 121276 154634 121328 154640
rect 121380 150754 121408 157306
rect 121736 156732 121788 156738
rect 121736 156674 121788 156680
rect 121368 150748 121420 150754
rect 121368 150690 121420 150696
rect 121748 150090 121776 156674
rect 122116 153882 122144 159200
rect 122748 156800 122800 156806
rect 122748 156742 122800 156748
rect 122760 155446 122788 156742
rect 122748 155440 122800 155446
rect 122748 155382 122800 155388
rect 122944 154698 122972 159200
rect 123484 155440 123536 155446
rect 123484 155382 123536 155388
rect 123392 155032 123444 155038
rect 123392 154974 123444 154980
rect 122932 154692 122984 154698
rect 122932 154634 122984 154640
rect 122380 153944 122432 153950
rect 122380 153886 122432 153892
rect 122104 153876 122156 153882
rect 122104 153818 122156 153824
rect 122392 150090 122420 153886
rect 123404 152046 123432 154974
rect 123496 154630 123524 155382
rect 123772 155038 123800 159200
rect 124312 156732 124364 156738
rect 124312 156674 124364 156680
rect 123760 155032 123812 155038
rect 123760 154974 123812 154980
rect 123484 154624 123536 154630
rect 123484 154566 123536 154572
rect 123666 152416 123722 152425
rect 123666 152351 123722 152360
rect 123392 152040 123444 152046
rect 123392 151982 123444 151988
rect 123024 151088 123076 151094
rect 123024 151030 123076 151036
rect 123036 150090 123064 151030
rect 123680 150090 123708 152351
rect 124324 150090 124352 156674
rect 124600 156670 124628 159200
rect 124588 156664 124640 156670
rect 124588 156606 124640 156612
rect 124954 156088 125010 156097
rect 124954 156023 125010 156032
rect 124968 150090 124996 156023
rect 125520 153882 125548 159200
rect 126242 155272 126298 155281
rect 126242 155207 126298 155216
rect 125508 153876 125560 153882
rect 125508 153818 125560 153824
rect 125692 153468 125744 153474
rect 125692 153410 125744 153416
rect 125598 152280 125654 152289
rect 125598 152215 125654 152224
rect 125612 150090 125640 152215
rect 125704 151978 125732 153410
rect 125692 151972 125744 151978
rect 125692 151914 125744 151920
rect 126256 150090 126284 155207
rect 126348 152289 126376 159200
rect 127176 154902 127204 159200
rect 127164 154896 127216 154902
rect 127164 154838 127216 154844
rect 126334 152280 126390 152289
rect 126334 152215 126390 152224
rect 126888 151904 126940 151910
rect 126888 151846 126940 151852
rect 126900 150090 126928 151846
rect 127532 151156 127584 151162
rect 127532 151098 127584 151104
rect 127544 150090 127572 151098
rect 128004 151094 128032 159200
rect 128268 155032 128320 155038
rect 128268 154974 128320 154980
rect 128176 152040 128228 152046
rect 128176 151982 128228 151988
rect 128280 151994 128308 154974
rect 128544 154964 128596 154970
rect 128544 154906 128596 154912
rect 128452 152040 128504 152046
rect 128280 151988 128452 151994
rect 128280 151982 128504 151988
rect 128188 151858 128216 151982
rect 128280 151966 128492 151982
rect 128556 151910 128584 154906
rect 128832 154698 128860 159200
rect 129660 154698 129688 159200
rect 130108 156868 130160 156874
rect 130108 156810 130160 156816
rect 128820 154692 128872 154698
rect 128820 154634 128872 154640
rect 129556 154692 129608 154698
rect 129556 154634 129608 154640
rect 129648 154692 129700 154698
rect 129648 154634 129700 154640
rect 129568 154086 129596 154634
rect 129464 154080 129516 154086
rect 129464 154022 129516 154028
rect 129556 154080 129608 154086
rect 129556 154022 129608 154028
rect 128820 152516 128872 152522
rect 128820 152458 128872 152464
rect 128544 151904 128596 151910
rect 128188 151842 128308 151858
rect 128544 151846 128596 151852
rect 128084 151836 128136 151842
rect 128188 151836 128320 151842
rect 128188 151830 128268 151836
rect 128084 151778 128136 151784
rect 128268 151778 128320 151784
rect 127992 151088 128044 151094
rect 127992 151030 128044 151036
rect 128096 150226 128124 151778
rect 128832 150226 128860 152458
rect 129476 150226 129504 154022
rect 130120 150226 130148 156810
rect 130488 155038 130516 159200
rect 131408 156738 131436 159200
rect 131396 156732 131448 156738
rect 131396 156674 131448 156680
rect 131118 155952 131174 155961
rect 131118 155887 131174 155896
rect 131026 155544 131082 155553
rect 131026 155479 131082 155488
rect 130476 155032 130528 155038
rect 130476 154974 130528 154980
rect 130750 153096 130806 153105
rect 130750 153031 130806 153040
rect 130764 150226 130792 153031
rect 131040 151814 131068 155479
rect 131132 153105 131160 155887
rect 132236 154018 132264 159200
rect 133064 155310 133092 159200
rect 132960 155304 133012 155310
rect 132958 155272 132960 155281
rect 133052 155304 133104 155310
rect 133012 155272 133014 155281
rect 133052 155246 133104 155252
rect 132958 155207 133014 155216
rect 133892 155038 133920 159200
rect 134522 155680 134578 155689
rect 134720 155650 134748 159200
rect 135352 156936 135404 156942
rect 135352 156878 135404 156884
rect 134522 155615 134578 155624
rect 134616 155644 134668 155650
rect 133236 155032 133288 155038
rect 133236 154974 133288 154980
rect 133880 155032 133932 155038
rect 133880 154974 133932 154980
rect 132040 154012 132092 154018
rect 132040 153954 132092 153960
rect 132224 154012 132276 154018
rect 132224 153954 132276 153960
rect 131118 153096 131174 153105
rect 131118 153031 131174 153040
rect 131040 151786 131436 151814
rect 131408 150226 131436 151786
rect 132052 150226 132080 153954
rect 133248 152561 133276 154974
rect 134536 152697 134564 155615
rect 134616 155586 134668 155592
rect 134708 155644 134760 155650
rect 134708 155586 134760 155592
rect 135168 155644 135220 155650
rect 135168 155586 135220 155592
rect 134628 154970 134656 155586
rect 134616 154964 134668 154970
rect 134616 154906 134668 154912
rect 134614 153912 134670 153921
rect 134614 153847 134670 153856
rect 133970 152688 134026 152697
rect 133970 152623 134026 152632
rect 134522 152688 134578 152697
rect 134522 152623 134578 152632
rect 133234 152552 133290 152561
rect 133234 152487 133290 152496
rect 133326 152416 133382 152425
rect 133326 152351 133382 152360
rect 132684 151224 132736 151230
rect 132684 151166 132736 151172
rect 128096 150198 128262 150226
rect 128832 150198 128906 150226
rect 129476 150198 129550 150226
rect 130120 150198 130194 150226
rect 130764 150198 130838 150226
rect 131408 150198 131482 150226
rect 132052 150198 132126 150226
rect 119816 150062 119890 150090
rect 120460 150062 120534 150090
rect 121104 150062 121178 150090
rect 121748 150062 121822 150090
rect 122392 150062 122466 150090
rect 123036 150062 123110 150090
rect 123680 150062 123754 150090
rect 124324 150062 124398 150090
rect 124968 150062 125042 150090
rect 125612 150062 125686 150090
rect 126256 150062 126330 150090
rect 126900 150062 126974 150090
rect 127544 150062 127618 150090
rect 118988 149926 119324 149954
rect 119862 149940 119890 150062
rect 120506 149940 120534 150062
rect 121150 149940 121178 150062
rect 121794 149940 121822 150062
rect 122438 149940 122466 150062
rect 123082 149940 123110 150062
rect 123726 149940 123754 150062
rect 124370 149940 124398 150062
rect 125014 149940 125042 150062
rect 125658 149940 125686 150062
rect 126302 149940 126330 150062
rect 126946 149940 126974 150062
rect 127590 149940 127618 150062
rect 128234 149940 128262 150198
rect 128878 149940 128906 150198
rect 129522 149940 129550 150198
rect 130166 149940 130194 150198
rect 130810 149940 130838 150198
rect 131454 149940 131482 150198
rect 132098 149940 132126 150198
rect 132696 150090 132724 151166
rect 133340 150226 133368 152351
rect 133984 150226 134012 152623
rect 134628 150226 134656 153847
rect 135180 151162 135208 155586
rect 135168 151156 135220 151162
rect 135168 151098 135220 151104
rect 135364 150226 135392 156878
rect 135548 153474 135576 159200
rect 136376 155650 136404 159200
rect 137100 157004 137152 157010
rect 137100 156946 137152 156952
rect 136364 155644 136416 155650
rect 136364 155586 136416 155592
rect 137008 155304 137060 155310
rect 137008 155246 137060 155252
rect 135904 155236 135956 155242
rect 135904 155178 135956 155184
rect 135536 153468 135588 153474
rect 135536 153410 135588 153416
rect 133340 150198 133414 150226
rect 133984 150198 134058 150226
rect 134628 150198 134702 150226
rect 132696 150062 132770 150090
rect 132742 149940 132770 150062
rect 133386 149940 133414 150198
rect 134030 149940 134058 150198
rect 134674 149940 134702 150198
rect 135318 150198 135392 150226
rect 135916 150226 135944 155178
rect 136916 154964 136968 154970
rect 136916 154906 136968 154912
rect 136928 154873 136956 154906
rect 136914 154864 136970 154873
rect 136914 154799 136970 154808
rect 136546 152688 136602 152697
rect 136546 152623 136602 152632
rect 136560 150226 136588 152623
rect 137020 152522 137048 155246
rect 137008 152516 137060 152522
rect 137008 152458 137060 152464
rect 137112 151814 137140 156946
rect 137204 155242 137232 159200
rect 138124 156942 138152 159200
rect 138112 156936 138164 156942
rect 138112 156878 138164 156884
rect 138018 155816 138074 155825
rect 138018 155751 138074 155760
rect 137376 155304 137428 155310
rect 137374 155272 137376 155281
rect 137428 155272 137430 155281
rect 137192 155236 137244 155242
rect 137374 155207 137430 155216
rect 137192 155178 137244 155184
rect 137652 155032 137704 155038
rect 137652 154974 137704 154980
rect 137376 154896 137428 154902
rect 137560 154896 137612 154902
rect 137376 154838 137428 154844
rect 137558 154864 137560 154873
rect 137612 154864 137614 154873
rect 137388 154714 137416 154838
rect 137558 154799 137614 154808
rect 137664 154714 137692 154974
rect 137388 154686 137692 154714
rect 138032 152522 138060 155751
rect 138952 153785 138980 159200
rect 138938 153776 138994 153785
rect 138938 153711 138994 153720
rect 139780 152726 139808 159200
rect 140412 157072 140464 157078
rect 140412 157014 140464 157020
rect 139124 152720 139176 152726
rect 139124 152662 139176 152668
rect 139768 152720 139820 152726
rect 139768 152662 139820 152668
rect 138480 152584 138532 152590
rect 138480 152526 138532 152532
rect 137284 152516 137336 152522
rect 137284 152458 137336 152464
rect 138020 152516 138072 152522
rect 138020 152458 138072 152464
rect 137112 151786 137232 151814
rect 137204 150226 137232 151786
rect 137296 151230 137324 152458
rect 137836 151292 137888 151298
rect 137836 151234 137888 151240
rect 137284 151224 137336 151230
rect 137284 151166 137336 151172
rect 135916 150198 135990 150226
rect 136560 150198 136634 150226
rect 137204 150198 137278 150226
rect 135318 149940 135346 150198
rect 135962 149940 135990 150198
rect 136606 149940 136634 150198
rect 137250 149940 137278 150198
rect 137848 150090 137876 151234
rect 138492 150226 138520 152526
rect 139136 150226 139164 152662
rect 139768 151972 139820 151978
rect 139768 151914 139820 151920
rect 139780 150226 139808 151914
rect 140424 150226 140452 157014
rect 140608 155281 140636 159200
rect 141436 156874 141464 159200
rect 141424 156868 141476 156874
rect 141424 156810 141476 156816
rect 142264 156754 142292 159200
rect 142712 158568 142764 158574
rect 142712 158510 142764 158516
rect 142264 156726 142476 156754
rect 140780 155304 140832 155310
rect 140594 155272 140650 155281
rect 140780 155246 140832 155252
rect 140594 155207 140650 155216
rect 140792 152590 140820 155246
rect 142448 154154 142476 156726
rect 142620 155236 142672 155242
rect 142620 155178 142672 155184
rect 142344 154148 142396 154154
rect 142344 154090 142396 154096
rect 142436 154148 142488 154154
rect 142436 154090 142488 154096
rect 141054 153096 141110 153105
rect 141054 153031 141110 153040
rect 140780 152584 140832 152590
rect 140780 152526 140832 152532
rect 141068 150226 141096 153031
rect 141792 152720 141844 152726
rect 141792 152662 141844 152668
rect 141804 152522 141832 152662
rect 141700 152516 141752 152522
rect 141700 152458 141752 152464
rect 141792 152516 141844 152522
rect 141792 152458 141844 152464
rect 141712 150226 141740 152458
rect 142356 150226 142384 154090
rect 142632 151978 142660 155178
rect 142620 151972 142672 151978
rect 142620 151914 142672 151920
rect 142724 151814 142752 158510
rect 143092 155310 143120 159200
rect 143448 157004 143500 157010
rect 143448 156946 143500 156952
rect 143460 156806 143488 156946
rect 143448 156800 143500 156806
rect 143448 156742 143500 156748
rect 143080 155304 143132 155310
rect 143080 155246 143132 155252
rect 143920 155242 143948 159200
rect 144840 157078 144868 159200
rect 144828 157072 144880 157078
rect 144828 157014 144880 157020
rect 145194 156632 145250 156641
rect 145194 156567 145250 156576
rect 143908 155236 143960 155242
rect 143908 155178 143960 155184
rect 144828 154896 144880 154902
rect 144828 154838 144880 154844
rect 144840 152794 144868 154838
rect 144276 152788 144328 152794
rect 144276 152730 144328 152736
rect 144828 152788 144880 152794
rect 144828 152730 144880 152736
rect 143632 152652 143684 152658
rect 143632 152594 143684 152600
rect 142724 151786 143028 151814
rect 143000 150226 143028 151786
rect 143644 150226 143672 152594
rect 144288 150226 144316 152730
rect 145208 151814 145236 156567
rect 145668 154290 145696 159200
rect 146208 157480 146260 157486
rect 146208 157422 146260 157428
rect 145564 154284 145616 154290
rect 145564 154226 145616 154232
rect 145656 154284 145708 154290
rect 145656 154226 145708 154232
rect 145024 151786 145236 151814
rect 145024 150226 145052 151786
rect 138492 150198 138566 150226
rect 139136 150198 139210 150226
rect 139780 150198 139854 150226
rect 140424 150198 140498 150226
rect 141068 150198 141142 150226
rect 141712 150198 141786 150226
rect 142356 150198 142430 150226
rect 143000 150198 143074 150226
rect 143644 150198 143718 150226
rect 144288 150198 144362 150226
rect 137848 150062 137922 150090
rect 137894 149940 137922 150062
rect 138538 149940 138566 150198
rect 139182 149940 139210 150198
rect 139826 149940 139854 150198
rect 140470 149940 140498 150198
rect 141114 149940 141142 150198
rect 141758 149940 141786 150198
rect 142402 149940 142430 150198
rect 143046 149940 143074 150198
rect 143690 149940 143718 150198
rect 144334 149940 144362 150198
rect 144978 150198 145052 150226
rect 145576 150226 145604 154226
rect 146220 150226 146248 157422
rect 146496 152658 146524 159200
rect 146852 157208 146904 157214
rect 146852 157150 146904 157156
rect 146484 152652 146536 152658
rect 146484 152594 146536 152600
rect 146760 152380 146812 152386
rect 146760 152322 146812 152328
rect 146772 150498 146800 152322
rect 146864 151814 146892 157150
rect 146944 155644 146996 155650
rect 146944 155586 146996 155592
rect 146956 154902 146984 155586
rect 147324 155553 147352 159200
rect 147680 157548 147732 157554
rect 147680 157490 147732 157496
rect 147310 155544 147366 155553
rect 147310 155479 147366 155488
rect 147588 155236 147640 155242
rect 147588 155178 147640 155184
rect 146944 154896 146996 154902
rect 146944 154838 146996 154844
rect 147600 152726 147628 155178
rect 147588 152720 147640 152726
rect 147588 152662 147640 152668
rect 146864 151786 147536 151814
rect 146772 150470 146892 150498
rect 146864 150226 146892 150470
rect 147508 150226 147536 151786
rect 145576 150198 145650 150226
rect 146220 150198 146294 150226
rect 146864 150198 146938 150226
rect 147508 150198 147582 150226
rect 147692 150210 147720 157490
rect 148152 157146 148180 159200
rect 148140 157140 148192 157146
rect 148140 157082 148192 157088
rect 148324 157072 148376 157078
rect 148152 157020 148324 157026
rect 148152 157014 148376 157020
rect 148152 157010 148364 157014
rect 148140 157004 148364 157010
rect 148192 156998 148364 157004
rect 148140 156946 148192 156952
rect 148980 154222 149008 159200
rect 149808 155242 149836 159200
rect 149980 157208 150032 157214
rect 149980 157150 150032 157156
rect 149796 155236 149848 155242
rect 149796 155178 149848 155184
rect 148140 154216 148192 154222
rect 148140 154158 148192 154164
rect 148968 154216 149020 154222
rect 148968 154158 149020 154164
rect 148152 150226 148180 154158
rect 149428 152584 149480 152590
rect 149428 152526 149480 152532
rect 149440 150226 149468 152526
rect 149992 150226 150020 157150
rect 150636 155258 150664 159200
rect 151268 157616 151320 157622
rect 151268 157558 151320 157564
rect 150636 155230 150756 155258
rect 150624 154352 150676 154358
rect 150624 154294 150676 154300
rect 150636 150226 150664 154294
rect 150728 152658 150756 155230
rect 150716 152652 150768 152658
rect 150716 152594 150768 152600
rect 151280 150226 151308 157558
rect 151556 157078 151584 159200
rect 151544 157072 151596 157078
rect 151544 157014 151596 157020
rect 152384 154358 152412 159200
rect 152556 157276 152608 157282
rect 152556 157218 152608 157224
rect 152372 154352 152424 154358
rect 152372 154294 152424 154300
rect 151912 152856 151964 152862
rect 151912 152798 151964 152804
rect 151924 150226 151952 152798
rect 152568 150226 152596 157218
rect 152924 157208 152976 157214
rect 152924 157150 152976 157156
rect 152936 156602 152964 157150
rect 152924 156596 152976 156602
rect 152924 156538 152976 156544
rect 153016 156596 153068 156602
rect 153016 156538 153068 156544
rect 152924 155780 152976 155786
rect 152924 155722 152976 155728
rect 152936 154714 152964 155722
rect 153028 154834 153056 156538
rect 153212 155632 153240 159200
rect 153752 157752 153804 157758
rect 153752 157694 153804 157700
rect 153660 155780 153712 155786
rect 153660 155722 153712 155728
rect 153292 155644 153344 155650
rect 153212 155604 153292 155632
rect 153292 155586 153344 155592
rect 153672 155582 153700 155722
rect 153660 155576 153712 155582
rect 153660 155518 153712 155524
rect 153016 154828 153068 154834
rect 153016 154770 153068 154776
rect 153108 154828 153160 154834
rect 153108 154770 153160 154776
rect 153120 154714 153148 154770
rect 152936 154686 153148 154714
rect 153198 154048 153254 154057
rect 153198 153983 153254 153992
rect 153212 150226 153240 153983
rect 153764 151814 153792 157694
rect 154040 155378 154068 159200
rect 154868 155582 154896 159200
rect 155132 157344 155184 157350
rect 155132 157286 155184 157292
rect 154856 155576 154908 155582
rect 154856 155518 154908 155524
rect 153936 155372 153988 155378
rect 153936 155314 153988 155320
rect 154028 155372 154080 155378
rect 154028 155314 154080 155320
rect 153948 152862 153976 155314
rect 154488 152924 154540 152930
rect 154488 152866 154540 152872
rect 153936 152856 153988 152862
rect 153936 152798 153988 152804
rect 153764 151786 153884 151814
rect 153856 150226 153884 151786
rect 154500 150226 154528 152866
rect 155144 150226 155172 157286
rect 155696 155666 155724 159200
rect 156328 157684 156380 157690
rect 156328 157626 156380 157632
rect 156052 157344 156104 157350
rect 156052 157286 156104 157292
rect 155868 157276 155920 157282
rect 155868 157218 155920 157224
rect 155696 155638 155816 155666
rect 155684 155576 155736 155582
rect 155684 155518 155736 155524
rect 155592 154420 155644 154426
rect 155592 154362 155644 154368
rect 155604 150498 155632 154362
rect 155696 151298 155724 155518
rect 155788 154426 155816 155638
rect 155880 154902 155908 157218
rect 156064 156534 156092 157286
rect 156052 156528 156104 156534
rect 156052 156470 156104 156476
rect 155868 154896 155920 154902
rect 155868 154838 155920 154844
rect 155776 154420 155828 154426
rect 155776 154362 155828 154368
rect 156340 151814 156368 157626
rect 156420 157004 156472 157010
rect 156420 156946 156472 156952
rect 156432 156534 156460 156946
rect 156420 156528 156472 156534
rect 156420 156470 156472 156476
rect 156524 155582 156552 159200
rect 156696 155780 156748 155786
rect 156696 155722 156748 155728
rect 156512 155576 156564 155582
rect 156512 155518 156564 155524
rect 156604 155236 156656 155242
rect 156604 155178 156656 155184
rect 156616 154834 156644 155178
rect 156604 154828 156656 154834
rect 156604 154770 156656 154776
rect 156708 152930 156736 155722
rect 156696 152924 156748 152930
rect 156696 152866 156748 152872
rect 157352 152794 157380 159200
rect 157708 157208 157760 157214
rect 157708 157150 157760 157156
rect 157064 152788 157116 152794
rect 157064 152730 157116 152736
rect 157340 152788 157392 152794
rect 157340 152730 157392 152736
rect 156340 151786 156460 151814
rect 155684 151292 155736 151298
rect 155684 151234 155736 151240
rect 155604 150470 155816 150498
rect 155788 150226 155816 150470
rect 156432 150226 156460 151786
rect 157076 150226 157104 152730
rect 144978 149940 145006 150198
rect 145622 149940 145650 150198
rect 146266 149940 146294 150198
rect 146910 149940 146938 150198
rect 147554 149940 147582 150198
rect 147680 150204 147732 150210
rect 148152 150198 148226 150226
rect 147680 150146 147732 150152
rect 148198 149940 148226 150198
rect 148830 150204 148882 150210
rect 149440 150198 149514 150226
rect 149992 150198 150066 150226
rect 150636 150198 150710 150226
rect 151280 150198 151354 150226
rect 151924 150198 151998 150226
rect 152568 150198 152642 150226
rect 153212 150198 153286 150226
rect 153856 150198 153930 150226
rect 154500 150198 154574 150226
rect 155144 150198 155218 150226
rect 155788 150198 155862 150226
rect 156432 150198 156506 150226
rect 157076 150198 157150 150226
rect 148830 150146 148882 150152
rect 148842 149940 148870 150146
rect 149486 149940 149514 150198
rect 150038 149940 150066 150198
rect 150682 149940 150710 150198
rect 151326 149940 151354 150198
rect 151970 149940 151998 150198
rect 152614 149940 152642 150198
rect 153258 149940 153286 150198
rect 153902 149940 153930 150198
rect 154546 149940 154574 150198
rect 155190 149940 155218 150198
rect 155834 149940 155862 150198
rect 156478 149940 156506 150198
rect 157122 149940 157150 150198
rect 157720 150090 157748 157150
rect 158272 157146 158300 159200
rect 158996 157820 159048 157826
rect 158996 157762 159048 157768
rect 158260 157140 158312 157146
rect 158260 157082 158312 157088
rect 158812 155780 158864 155786
rect 158812 155722 158864 155728
rect 158824 155582 158852 155722
rect 158812 155576 158864 155582
rect 158812 155518 158864 155524
rect 158352 154556 158404 154562
rect 158352 154498 158404 154504
rect 158364 150090 158392 154498
rect 159008 150226 159036 157762
rect 159100 154562 159128 159200
rect 159928 155582 159956 159200
rect 160284 157344 160336 157350
rect 160284 157286 160336 157292
rect 159916 155576 159968 155582
rect 159916 155518 159968 155524
rect 159088 154556 159140 154562
rect 159088 154498 159140 154504
rect 159640 152856 159692 152862
rect 159640 152798 159692 152804
rect 159008 150198 159082 150226
rect 157720 150062 157794 150090
rect 158364 150062 158438 150090
rect 157766 149940 157794 150062
rect 158410 149940 158438 150062
rect 159054 149940 159082 150198
rect 159652 150090 159680 152798
rect 160296 150090 160324 157286
rect 160756 155378 160784 159200
rect 161584 157214 161612 159200
rect 161664 157888 161716 157894
rect 161664 157830 161716 157836
rect 161572 157208 161624 157214
rect 161572 157150 161624 157156
rect 160652 155372 160704 155378
rect 160652 155314 160704 155320
rect 160744 155372 160796 155378
rect 160744 155314 160796 155320
rect 160664 155258 160692 155314
rect 160664 155242 160876 155258
rect 160664 155236 160888 155242
rect 160664 155230 160836 155236
rect 160836 155178 160888 155184
rect 161204 154896 161256 154902
rect 161204 154838 161256 154844
rect 161296 154896 161348 154902
rect 161296 154838 161348 154844
rect 160928 154488 160980 154494
rect 160928 154430 160980 154436
rect 160940 150090 160968 154430
rect 161216 152386 161244 154838
rect 161308 154766 161336 154838
rect 161296 154760 161348 154766
rect 161296 154702 161348 154708
rect 161204 152380 161256 152386
rect 161204 152322 161256 152328
rect 161676 150226 161704 157830
rect 161940 157344 161992 157350
rect 162412 157334 162440 159200
rect 161940 157286 161992 157292
rect 162044 157306 162440 157334
rect 161952 156466 161980 157286
rect 161940 156460 161992 156466
rect 161940 156402 161992 156408
rect 162044 154494 162072 157306
rect 162584 157276 162636 157282
rect 162584 157218 162636 157224
rect 162124 156528 162176 156534
rect 162124 156470 162176 156476
rect 162136 156346 162164 156470
rect 162596 156466 162624 157218
rect 162584 156460 162636 156466
rect 162584 156402 162636 156408
rect 162492 156392 162544 156398
rect 162136 156340 162492 156346
rect 162136 156334 162544 156340
rect 162136 156318 162532 156334
rect 162124 155508 162176 155514
rect 162124 155450 162176 155456
rect 162136 154766 162164 155450
rect 162124 154760 162176 154766
rect 162124 154702 162176 154708
rect 162032 154488 162084 154494
rect 162032 154430 162084 154436
rect 162216 152992 162268 152998
rect 162216 152934 162268 152940
rect 162858 152960 162914 152969
rect 161630 150198 161704 150226
rect 159652 150062 159726 150090
rect 160296 150062 160370 150090
rect 160940 150062 161014 150090
rect 159698 149940 159726 150062
rect 160342 149940 160370 150062
rect 160986 149940 161014 150062
rect 161630 149940 161658 150198
rect 162228 150090 162256 152934
rect 162858 152895 162914 152904
rect 162872 150090 162900 152895
rect 163240 152862 163268 159200
rect 163872 157956 163924 157962
rect 163872 157898 163924 157904
rect 163884 157334 163912 157898
rect 163884 157306 164096 157334
rect 163504 153808 163556 153814
rect 163504 153750 163556 153756
rect 163228 152856 163280 152862
rect 163228 152798 163280 152804
rect 163516 150090 163544 153750
rect 164068 150226 164096 157306
rect 164160 155514 164188 159200
rect 164240 155712 164292 155718
rect 164292 155660 164464 155666
rect 164240 155654 164464 155660
rect 164252 155638 164464 155654
rect 164436 155582 164464 155638
rect 164332 155576 164384 155582
rect 164332 155518 164384 155524
rect 164424 155576 164476 155582
rect 164424 155518 164476 155524
rect 164148 155508 164200 155514
rect 164148 155450 164200 155456
rect 164344 154902 164372 155518
rect 164240 154896 164292 154902
rect 164240 154838 164292 154844
rect 164332 154896 164384 154902
rect 164332 154838 164384 154844
rect 164252 153921 164280 154838
rect 164238 153912 164294 153921
rect 164238 153847 164294 153856
rect 164792 152924 164844 152930
rect 164792 152866 164844 152872
rect 164068 150198 164234 150226
rect 162228 150062 162302 150090
rect 162872 150062 162946 150090
rect 163516 150062 163590 150090
rect 162274 149940 162302 150062
rect 162918 149940 162946 150062
rect 163562 149940 163590 150062
rect 164206 149940 164234 150198
rect 164804 150090 164832 152866
rect 164988 150618 165016 159200
rect 165436 157344 165488 157350
rect 165436 157286 165488 157292
rect 164976 150612 165028 150618
rect 164976 150554 165028 150560
rect 165448 150090 165476 157286
rect 165620 155508 165672 155514
rect 165620 155450 165672 155456
rect 165632 152930 165660 155450
rect 165816 153814 165844 159200
rect 165988 158024 166040 158030
rect 165988 157966 166040 157972
rect 166000 157334 166028 157966
rect 166000 157306 166580 157334
rect 166078 154184 166134 154193
rect 166078 154119 166134 154128
rect 165804 153808 165856 153814
rect 165804 153750 165856 153756
rect 165620 152924 165672 152930
rect 165620 152866 165672 152872
rect 166092 150090 166120 154119
rect 166552 150226 166580 157306
rect 166644 155514 166672 159200
rect 167472 155718 167500 159200
rect 167460 155712 167512 155718
rect 167460 155654 167512 155660
rect 166632 155508 166684 155514
rect 166632 155450 166684 155456
rect 167644 154760 167696 154766
rect 167644 154702 167696 154708
rect 167368 153060 167420 153066
rect 167368 153002 167420 153008
rect 167380 150226 167408 153002
rect 167656 151842 167684 154702
rect 167552 151836 167604 151842
rect 167552 151778 167604 151784
rect 167644 151836 167696 151842
rect 167644 151778 167696 151784
rect 167564 150498 167592 151778
rect 168300 150686 168328 159200
rect 169128 153678 169156 159200
rect 169300 158092 169352 158098
rect 169300 158034 169352 158040
rect 168656 153672 168708 153678
rect 168656 153614 168708 153620
rect 169116 153672 169168 153678
rect 169116 153614 169168 153620
rect 168288 150680 168340 150686
rect 168288 150622 168340 150628
rect 167564 150470 168052 150498
rect 168024 150226 168052 150470
rect 168668 150226 168696 153614
rect 169312 150226 169340 158034
rect 169760 155576 169812 155582
rect 169760 155518 169812 155524
rect 169772 153066 169800 155518
rect 169760 153060 169812 153066
rect 169760 153002 169812 153008
rect 169956 152998 169984 159200
rect 170876 155582 170904 159200
rect 171704 157282 171732 159200
rect 171876 158228 171928 158234
rect 171876 158170 171928 158176
rect 171692 157276 171744 157282
rect 171692 157218 171744 157224
rect 171060 155774 171180 155802
rect 171060 155718 171088 155774
rect 171152 155718 171180 155774
rect 171048 155712 171100 155718
rect 171048 155654 171100 155660
rect 171140 155712 171192 155718
rect 171140 155654 171192 155660
rect 170864 155576 170916 155582
rect 170864 155518 170916 155524
rect 171232 153740 171284 153746
rect 171232 153682 171284 153688
rect 169944 152992 169996 152998
rect 169944 152934 169996 152940
rect 169944 152380 169996 152386
rect 169944 152322 169996 152328
rect 169956 150226 169984 152322
rect 170586 151056 170642 151065
rect 170586 150991 170642 151000
rect 166552 150198 166810 150226
rect 167380 150198 167454 150226
rect 168024 150198 168098 150226
rect 168668 150198 168742 150226
rect 169312 150198 169386 150226
rect 169956 150198 170030 150226
rect 164804 150062 164878 150090
rect 165448 150062 165522 150090
rect 166092 150062 166166 150090
rect 164850 149940 164878 150062
rect 165494 149940 165522 150062
rect 166138 149940 166166 150062
rect 166782 149940 166810 150198
rect 167426 149940 167454 150198
rect 168070 149940 168098 150198
rect 168714 149940 168742 150198
rect 169358 149940 169386 150198
rect 170002 149940 170030 150198
rect 170600 150090 170628 150991
rect 171244 150226 171272 153682
rect 171888 150226 171916 158170
rect 172532 157350 172560 159200
rect 172520 157344 172572 157350
rect 172520 157286 172572 157292
rect 173072 156528 173124 156534
rect 173072 156470 173124 156476
rect 172520 151836 172572 151842
rect 173084 151814 173112 156470
rect 173360 155582 173388 159200
rect 173440 155848 173492 155854
rect 173438 155816 173440 155825
rect 173492 155816 173494 155825
rect 174188 155786 174216 159200
rect 174452 158160 174504 158166
rect 174452 158102 174504 158108
rect 173438 155751 173494 155760
rect 174176 155780 174228 155786
rect 174176 155722 174228 155728
rect 173256 155576 173308 155582
rect 173256 155518 173308 155524
rect 173348 155576 173400 155582
rect 173348 155518 173400 155524
rect 173268 152386 173296 155518
rect 173256 152380 173308 152386
rect 173256 152322 173308 152328
rect 173084 151786 173204 151814
rect 172520 151778 172572 151784
rect 172532 150226 172560 151778
rect 173176 150226 173204 151786
rect 173808 151360 173860 151366
rect 173808 151302 173860 151308
rect 171244 150198 171318 150226
rect 171888 150198 171962 150226
rect 172532 150198 172606 150226
rect 173176 150198 173250 150226
rect 170600 150062 170674 150090
rect 170646 149940 170674 150062
rect 171290 149940 171318 150198
rect 171934 149940 171962 150198
rect 172578 149940 172606 150198
rect 173222 149940 173250 150198
rect 173820 150090 173848 151302
rect 174464 150226 174492 158102
rect 174544 156528 174596 156534
rect 174544 156470 174596 156476
rect 174556 155990 174584 156470
rect 174544 155984 174596 155990
rect 174544 155926 174596 155932
rect 175016 155564 175044 159200
rect 175844 156482 175872 159200
rect 175752 156454 175872 156482
rect 175936 156590 176332 156618
rect 175648 155848 175700 155854
rect 175648 155790 175700 155796
rect 175016 155536 175228 155564
rect 175096 153128 175148 153134
rect 175096 153070 175148 153076
rect 175108 150226 175136 153070
rect 175200 151366 175228 155536
rect 175660 151434 175688 155790
rect 175752 153746 175780 156454
rect 175832 156392 175884 156398
rect 175832 156334 175884 156340
rect 175844 155990 175872 156334
rect 175936 156330 175964 156590
rect 176304 156466 176332 156590
rect 176200 156460 176252 156466
rect 176200 156402 176252 156408
rect 176292 156460 176344 156466
rect 176292 156402 176344 156408
rect 175924 156324 175976 156330
rect 175924 156266 175976 156272
rect 176212 156262 176240 156402
rect 176200 156256 176252 156262
rect 176200 156198 176252 156204
rect 175832 155984 175884 155990
rect 175832 155926 175884 155932
rect 175832 155848 175884 155854
rect 175830 155816 175832 155825
rect 175884 155816 175886 155825
rect 175830 155751 175886 155760
rect 176016 155712 176068 155718
rect 176016 155654 176068 155660
rect 176028 155378 176056 155654
rect 175924 155372 175976 155378
rect 175924 155314 175976 155320
rect 176016 155372 176068 155378
rect 176016 155314 176068 155320
rect 175936 155174 175964 155314
rect 175832 155168 175884 155174
rect 175832 155110 175884 155116
rect 175924 155168 175976 155174
rect 175924 155110 175976 155116
rect 175844 154766 175872 155110
rect 175832 154760 175884 154766
rect 175832 154702 175884 154708
rect 175740 153740 175792 153746
rect 175740 153682 175792 153688
rect 176384 153536 176436 153542
rect 176384 153478 176436 153484
rect 175556 151428 175608 151434
rect 175556 151370 175608 151376
rect 175648 151428 175700 151434
rect 175648 151370 175700 151376
rect 175188 151360 175240 151366
rect 175188 151302 175240 151308
rect 175568 150226 175596 151370
rect 176396 150226 176424 153478
rect 176672 153134 176700 159200
rect 177028 158296 177080 158302
rect 177028 158238 177080 158244
rect 176660 153128 176712 153134
rect 176660 153070 176712 153076
rect 177040 150226 177068 158238
rect 177592 155786 177620 159200
rect 178040 156528 178092 156534
rect 178040 156470 178092 156476
rect 177764 155848 177816 155854
rect 177764 155790 177816 155796
rect 177580 155780 177632 155786
rect 177580 155722 177632 155728
rect 177776 153066 177804 155790
rect 177672 153060 177724 153066
rect 177672 153002 177724 153008
rect 177764 153060 177816 153066
rect 177764 153002 177816 153008
rect 177684 150226 177712 153002
rect 178052 151814 178080 156470
rect 178420 156330 178448 159200
rect 179248 156534 179276 159200
rect 179236 156528 179288 156534
rect 179236 156470 179288 156476
rect 178960 156460 179012 156466
rect 178960 156402 179012 156408
rect 178408 156324 178460 156330
rect 178408 156266 178460 156272
rect 178052 151786 178356 151814
rect 178328 150226 178356 151786
rect 178972 150226 179000 156402
rect 180076 155854 180104 159200
rect 180064 155848 180116 155854
rect 180064 155790 180116 155796
rect 180904 155582 180932 159200
rect 181732 159174 181852 159200
rect 181168 156392 181220 156398
rect 181168 156334 181220 156340
rect 180064 155576 180116 155582
rect 180064 155518 180116 155524
rect 180892 155576 180944 155582
rect 180892 155518 180944 155524
rect 180076 150482 180104 155518
rect 180248 153196 180300 153202
rect 180248 153138 180300 153144
rect 179604 150476 179656 150482
rect 179604 150418 179656 150424
rect 180064 150476 180116 150482
rect 180064 150418 180116 150424
rect 174464 150198 174538 150226
rect 175108 150198 175182 150226
rect 175568 150198 175826 150226
rect 176396 150198 176470 150226
rect 177040 150198 177114 150226
rect 177684 150198 177758 150226
rect 178328 150198 178402 150226
rect 178972 150198 179046 150226
rect 173820 150062 173894 150090
rect 173866 149940 173894 150062
rect 174510 149940 174538 150198
rect 175154 149940 175182 150198
rect 175798 149940 175826 150198
rect 176442 149940 176470 150198
rect 177086 149940 177114 150198
rect 177730 149940 177758 150198
rect 178374 149940 178402 150198
rect 179018 149940 179046 150198
rect 179616 150090 179644 150418
rect 180260 150226 180288 153138
rect 181180 151814 181208 156334
rect 180904 151786 181208 151814
rect 180904 150226 180932 151786
rect 182008 151502 182036 159310
rect 182546 159200 182602 160400
rect 183374 159200 183430 160400
rect 184294 159200 184350 160400
rect 185122 159200 185178 160400
rect 185950 159202 186006 160400
rect 186056 159310 186268 159338
rect 186056 159202 186084 159310
rect 185950 159200 186084 159202
rect 182088 158364 182140 158370
rect 182088 158306 182140 158312
rect 181444 151496 181496 151502
rect 181444 151438 181496 151444
rect 181996 151496 182048 151502
rect 181996 151438 182048 151444
rect 180260 150198 180334 150226
rect 179616 150062 179690 150090
rect 179662 149940 179690 150062
rect 180306 149940 180334 150198
rect 180858 150198 180932 150226
rect 180858 149940 180886 150198
rect 181456 150090 181484 151438
rect 182100 150226 182128 158306
rect 182560 153542 182588 159200
rect 183388 156466 183416 159200
rect 183376 156460 183428 156466
rect 183376 156402 183428 156408
rect 184308 155106 184336 159200
rect 185136 156398 185164 159200
rect 185964 159174 186084 159200
rect 185124 156392 185176 156398
rect 185124 156334 185176 156340
rect 185320 156330 185808 156346
rect 185320 156324 185820 156330
rect 185320 156318 185768 156324
rect 185320 156194 185348 156318
rect 185768 156266 185820 156272
rect 185676 156256 185728 156262
rect 185676 156198 185728 156204
rect 185308 156188 185360 156194
rect 185308 156130 185360 156136
rect 185400 156120 185452 156126
rect 185400 156062 185452 156068
rect 184204 155100 184256 155106
rect 184204 155042 184256 155048
rect 184296 155100 184348 155106
rect 184296 155042 184348 155048
rect 184216 154766 184244 155042
rect 183284 154760 183336 154766
rect 183284 154702 183336 154708
rect 184204 154760 184256 154766
rect 184204 154702 184256 154708
rect 182548 153536 182600 153542
rect 182548 153478 182600 153484
rect 183296 153202 183324 154702
rect 184952 154698 185164 154714
rect 184940 154692 185176 154698
rect 184992 154686 185124 154692
rect 184940 154634 184992 154640
rect 185124 154634 185176 154640
rect 184848 154624 184900 154630
rect 184848 154566 184900 154572
rect 184860 153406 184888 154566
rect 184020 153400 184072 153406
rect 184020 153342 184072 153348
rect 184848 153400 184900 153406
rect 184848 153342 184900 153348
rect 183284 153196 183336 153202
rect 183284 153138 183336 153144
rect 182732 153060 182784 153066
rect 182732 153002 182784 153008
rect 182744 150226 182772 153002
rect 183376 151632 183428 151638
rect 183376 151574 183428 151580
rect 182100 150198 182174 150226
rect 182744 150198 182818 150226
rect 181456 150062 181530 150090
rect 181502 149940 181530 150062
rect 182146 149940 182174 150198
rect 182790 149940 182818 150198
rect 183388 150090 183416 151574
rect 184032 150226 184060 153342
rect 185308 152448 185360 152454
rect 185308 152390 185360 152396
rect 184662 151464 184718 151473
rect 184662 151399 184718 151408
rect 184032 150198 184106 150226
rect 183388 150062 183462 150090
rect 183434 149940 183462 150062
rect 184078 149940 184106 150198
rect 184676 150090 184704 151399
rect 185320 150226 185348 152390
rect 185412 151814 185440 156062
rect 185688 156058 185716 156198
rect 185676 156052 185728 156058
rect 185676 155994 185728 156000
rect 185492 155848 185544 155854
rect 185492 155790 185544 155796
rect 185504 154766 185532 155790
rect 185676 155780 185728 155786
rect 185676 155722 185728 155728
rect 185688 155582 185716 155722
rect 185676 155576 185728 155582
rect 185676 155518 185728 155524
rect 186136 155100 186188 155106
rect 186136 155042 186188 155048
rect 185492 154760 185544 154766
rect 185492 154702 185544 154708
rect 186148 153134 186176 155042
rect 186136 153128 186188 153134
rect 186136 153070 186188 153076
rect 185412 151786 185992 151814
rect 185964 150226 185992 151786
rect 186240 151638 186268 159310
rect 186778 159200 186834 160400
rect 187606 159200 187662 160400
rect 188434 159200 188490 160400
rect 189262 159200 189318 160400
rect 190090 159200 190146 160400
rect 191010 159200 191066 160400
rect 191838 159200 191894 160400
rect 192666 159200 192722 160400
rect 193494 159200 193550 160400
rect 194322 159200 194378 160400
rect 195150 159200 195206 160400
rect 195978 159200 196034 160400
rect 196898 159200 196954 160400
rect 197726 159200 197782 160400
rect 198554 159200 198610 160400
rect 199382 159200 199438 160400
rect 200210 159200 200266 160400
rect 201038 159200 201094 160400
rect 201866 159200 201922 160400
rect 202694 159200 202750 160400
rect 203614 159200 203670 160400
rect 204442 159200 204498 160400
rect 205270 159200 205326 160400
rect 206098 159200 206154 160400
rect 206926 159200 206982 160400
rect 207754 159200 207810 160400
rect 208582 159200 208638 160400
rect 209410 159200 209466 160400
rect 210330 159200 210386 160400
rect 211158 159200 211214 160400
rect 211986 159200 212042 160400
rect 212814 159200 212870 160400
rect 213642 159200 213698 160400
rect 214470 159200 214526 160400
rect 215298 159200 215354 160400
rect 216126 159200 216182 160400
rect 217046 159200 217102 160400
rect 217874 159200 217930 160400
rect 218702 159200 218758 160400
rect 219530 159200 219586 160400
rect 220358 159202 220414 160400
rect 220464 159310 220768 159338
rect 220464 159202 220492 159310
rect 220358 159200 220492 159202
rect 186688 158432 186740 158438
rect 186688 158374 186740 158380
rect 186596 153332 186648 153338
rect 186596 153274 186648 153280
rect 186228 151632 186280 151638
rect 186228 151574 186280 151580
rect 185320 150198 185394 150226
rect 185964 150198 186038 150226
rect 184676 150062 184750 150090
rect 184722 149940 184750 150062
rect 185366 149940 185394 150198
rect 186010 149940 186038 150198
rect 186608 150090 186636 153274
rect 186700 150634 186728 158374
rect 186792 155514 186820 159200
rect 187620 155854 187648 159200
rect 188448 157334 188476 159200
rect 188448 157306 188660 157334
rect 187516 155848 187568 155854
rect 187516 155790 187568 155796
rect 187608 155848 187660 155854
rect 187608 155790 187660 155796
rect 186780 155508 186832 155514
rect 186780 155450 186832 155456
rect 187528 155106 187556 155790
rect 187516 155100 187568 155106
rect 187516 155042 187568 155048
rect 187884 153196 187936 153202
rect 187884 153138 187936 153144
rect 186700 150606 187280 150634
rect 187252 150226 187280 150606
rect 187252 150198 187326 150226
rect 186608 150062 186682 150090
rect 186654 149940 186682 150062
rect 187298 149940 187326 150198
rect 187896 150090 187924 153138
rect 188632 151570 188660 157306
rect 189170 156768 189226 156777
rect 189170 156703 189226 156712
rect 188988 154624 189040 154630
rect 188988 154566 189040 154572
rect 189000 152454 189028 154566
rect 188988 152448 189040 152454
rect 188988 152390 189040 152396
rect 188528 151564 188580 151570
rect 188528 151506 188580 151512
rect 188620 151564 188672 151570
rect 188620 151506 188672 151512
rect 188540 150090 188568 151506
rect 189184 150090 189212 156703
rect 189276 153406 189304 159200
rect 189816 156324 189868 156330
rect 189816 156266 189868 156272
rect 189264 153400 189316 153406
rect 189264 153342 189316 153348
rect 189828 150090 189856 156266
rect 190104 153202 190132 159200
rect 191024 157334 191052 159200
rect 190932 157306 191052 157334
rect 191852 157334 191880 159200
rect 192392 158500 192444 158506
rect 192392 158442 192444 158448
rect 191852 157306 191972 157334
rect 190828 155100 190880 155106
rect 190828 155042 190880 155048
rect 190840 154737 190868 155042
rect 190826 154728 190882 154737
rect 190826 154663 190882 154672
rect 190932 154630 190960 157306
rect 191288 156256 191340 156262
rect 191288 156198 191340 156204
rect 191104 155780 191156 155786
rect 191104 155722 191156 155728
rect 191116 155514 191144 155722
rect 191012 155508 191064 155514
rect 191012 155450 191064 155456
rect 191104 155508 191156 155514
rect 191104 155450 191156 155456
rect 191024 155394 191052 155450
rect 191024 155366 191236 155394
rect 191012 155304 191064 155310
rect 191012 155246 191064 155252
rect 191104 155304 191156 155310
rect 191104 155246 191156 155252
rect 191024 155106 191052 155246
rect 191116 155174 191144 155246
rect 191208 155174 191236 155366
rect 191104 155168 191156 155174
rect 191104 155110 191156 155116
rect 191196 155168 191248 155174
rect 191196 155110 191248 155116
rect 191012 155100 191064 155106
rect 191012 155042 191064 155048
rect 190920 154624 190972 154630
rect 190920 154566 190972 154572
rect 190092 153196 190144 153202
rect 190092 153138 190144 153144
rect 190458 152824 190514 152833
rect 190458 152759 190514 152768
rect 190472 150090 190500 152759
rect 190736 151768 190788 151774
rect 190920 151768 190972 151774
rect 190788 151716 190920 151722
rect 190736 151710 190972 151716
rect 190748 151694 190960 151710
rect 191012 151700 191064 151706
rect 191012 151642 191064 151648
rect 191024 151434 191052 151642
rect 191104 151632 191156 151638
rect 191104 151574 191156 151580
rect 191116 151434 191144 151574
rect 191012 151428 191064 151434
rect 191012 151370 191064 151376
rect 191104 151428 191156 151434
rect 191104 151370 191156 151376
rect 191300 150226 191328 156198
rect 191840 154624 191892 154630
rect 191840 154566 191892 154572
rect 191852 152697 191880 154566
rect 191838 152688 191894 152697
rect 191838 152623 191894 152632
rect 191748 151768 191800 151774
rect 191748 151710 191800 151716
rect 191162 150198 191328 150226
rect 187896 150062 187970 150090
rect 188540 150062 188614 150090
rect 189184 150062 189258 150090
rect 189828 150062 189902 150090
rect 190472 150062 190546 150090
rect 187942 149940 187970 150062
rect 188586 149940 188614 150062
rect 189230 149940 189258 150062
rect 189874 149940 189902 150062
rect 190518 149940 190546 150062
rect 191162 149940 191190 150198
rect 191760 150090 191788 151710
rect 191944 151638 191972 157306
rect 192022 154728 192078 154737
rect 192022 154663 192078 154672
rect 192036 154630 192064 154663
rect 192024 154624 192076 154630
rect 192024 154566 192076 154572
rect 191932 151632 191984 151638
rect 191932 151574 191984 151580
rect 192404 150226 192432 158442
rect 192680 156262 192708 159200
rect 192668 156256 192720 156262
rect 192668 156198 192720 156204
rect 193508 154698 193536 159200
rect 194336 155854 194364 159200
rect 195164 156330 195192 159200
rect 195992 157334 196020 159200
rect 195992 157306 196112 157334
rect 195152 156324 195204 156330
rect 195152 156266 195204 156272
rect 195704 155916 195756 155922
rect 195704 155858 195756 155864
rect 194324 155848 194376 155854
rect 194324 155790 194376 155796
rect 195716 155530 195744 155858
rect 195716 155502 196020 155530
rect 193220 154692 193272 154698
rect 193220 154634 193272 154640
rect 193496 154692 193548 154698
rect 193496 154634 193548 154640
rect 193232 154329 193260 154634
rect 194600 154624 194652 154630
rect 194600 154566 194652 154572
rect 193218 154320 193274 154329
rect 193218 154255 193274 154264
rect 194322 154184 194378 154193
rect 194322 154119 194378 154128
rect 193036 152448 193088 152454
rect 193036 152390 193088 152396
rect 192404 150198 192478 150226
rect 191760 150062 191834 150090
rect 191806 149940 191834 150062
rect 192450 149940 192478 150198
rect 193048 150090 193076 152390
rect 193680 151768 193732 151774
rect 193680 151710 193732 151716
rect 193692 150090 193720 151710
rect 194336 150090 194364 154119
rect 194612 151842 194640 154566
rect 195992 152454 196020 155502
rect 195980 152448 196032 152454
rect 195980 152390 196032 152396
rect 195612 152312 195664 152318
rect 195612 152254 195664 152260
rect 194600 151836 194652 151842
rect 194600 151778 194652 151784
rect 195060 151700 195112 151706
rect 195060 151642 195112 151648
rect 195072 150550 195100 151642
rect 194968 150544 195020 150550
rect 194968 150486 195020 150492
rect 195060 150544 195112 150550
rect 195060 150486 195112 150492
rect 194980 150090 195008 150486
rect 195624 150090 195652 152254
rect 196084 151706 196112 157306
rect 196806 156904 196862 156913
rect 196806 156839 196862 156848
rect 196072 151700 196124 151706
rect 196072 151642 196124 151648
rect 196256 151020 196308 151026
rect 196256 150962 196308 150968
rect 196268 150090 196296 150962
rect 196820 150226 196848 156839
rect 196912 155718 196940 159200
rect 197544 157412 197596 157418
rect 197544 157354 197596 157360
rect 196900 155712 196952 155718
rect 196900 155654 196952 155660
rect 197556 150226 197584 157354
rect 197740 154630 197768 159200
rect 197728 154624 197780 154630
rect 197728 154566 197780 154572
rect 198188 152448 198240 152454
rect 198188 152390 198240 152396
rect 196820 150198 196986 150226
rect 197556 150198 197630 150226
rect 193048 150062 193122 150090
rect 193692 150062 193766 150090
rect 194336 150062 194410 150090
rect 194980 150062 195054 150090
rect 195624 150062 195698 150090
rect 196268 150062 196342 150090
rect 193094 149940 193122 150062
rect 193738 149940 193766 150062
rect 194382 149940 194410 150062
rect 195026 149940 195054 150062
rect 195670 149940 195698 150062
rect 196314 149940 196342 150062
rect 196958 149940 196986 150198
rect 197602 149940 197630 150198
rect 198200 150090 198228 152390
rect 198568 151638 198596 159200
rect 198830 157040 198886 157049
rect 198830 156975 198886 156984
rect 198556 151632 198608 151638
rect 198556 151574 198608 151580
rect 198844 150090 198872 156975
rect 199396 151026 199424 159200
rect 200224 157334 200252 159200
rect 200224 157306 200896 157334
rect 200672 155916 200724 155922
rect 200672 155858 200724 155864
rect 200764 155916 200816 155922
rect 200764 155858 200816 155864
rect 200304 155848 200356 155854
rect 200304 155790 200356 155796
rect 200316 155718 200344 155790
rect 200396 155780 200448 155786
rect 200580 155780 200632 155786
rect 200448 155740 200580 155768
rect 200396 155722 200448 155728
rect 200580 155722 200632 155728
rect 200212 155712 200264 155718
rect 200212 155654 200264 155660
rect 200304 155712 200356 155718
rect 200304 155654 200356 155660
rect 200118 153912 200174 153921
rect 200118 153847 200174 153856
rect 199476 153264 199528 153270
rect 199476 153206 199528 153212
rect 199384 151020 199436 151026
rect 199384 150962 199436 150968
rect 199488 150090 199516 153206
rect 200132 150090 200160 153847
rect 200224 152833 200252 155654
rect 200684 155258 200712 155858
rect 200776 155446 200804 155858
rect 200868 155446 200896 157306
rect 201052 155854 201080 159200
rect 201040 155848 201092 155854
rect 201040 155790 201092 155796
rect 200764 155440 200816 155446
rect 200764 155382 200816 155388
rect 200856 155440 200908 155446
rect 200856 155382 200908 155388
rect 200684 155230 200988 155258
rect 200488 155100 200540 155106
rect 200488 155042 200540 155048
rect 200764 155100 200816 155106
rect 200764 155042 200816 155048
rect 200500 153270 200528 155042
rect 200776 154698 200804 155042
rect 200960 154698 200988 155230
rect 200764 154692 200816 154698
rect 200764 154634 200816 154640
rect 200948 154692 201000 154698
rect 200948 154634 201000 154640
rect 201880 153921 201908 159200
rect 202050 154456 202106 154465
rect 202050 154391 202106 154400
rect 201866 153912 201922 153921
rect 201866 153847 201922 153856
rect 200488 153264 200540 153270
rect 200488 153206 200540 153212
rect 200210 152824 200266 152833
rect 200210 152759 200266 152768
rect 200764 152244 200816 152250
rect 200764 152186 200816 152192
rect 200776 150090 200804 152186
rect 201408 150952 201460 150958
rect 201408 150894 201460 150900
rect 201420 150090 201448 150894
rect 202064 150090 202092 154391
rect 202708 150958 202736 159200
rect 203628 152454 203656 159200
rect 203616 152448 203668 152454
rect 203616 152390 203668 152396
rect 204456 152318 204484 159200
rect 205180 155984 205232 155990
rect 205180 155926 205232 155932
rect 204628 153604 204680 153610
rect 204628 153546 204680 153552
rect 204444 152312 204496 152318
rect 204444 152254 204496 152260
rect 203340 152176 203392 152182
rect 203340 152118 203392 152124
rect 202696 150952 202748 150958
rect 202696 150894 202748 150900
rect 202742 150136 202794 150142
rect 198200 150062 198274 150090
rect 198844 150062 198918 150090
rect 199488 150062 199562 150090
rect 200132 150062 200206 150090
rect 200776 150062 200850 150090
rect 201420 150062 201494 150090
rect 202064 150062 202138 150090
rect 202742 150078 202794 150084
rect 203352 150090 203380 152118
rect 203982 151328 204038 151337
rect 203982 151263 204038 151272
rect 203996 150090 204024 151263
rect 204640 150090 204668 153546
rect 205192 150226 205220 155926
rect 205284 154057 205312 159200
rect 205916 155916 205968 155922
rect 205916 155858 205968 155864
rect 205270 154048 205326 154057
rect 205270 153983 205326 153992
rect 205192 150198 205358 150226
rect 198246 149940 198274 150062
rect 198890 149940 198918 150062
rect 199534 149940 199562 150062
rect 200178 149940 200206 150062
rect 200822 149940 200850 150062
rect 201466 149940 201494 150062
rect 202110 149940 202138 150062
rect 202754 149940 202782 150078
rect 203352 150062 203426 150090
rect 203996 150062 204070 150090
rect 204640 150062 204714 150090
rect 203398 149940 203426 150062
rect 204042 149940 204070 150062
rect 204686 149940 204714 150062
rect 205330 149940 205358 150198
rect 205928 150090 205956 155858
rect 206112 154193 206140 159200
rect 206940 155922 206968 159200
rect 206928 155916 206980 155922
rect 206928 155858 206980 155864
rect 207768 155689 207796 159200
rect 207848 156596 207900 156602
rect 207848 156538 207900 156544
rect 207754 155680 207810 155689
rect 207754 155615 207810 155624
rect 206098 154184 206154 154193
rect 206098 154119 206154 154128
rect 207202 151192 207258 151201
rect 207202 151127 207258 151136
rect 206560 150884 206612 150890
rect 206560 150826 206612 150832
rect 206572 150090 206600 150826
rect 207216 150090 207244 151127
rect 207860 150090 207888 156538
rect 208596 153610 208624 159200
rect 208674 155408 208730 155417
rect 208674 155343 208730 155352
rect 208584 153604 208636 153610
rect 208584 153546 208636 153552
rect 208688 151910 208716 155343
rect 208492 151904 208544 151910
rect 208492 151846 208544 151852
rect 208676 151904 208728 151910
rect 208676 151846 208728 151852
rect 208504 150090 208532 151846
rect 209424 150890 209452 159200
rect 209780 155984 209832 155990
rect 209780 155926 209832 155932
rect 209688 155848 209740 155854
rect 209688 155790 209740 155796
rect 209700 155530 209728 155790
rect 209608 155502 209728 155530
rect 209608 154698 209636 155502
rect 209792 155446 209820 155926
rect 209688 155440 209740 155446
rect 209688 155382 209740 155388
rect 209780 155440 209832 155446
rect 209780 155382 209832 155388
rect 209700 154698 209728 155382
rect 209596 154692 209648 154698
rect 209596 154634 209648 154640
rect 209688 154692 209740 154698
rect 209688 154634 209740 154640
rect 209778 153640 209834 153649
rect 209778 153575 209834 153584
rect 209412 150884 209464 150890
rect 209412 150826 209464 150832
rect 209136 150816 209188 150822
rect 209136 150758 209188 150764
rect 209148 150090 209176 150758
rect 209792 150226 209820 153575
rect 210344 152182 210372 159200
rect 211172 152182 211200 159200
rect 211894 155000 211950 155009
rect 212000 154970 212028 159200
rect 212538 155000 212594 155009
rect 211894 154935 211896 154944
rect 211948 154935 211950 154944
rect 211988 154964 212040 154970
rect 211896 154906 211948 154912
rect 211988 154906 212040 154912
rect 212448 154964 212500 154970
rect 212538 154935 212540 154944
rect 212448 154906 212500 154912
rect 212592 154935 212594 154944
rect 212540 154906 212592 154912
rect 212264 153944 212316 153950
rect 212264 153886 212316 153892
rect 210332 152176 210384 152182
rect 210332 152118 210384 152124
rect 211160 152176 211212 152182
rect 211160 152118 211212 152124
rect 210424 152108 210476 152114
rect 210424 152050 210476 152056
rect 210436 150226 210464 152050
rect 211068 151904 211120 151910
rect 211068 151846 211120 151852
rect 211080 150226 211108 151846
rect 211620 150748 211672 150754
rect 211620 150690 211672 150696
rect 209792 150198 209866 150226
rect 210436 150198 210510 150226
rect 211080 150198 211154 150226
rect 205928 150062 206002 150090
rect 206572 150062 206646 150090
rect 207216 150062 207290 150090
rect 207860 150062 207934 150090
rect 208504 150062 208578 150090
rect 209148 150062 209222 150090
rect 205974 149940 206002 150062
rect 206618 149940 206646 150062
rect 207262 149940 207290 150062
rect 207906 149940 207934 150062
rect 208550 149940 208578 150062
rect 209194 149940 209222 150062
rect 209838 149940 209866 150198
rect 210482 149940 210510 150198
rect 211126 149940 211154 150198
rect 211632 150090 211660 150690
rect 212276 150226 212304 153886
rect 212460 153490 212488 154906
rect 212828 153950 212856 159200
rect 213656 155038 213684 159200
rect 214196 156664 214248 156670
rect 214196 156606 214248 156612
rect 213092 155032 213144 155038
rect 213092 154974 213144 154980
rect 213644 155032 213696 155038
rect 213644 154974 213696 154980
rect 212816 153944 212868 153950
rect 212816 153886 212868 153892
rect 212460 153462 213040 153490
rect 213012 153338 213040 153462
rect 212908 153332 212960 153338
rect 212908 153274 212960 153280
rect 213000 153332 213052 153338
rect 213000 153274 213052 153280
rect 212920 150226 212948 153274
rect 213104 152250 213132 154974
rect 213092 152244 213144 152250
rect 213092 152186 213144 152192
rect 213552 152040 213604 152046
rect 213552 151982 213604 151988
rect 213564 150226 213592 151982
rect 214208 150226 214236 156606
rect 214484 155417 214512 159200
rect 214470 155408 214526 155417
rect 214470 155343 214526 155352
rect 214380 154964 214432 154970
rect 214380 154906 214432 154912
rect 214564 154964 214616 154970
rect 214564 154906 214616 154912
rect 214392 152046 214420 154906
rect 214576 154630 214604 154906
rect 214564 154624 214616 154630
rect 214564 154566 214616 154572
rect 215312 153882 215340 159200
rect 216140 156670 216168 159200
rect 216128 156664 216180 156670
rect 216128 156606 216180 156612
rect 216496 155032 216548 155038
rect 216496 154974 216548 154980
rect 216508 154630 216536 154974
rect 216496 154624 216548 154630
rect 216496 154566 216548 154572
rect 214840 153876 214892 153882
rect 214840 153818 214892 153824
rect 215300 153876 215352 153882
rect 215300 153818 215352 153824
rect 214380 152040 214432 152046
rect 214380 151982 214432 151988
rect 214852 150226 214880 153818
rect 215482 152416 215538 152425
rect 215482 152351 215538 152360
rect 215496 150226 215524 152351
rect 216128 152244 216180 152250
rect 216128 152186 216180 152192
rect 216140 150226 216168 152186
rect 217060 152114 217088 159200
rect 217416 154080 217468 154086
rect 217416 154022 217468 154028
rect 217508 154080 217560 154086
rect 217508 154022 217560 154028
rect 217048 152108 217100 152114
rect 217048 152050 217100 152056
rect 216772 151088 216824 151094
rect 216772 151030 216824 151036
rect 212276 150198 212350 150226
rect 212920 150198 212994 150226
rect 213564 150198 213638 150226
rect 214208 150198 214282 150226
rect 214852 150198 214926 150226
rect 215496 150198 215570 150226
rect 216140 150198 216214 150226
rect 211632 150062 211706 150090
rect 211678 149940 211706 150062
rect 212322 149940 212350 150198
rect 212966 149940 212994 150198
rect 213610 149940 213638 150198
rect 214254 149940 214282 150198
rect 214898 149940 214926 150198
rect 215542 149940 215570 150198
rect 216186 149940 216214 150198
rect 216784 150090 216812 151030
rect 217428 150226 217456 154022
rect 217520 153950 217548 154022
rect 217508 153944 217560 153950
rect 217508 153886 217560 153892
rect 217600 153944 217652 153950
rect 217600 153886 217652 153892
rect 217612 153338 217640 153886
rect 217692 153876 217744 153882
rect 217692 153818 217744 153824
rect 217704 153338 217732 153818
rect 217600 153332 217652 153338
rect 217600 153274 217652 153280
rect 217692 153332 217744 153338
rect 217692 153274 217744 153280
rect 217888 152425 217916 159200
rect 218244 156732 218296 156738
rect 218244 156674 218296 156680
rect 218058 154320 218114 154329
rect 218058 154255 218114 154264
rect 217874 152416 217930 152425
rect 217874 152351 217930 152360
rect 218072 150226 218100 154255
rect 217428 150198 217502 150226
rect 218072 150198 218146 150226
rect 218256 150210 218284 156674
rect 218716 153882 218744 159200
rect 219544 156738 219572 159200
rect 220372 159174 220492 159200
rect 219532 156732 219584 156738
rect 219532 156674 219584 156680
rect 220740 154986 220768 159310
rect 221186 159200 221242 160400
rect 222014 159200 222070 160400
rect 222842 159200 222898 160400
rect 223762 159200 223818 160400
rect 224590 159200 224646 160400
rect 225418 159200 225474 160400
rect 226246 159200 226302 160400
rect 227074 159200 227130 160400
rect 227902 159200 227958 160400
rect 228730 159200 228786 160400
rect 229650 159200 229706 160400
rect 230478 159200 230534 160400
rect 231306 159200 231362 160400
rect 232134 159202 232190 160400
rect 232240 159310 232544 159338
rect 232240 159202 232268 159310
rect 232134 159200 232268 159202
rect 221200 155038 221228 159200
rect 221188 155032 221240 155038
rect 220740 154958 220860 154986
rect 221188 154974 221240 154980
rect 220728 154828 220780 154834
rect 220728 154770 220780 154776
rect 220740 154329 220768 154770
rect 220726 154320 220782 154329
rect 220726 154255 220782 154264
rect 219992 154012 220044 154018
rect 219992 153954 220044 153960
rect 220728 154012 220780 154018
rect 220728 153954 220780 153960
rect 218704 153876 218756 153882
rect 218704 153818 218756 153824
rect 218702 152552 218758 152561
rect 218702 152487 218758 152496
rect 218716 150226 218744 152487
rect 220004 150226 220032 153954
rect 220740 153270 220768 153954
rect 220728 153264 220780 153270
rect 220728 153206 220780 153212
rect 220832 152561 220860 154958
rect 222028 154086 222056 159200
rect 222856 155650 222884 159200
rect 223212 156120 223264 156126
rect 223212 156062 223264 156068
rect 222752 155644 222804 155650
rect 222752 155586 222804 155592
rect 222844 155644 222896 155650
rect 222844 155586 222896 155592
rect 222764 155553 222792 155586
rect 222566 155544 222622 155553
rect 222566 155479 222622 155488
rect 222750 155544 222806 155553
rect 222750 155479 222806 155488
rect 222580 155145 222608 155479
rect 222566 155136 222622 155145
rect 222566 155071 222622 155080
rect 221924 154080 221976 154086
rect 221924 154022 221976 154028
rect 222016 154080 222068 154086
rect 222016 154022 222068 154028
rect 221936 153338 221964 154022
rect 222568 153468 222620 153474
rect 222568 153410 222620 153416
rect 221924 153332 221976 153338
rect 221924 153274 221976 153280
rect 220818 152552 220874 152561
rect 220818 152487 220874 152496
rect 221280 152040 221332 152046
rect 221280 151982 221332 151988
rect 220636 151224 220688 151230
rect 220636 151166 220688 151172
rect 216784 150062 216858 150090
rect 216830 149940 216858 150062
rect 217474 149940 217502 150198
rect 218118 149940 218146 150198
rect 218244 150204 218296 150210
rect 218716 150198 218790 150226
rect 218244 150146 218296 150152
rect 218762 149940 218790 150198
rect 219394 150204 219446 150210
rect 220004 150198 220078 150226
rect 219394 150146 219446 150152
rect 219406 149940 219434 150146
rect 220050 149940 220078 150198
rect 220648 150090 220676 151166
rect 221292 150226 221320 151982
rect 221924 151156 221976 151162
rect 221924 151098 221976 151104
rect 221292 150198 221366 150226
rect 220648 150062 220722 150090
rect 220694 149940 220722 150062
rect 221338 149940 221366 150198
rect 221936 150090 221964 151098
rect 222580 150226 222608 153410
rect 223224 150226 223252 156062
rect 223488 155644 223540 155650
rect 223488 155586 223540 155592
rect 223580 155644 223632 155650
rect 223580 155586 223632 155592
rect 223500 151094 223528 155586
rect 223592 155553 223620 155586
rect 223578 155544 223634 155553
rect 223578 155479 223634 155488
rect 223578 155272 223634 155281
rect 223578 155207 223634 155216
rect 223592 152046 223620 155207
rect 223776 154834 223804 159200
rect 224132 156868 224184 156874
rect 224132 156810 224184 156816
rect 223764 154828 223816 154834
rect 223764 154770 223816 154776
rect 223580 152040 223632 152046
rect 223580 151982 223632 151988
rect 223856 151972 223908 151978
rect 223856 151914 223908 151920
rect 223488 151088 223540 151094
rect 223488 151030 223540 151036
rect 223868 150226 223896 151914
rect 224144 151814 224172 156810
rect 224604 151978 224632 159200
rect 225432 154086 225460 159200
rect 226260 156874 226288 159200
rect 226248 156868 226300 156874
rect 226248 156810 226300 156816
rect 226892 156800 226944 156806
rect 226892 156742 226944 156748
rect 225328 154080 225380 154086
rect 225328 154022 225380 154028
rect 225420 154080 225472 154086
rect 225420 154022 225472 154028
rect 225142 153776 225198 153785
rect 225142 153711 225198 153720
rect 224592 151972 224644 151978
rect 224592 151914 224644 151920
rect 224144 151786 224540 151814
rect 224512 150226 224540 151786
rect 225156 150226 225184 153711
rect 225340 153474 225368 154022
rect 225328 153468 225380 153474
rect 225328 153410 225380 153416
rect 225788 152516 225840 152522
rect 225788 152458 225840 152464
rect 225800 150226 225828 152458
rect 226432 152040 226484 152046
rect 226432 151982 226484 151988
rect 226444 150226 226472 151982
rect 226904 151814 226932 156742
rect 227088 154834 227116 159200
rect 227916 155281 227944 159200
rect 228456 155644 228508 155650
rect 228456 155586 228508 155592
rect 227902 155272 227958 155281
rect 227902 155207 227958 155216
rect 227810 155136 227866 155145
rect 227810 155071 227866 155080
rect 226984 154828 227036 154834
rect 226984 154770 227036 154776
rect 227076 154828 227128 154834
rect 227076 154770 227128 154776
rect 226996 151978 227024 154770
rect 227720 154148 227772 154154
rect 227720 154090 227772 154096
rect 226984 151972 227036 151978
rect 226984 151914 227036 151920
rect 226904 151786 227116 151814
rect 227088 150226 227116 151786
rect 227732 150226 227760 154090
rect 227824 151910 227852 155071
rect 228272 154012 228324 154018
rect 228272 153954 228324 153960
rect 228364 154012 228416 154018
rect 228364 153954 228416 153960
rect 227812 151904 227864 151910
rect 227812 151846 227864 151852
rect 228284 151814 228312 153954
rect 228376 153474 228404 153954
rect 228468 153474 228496 155586
rect 228744 154154 228772 159200
rect 229560 156936 229612 156942
rect 229560 156878 229612 156884
rect 228732 154148 228784 154154
rect 228732 154090 228784 154096
rect 228364 153468 228416 153474
rect 228364 153410 228416 153416
rect 228456 153468 228508 153474
rect 228456 153410 228508 153416
rect 229008 152720 229060 152726
rect 229008 152662 229060 152668
rect 228284 151786 228404 151814
rect 228376 150226 228404 151786
rect 229020 150226 229048 152662
rect 229572 151814 229600 156878
rect 229664 153785 229692 159200
rect 230388 155644 230440 155650
rect 230388 155586 230440 155592
rect 230400 155310 230428 155586
rect 230492 155310 230520 159200
rect 230388 155304 230440 155310
rect 230388 155246 230440 155252
rect 230480 155304 230532 155310
rect 230480 155246 230532 155252
rect 230296 154284 230348 154290
rect 230296 154226 230348 154232
rect 229650 153776 229706 153785
rect 229650 153711 229706 153720
rect 229572 151786 229692 151814
rect 229664 150226 229692 151786
rect 230308 150226 230336 154226
rect 230940 152584 230992 152590
rect 230940 152526 230992 152532
rect 230952 150226 230980 152526
rect 231320 152522 231348 159200
rect 232148 159174 232268 159200
rect 232228 157072 232280 157078
rect 232228 157014 232280 157020
rect 232042 155000 232098 155009
rect 232042 154935 232044 154944
rect 232096 154935 232098 154944
rect 232044 154906 232096 154912
rect 231308 152516 231360 152522
rect 231308 152458 231360 152464
rect 231584 151904 231636 151910
rect 231584 151846 231636 151852
rect 231596 150226 231624 151846
rect 232240 150226 232268 157014
rect 232516 155582 232544 159310
rect 232962 159200 233018 160400
rect 233790 159200 233846 160400
rect 234618 159200 234674 160400
rect 235446 159200 235502 160400
rect 236366 159200 236422 160400
rect 237194 159200 237250 160400
rect 238022 159200 238078 160400
rect 238850 159200 238906 160400
rect 239678 159200 239734 160400
rect 240506 159200 240562 160400
rect 241334 159200 241390 160400
rect 242162 159200 242218 160400
rect 243082 159200 243138 160400
rect 243910 159202 243966 160400
rect 244016 159310 244228 159338
rect 244016 159202 244044 159310
rect 243910 159200 244044 159202
rect 232976 156806 233004 159200
rect 232964 156800 233016 156806
rect 232964 156742 233016 156748
rect 232320 155576 232372 155582
rect 232320 155518 232372 155524
rect 232504 155576 232556 155582
rect 232504 155518 232556 155524
rect 233148 155576 233200 155582
rect 233148 155518 233200 155524
rect 232332 154970 232360 155518
rect 232320 154964 232372 154970
rect 232320 154906 232372 154912
rect 232964 154352 233016 154358
rect 232964 154294 233016 154300
rect 232976 154222 233004 154294
rect 233160 154290 233188 155518
rect 233238 155000 233294 155009
rect 233238 154935 233294 154944
rect 233148 154284 233200 154290
rect 233148 154226 233200 154232
rect 232872 154216 232924 154222
rect 232872 154158 232924 154164
rect 232964 154216 233016 154222
rect 232964 154158 233016 154164
rect 232884 150226 232912 154158
rect 233252 152726 233280 154935
rect 233804 154902 233832 159200
rect 234632 155650 234660 159200
rect 234804 157004 234856 157010
rect 234804 156946 234856 156952
rect 233976 155644 234028 155650
rect 233976 155586 234028 155592
rect 234620 155644 234672 155650
rect 234620 155586 234672 155592
rect 233884 155576 233936 155582
rect 233884 155518 233936 155524
rect 233700 154896 233752 154902
rect 233700 154838 233752 154844
rect 233792 154896 233844 154902
rect 233792 154838 233844 154844
rect 233712 154358 233740 154838
rect 233896 154834 233924 155518
rect 233988 154834 234016 155586
rect 234620 155236 234672 155242
rect 234620 155178 234672 155184
rect 233884 154828 233936 154834
rect 233884 154770 233936 154776
rect 233976 154828 234028 154834
rect 233976 154770 234028 154776
rect 233700 154352 233752 154358
rect 233514 154320 233570 154329
rect 233700 154294 233752 154300
rect 233514 154255 233570 154264
rect 233240 152720 233292 152726
rect 233240 152662 233292 152668
rect 233528 150226 233556 154255
rect 234632 152726 234660 155178
rect 233976 152720 234028 152726
rect 233976 152662 234028 152668
rect 234620 152720 234672 152726
rect 234620 152662 234672 152668
rect 233988 151978 234016 152662
rect 234160 152652 234212 152658
rect 234160 152594 234212 152600
rect 233976 151972 234028 151978
rect 233976 151914 234028 151920
rect 234172 150226 234200 152594
rect 234816 150226 234844 156946
rect 235264 154420 235316 154426
rect 235264 154362 235316 154368
rect 235356 154420 235408 154426
rect 235356 154362 235408 154368
rect 235276 151814 235304 154362
rect 235368 154222 235396 154362
rect 235460 154222 235488 159200
rect 236380 154358 236408 159200
rect 237208 155242 237236 159200
rect 237196 155236 237248 155242
rect 237196 155178 237248 155184
rect 238036 154902 238064 159200
rect 238668 155304 238720 155310
rect 238668 155246 238720 155252
rect 238760 155304 238812 155310
rect 238760 155246 238812 155252
rect 238024 154896 238076 154902
rect 238024 154838 238076 154844
rect 238574 154864 238630 154873
rect 237380 154828 237432 154834
rect 238680 154834 238708 155246
rect 238772 154902 238800 155246
rect 238864 155122 238892 159200
rect 239692 156942 239720 159200
rect 239956 157140 240008 157146
rect 239956 157082 240008 157088
rect 239680 156936 239732 156942
rect 239680 156878 239732 156884
rect 238864 155094 238984 155122
rect 238760 154896 238812 154902
rect 238760 154838 238812 154844
rect 238852 154896 238904 154902
rect 238852 154838 238904 154844
rect 238574 154799 238576 154808
rect 237380 154770 237432 154776
rect 238628 154799 238630 154808
rect 238668 154828 238720 154834
rect 238576 154770 238628 154776
rect 238668 154770 238720 154776
rect 236184 154352 236236 154358
rect 236184 154294 236236 154300
rect 236368 154352 236420 154358
rect 236368 154294 236420 154300
rect 235356 154216 235408 154222
rect 235356 154158 235408 154164
rect 235448 154216 235500 154222
rect 235448 154158 235500 154164
rect 236196 153474 236224 154294
rect 236092 153468 236144 153474
rect 236092 153410 236144 153416
rect 236184 153468 236236 153474
rect 236184 153410 236236 153416
rect 235276 151786 235488 151814
rect 235460 150226 235488 151786
rect 236104 150226 236132 153410
rect 236736 152720 236788 152726
rect 236736 152662 236788 152668
rect 236748 150226 236776 152662
rect 237392 152590 237420 154770
rect 238760 154760 238812 154766
rect 238864 154714 238892 154838
rect 238812 154708 238892 154714
rect 238760 154702 238892 154708
rect 238772 154686 238892 154702
rect 238036 154562 238248 154574
rect 238024 154556 238248 154562
rect 238076 154546 238248 154556
rect 238024 154498 238076 154504
rect 238220 154426 238248 154546
rect 238956 154494 238984 155094
rect 239034 154864 239090 154873
rect 239034 154799 239036 154808
rect 239088 154799 239090 154808
rect 239036 154770 239088 154776
rect 238944 154488 238996 154494
rect 238944 154430 238996 154436
rect 238116 154420 238168 154426
rect 238116 154362 238168 154368
rect 238208 154420 238260 154426
rect 238208 154362 238260 154368
rect 237380 152584 237432 152590
rect 237380 152526 237432 152532
rect 237380 151292 237432 151298
rect 237380 151234 237432 151240
rect 222580 150198 222654 150226
rect 223224 150198 223298 150226
rect 223868 150198 223942 150226
rect 224512 150198 224586 150226
rect 225156 150198 225230 150226
rect 225800 150198 225874 150226
rect 226444 150198 226518 150226
rect 227088 150198 227162 150226
rect 227732 150198 227806 150226
rect 228376 150198 228450 150226
rect 229020 150198 229094 150226
rect 229664 150198 229738 150226
rect 230308 150198 230382 150226
rect 230952 150198 231026 150226
rect 231596 150198 231670 150226
rect 232240 150198 232314 150226
rect 232884 150198 232958 150226
rect 233528 150198 233602 150226
rect 234172 150198 234246 150226
rect 234816 150198 234890 150226
rect 235460 150198 235534 150226
rect 236104 150198 236178 150226
rect 236748 150198 236822 150226
rect 221936 150062 222010 150090
rect 221982 149940 222010 150062
rect 222626 149940 222654 150198
rect 223270 149940 223298 150198
rect 223914 149940 223942 150198
rect 224558 149940 224586 150198
rect 225202 149940 225230 150198
rect 225846 149940 225874 150198
rect 226490 149940 226518 150198
rect 227134 149940 227162 150198
rect 227778 149940 227806 150198
rect 228422 149940 228450 150198
rect 229066 149940 229094 150198
rect 229710 149940 229738 150198
rect 230354 149940 230382 150198
rect 230998 149940 231026 150198
rect 231642 149940 231670 150198
rect 232286 149940 232314 150198
rect 232930 149940 232958 150198
rect 233574 149940 233602 150198
rect 234218 149940 234246 150198
rect 234862 149940 234890 150198
rect 235506 149940 235534 150198
rect 236150 149940 236178 150198
rect 236794 149940 236822 150198
rect 237392 150090 237420 151234
rect 238128 150226 238156 154362
rect 239312 152788 239364 152794
rect 239312 152730 239364 152736
rect 238668 150544 238720 150550
rect 238668 150486 238720 150492
rect 238082 150198 238156 150226
rect 237392 150062 237466 150090
rect 237438 149940 237466 150062
rect 238082 149940 238110 150198
rect 238680 150090 238708 150486
rect 239324 150226 239352 152730
rect 239968 150226 239996 157082
rect 240520 155786 240548 159200
rect 240416 155780 240468 155786
rect 240416 155722 240468 155728
rect 240508 155780 240560 155786
rect 240508 155722 240560 155728
rect 240428 155553 240456 155722
rect 240414 155544 240470 155553
rect 240414 155479 240470 155488
rect 241348 155242 241376 159200
rect 240508 155236 240560 155242
rect 240508 155178 240560 155184
rect 241336 155236 241388 155242
rect 241336 155178 241388 155184
rect 240520 152726 240548 155178
rect 241428 154964 241480 154970
rect 241428 154906 241480 154912
rect 240600 154420 240652 154426
rect 240600 154362 240652 154368
rect 240508 152720 240560 152726
rect 240508 152662 240560 152668
rect 240612 150226 240640 154362
rect 241440 153474 241468 154906
rect 242176 154426 242204 159200
rect 242440 157208 242492 157214
rect 242440 157150 242492 157156
rect 242164 154420 242216 154426
rect 242164 154362 242216 154368
rect 241244 153468 241296 153474
rect 241244 153410 241296 153416
rect 241428 153468 241480 153474
rect 241428 153410 241480 153416
rect 241256 150226 241284 153410
rect 241888 152584 241940 152590
rect 241888 152526 241940 152532
rect 241900 150226 241928 152526
rect 242452 150226 242480 157150
rect 243096 157010 243124 159200
rect 243924 159174 244044 159200
rect 243084 157004 243136 157010
rect 243084 156946 243136 156952
rect 243544 155644 243596 155650
rect 243544 155586 243596 155592
rect 242990 155544 243046 155553
rect 242990 155479 243046 155488
rect 243004 155378 243032 155479
rect 242900 155372 242952 155378
rect 242900 155314 242952 155320
rect 242992 155372 243044 155378
rect 242992 155314 243044 155320
rect 242912 152794 242940 155314
rect 243556 154970 243584 155586
rect 243544 154964 243596 154970
rect 243544 154906 243596 154912
rect 244200 154578 244228 159310
rect 244738 159200 244794 160400
rect 245566 159200 245622 160400
rect 246394 159200 246450 160400
rect 247222 159200 247278 160400
rect 248050 159200 248106 160400
rect 248878 159200 248934 160400
rect 249798 159200 249854 160400
rect 250626 159200 250682 160400
rect 251454 159200 251510 160400
rect 252282 159200 252338 160400
rect 253110 159200 253166 160400
rect 253938 159200 253994 160400
rect 254766 159200 254822 160400
rect 255594 159200 255650 160400
rect 256514 159200 256570 160400
rect 257342 159200 257398 160400
rect 258170 159200 258226 160400
rect 258998 159200 259054 160400
rect 259826 159200 259882 160400
rect 260654 159200 260710 160400
rect 261482 159200 261538 160400
rect 262402 159200 262458 160400
rect 263230 159202 263286 160400
rect 263336 159310 263548 159338
rect 263336 159202 263364 159310
rect 263230 159200 263364 159202
rect 244556 155984 244608 155990
rect 244556 155926 244608 155932
rect 244568 155718 244596 155926
rect 244556 155712 244608 155718
rect 244556 155654 244608 155660
rect 244752 155378 244780 159200
rect 244832 155780 244884 155786
rect 244832 155722 244884 155728
rect 244648 155372 244700 155378
rect 244648 155314 244700 155320
rect 244740 155372 244792 155378
rect 244740 155314 244792 155320
rect 244660 155258 244688 155314
rect 244844 155258 244872 155722
rect 244660 155230 244872 155258
rect 245476 155304 245528 155310
rect 245476 155246 245528 155252
rect 243084 154556 243136 154562
rect 244200 154550 244320 154578
rect 243084 154498 243136 154504
rect 242900 152788 242952 152794
rect 242900 152730 242952 152736
rect 243096 150226 243124 154498
rect 243728 152856 243780 152862
rect 243728 152798 243780 152804
rect 243544 152584 243596 152590
rect 243544 152526 243596 152532
rect 243556 152386 243584 152526
rect 243544 152380 243596 152386
rect 243544 152322 243596 152328
rect 243740 150226 243768 152798
rect 244292 152658 244320 154550
rect 245488 152930 245516 155246
rect 245580 154562 245608 159200
rect 246304 155984 246356 155990
rect 246304 155926 246356 155932
rect 246316 155718 246344 155926
rect 246304 155712 246356 155718
rect 246304 155654 246356 155660
rect 245568 154556 245620 154562
rect 245568 154498 245620 154504
rect 245660 153808 245712 153814
rect 245660 153750 245712 153756
rect 244372 152924 244424 152930
rect 244372 152866 244424 152872
rect 245476 152924 245528 152930
rect 245476 152866 245528 152872
rect 244280 152652 244332 152658
rect 244280 152594 244332 152600
rect 239324 150198 239398 150226
rect 239968 150198 240042 150226
rect 240612 150198 240686 150226
rect 241256 150198 241330 150226
rect 241900 150198 241974 150226
rect 242452 150198 242526 150226
rect 243096 150198 243170 150226
rect 243740 150198 243814 150226
rect 238680 150062 238754 150090
rect 238726 149940 238754 150062
rect 239370 149940 239398 150198
rect 240014 149940 240042 150198
rect 240658 149940 240686 150198
rect 241302 149940 241330 150198
rect 241946 149940 241974 150198
rect 242498 149940 242526 150198
rect 243142 149940 243170 150198
rect 243786 149940 243814 150198
rect 244384 150090 244412 152866
rect 245016 150612 245068 150618
rect 245016 150554 245068 150560
rect 245028 150090 245056 150554
rect 245672 150090 245700 153750
rect 246304 153468 246356 153474
rect 246304 153410 246356 153416
rect 246316 150090 246344 153410
rect 246408 151162 246436 159200
rect 247236 154902 247264 159200
rect 248064 155310 248092 159200
rect 248144 155780 248196 155786
rect 248144 155722 248196 155728
rect 248052 155304 248104 155310
rect 248052 155246 248104 155252
rect 247132 154896 247184 154902
rect 247132 154838 247184 154844
rect 247224 154896 247276 154902
rect 247224 154838 247276 154844
rect 247144 153678 247172 154838
rect 247132 153672 247184 153678
rect 247132 153614 247184 153620
rect 246948 152788 247000 152794
rect 246948 152730 247000 152736
rect 246396 151156 246448 151162
rect 246396 151098 246448 151104
rect 246960 150090 246988 152730
rect 248156 152386 248184 155722
rect 248892 154562 248920 159200
rect 249812 157078 249840 159200
rect 250168 157276 250220 157282
rect 250168 157218 250220 157224
rect 249800 157072 249852 157078
rect 249800 157014 249852 157020
rect 249064 155780 249116 155786
rect 249064 155722 249116 155728
rect 249076 155514 249104 155722
rect 249064 155508 249116 155514
rect 249064 155450 249116 155456
rect 249156 155508 249208 155514
rect 249156 155450 249208 155456
rect 249168 155174 249196 155450
rect 249156 155168 249208 155174
rect 249156 155110 249208 155116
rect 248788 154556 248840 154562
rect 248788 154498 248840 154504
rect 248880 154556 248932 154562
rect 248880 154498 248932 154504
rect 248984 154550 249196 154578
rect 248800 154442 248828 154498
rect 248984 154442 249012 154550
rect 249168 154494 249196 154550
rect 248800 154414 249012 154442
rect 249064 154488 249116 154494
rect 249064 154430 249116 154436
rect 249156 154488 249208 154494
rect 249156 154430 249208 154436
rect 248236 153740 248288 153746
rect 248236 153682 248288 153688
rect 248144 152380 248196 152386
rect 248144 152322 248196 152328
rect 247592 150680 247644 150686
rect 247592 150622 247644 150628
rect 247604 150090 247632 150622
rect 248248 150090 248276 153682
rect 249076 153474 249104 154430
rect 249064 153468 249116 153474
rect 249064 153410 249116 153416
rect 248880 152992 248932 152998
rect 248880 152934 248932 152940
rect 248892 150090 248920 152934
rect 249524 152584 249576 152590
rect 249524 152526 249576 152532
rect 249536 150090 249564 152526
rect 250180 150090 250208 157218
rect 250640 152998 250668 159200
rect 250812 157344 250864 157350
rect 250812 157286 250864 157292
rect 250628 152992 250680 152998
rect 250628 152934 250680 152940
rect 250824 150090 250852 157286
rect 251468 152862 251496 159200
rect 252296 153814 252324 159200
rect 252560 155372 252612 155378
rect 252560 155314 252612 155320
rect 252284 153808 252336 153814
rect 252284 153750 252336 153756
rect 251456 152856 251508 152862
rect 251456 152798 251508 152804
rect 252572 152386 252600 155314
rect 253124 155174 253152 159200
rect 253952 155378 253980 159200
rect 254780 155553 254808 159200
rect 255412 156188 255464 156194
rect 255412 156130 255464 156136
rect 254766 155544 254822 155553
rect 254124 155508 254176 155514
rect 254766 155479 254822 155488
rect 254124 155450 254176 155456
rect 253940 155372 253992 155378
rect 253940 155314 253992 155320
rect 253112 155168 253164 155174
rect 253112 155110 253164 155116
rect 253388 153740 253440 153746
rect 253388 153682 253440 153688
rect 252100 152380 252152 152386
rect 252100 152322 252152 152328
rect 252560 152380 252612 152386
rect 252560 152322 252612 152328
rect 251456 150476 251508 150482
rect 251456 150418 251508 150424
rect 251468 150090 251496 150418
rect 252112 150090 252140 152322
rect 252744 151360 252796 151366
rect 252744 151302 252796 151308
rect 252756 150090 252784 151302
rect 253400 150090 253428 153682
rect 254136 153066 254164 155450
rect 254032 153060 254084 153066
rect 254032 153002 254084 153008
rect 254124 153060 254176 153066
rect 254124 153002 254176 153008
rect 254044 150226 254072 153002
rect 254308 152992 254360 152998
rect 254308 152934 254360 152940
rect 254320 152658 254348 152934
rect 254308 152652 254360 152658
rect 254308 152594 254360 152600
rect 254676 151836 254728 151842
rect 254676 151778 254728 151784
rect 254688 150226 254716 151778
rect 255424 150226 255452 156130
rect 255608 153746 255636 159200
rect 255964 156528 256016 156534
rect 255964 156470 256016 156476
rect 255596 153740 255648 153746
rect 255596 153682 255648 153688
rect 254044 150198 254118 150226
rect 254688 150198 254762 150226
rect 244384 150062 244458 150090
rect 245028 150062 245102 150090
rect 245672 150062 245746 150090
rect 246316 150062 246390 150090
rect 246960 150062 247034 150090
rect 247604 150062 247678 150090
rect 248248 150062 248322 150090
rect 248892 150062 248966 150090
rect 249536 150062 249610 150090
rect 250180 150062 250254 150090
rect 250824 150062 250898 150090
rect 251468 150062 251542 150090
rect 252112 150062 252186 150090
rect 252756 150062 252830 150090
rect 253400 150062 253474 150090
rect 244430 149940 244458 150062
rect 245074 149940 245102 150062
rect 245718 149940 245746 150062
rect 246362 149940 246390 150062
rect 247006 149940 247034 150062
rect 247650 149940 247678 150062
rect 248294 149940 248322 150062
rect 248938 149940 248966 150062
rect 249582 149940 249610 150062
rect 250226 149940 250254 150062
rect 250870 149940 250898 150062
rect 251514 149940 251542 150062
rect 252158 149940 252186 150062
rect 252802 149940 252830 150062
rect 253446 149940 253474 150062
rect 254090 149940 254118 150198
rect 254734 149940 254762 150198
rect 255378 150198 255452 150226
rect 255976 150226 256004 156470
rect 256528 155530 256556 159200
rect 257252 155780 257304 155786
rect 257252 155722 257304 155728
rect 256436 155502 256556 155530
rect 256436 151230 256464 155502
rect 256516 153672 256568 153678
rect 256516 153614 256568 153620
rect 256528 151814 256556 153614
rect 256528 151786 256648 151814
rect 256424 151224 256476 151230
rect 256424 151166 256476 151172
rect 256620 150226 256648 151786
rect 257264 150226 257292 155722
rect 257356 155514 257384 159200
rect 257344 155508 257396 155514
rect 257344 155450 257396 155456
rect 258184 152862 258212 159200
rect 259012 153678 259040 159200
rect 259184 156460 259236 156466
rect 259184 156402 259236 156408
rect 259000 153672 259052 153678
rect 259000 153614 259052 153620
rect 258540 153536 258592 153542
rect 258540 153478 258592 153484
rect 258172 152856 258224 152862
rect 258172 152798 258224 152804
rect 257896 151496 257948 151502
rect 257896 151438 257948 151444
rect 255976 150198 256050 150226
rect 256620 150198 256694 150226
rect 257264 150198 257338 150226
rect 255378 149940 255406 150198
rect 256022 149940 256050 150198
rect 256666 149940 256694 150198
rect 257310 149940 257338 150198
rect 257908 150090 257936 151438
rect 258552 150226 258580 153478
rect 259196 150226 259224 156402
rect 259840 155854 259868 159200
rect 260012 156392 260064 156398
rect 260012 156334 260064 156340
rect 259828 155848 259880 155854
rect 259828 155790 259880 155796
rect 259828 153128 259880 153134
rect 259828 153070 259880 153076
rect 259840 150226 259868 153070
rect 260024 151814 260052 156334
rect 260668 155514 260696 159200
rect 261496 155786 261524 159200
rect 261392 155780 261444 155786
rect 261392 155722 261444 155728
rect 261484 155780 261536 155786
rect 261484 155722 261536 155728
rect 260564 155508 260616 155514
rect 260564 155450 260616 155456
rect 260656 155508 260708 155514
rect 260656 155450 260708 155456
rect 260576 155145 260604 155450
rect 260562 155136 260618 155145
rect 260196 155100 260248 155106
rect 261404 155106 261432 155722
rect 262128 155712 262180 155718
rect 262128 155654 262180 155660
rect 260562 155071 260618 155080
rect 261392 155100 261444 155106
rect 260196 155042 260248 155048
rect 261392 155042 261444 155048
rect 260208 153134 260236 155042
rect 260196 153128 260248 153134
rect 260196 153070 260248 153076
rect 261760 153060 261812 153066
rect 261760 153002 261812 153008
rect 260024 151786 260512 151814
rect 260484 150226 260512 151786
rect 261116 151428 261168 151434
rect 261116 151370 261168 151376
rect 258552 150198 258626 150226
rect 259196 150198 259270 150226
rect 259840 150198 259914 150226
rect 260484 150198 260558 150226
rect 257908 150062 257982 150090
rect 257954 149940 257982 150062
rect 258598 149940 258626 150198
rect 259242 149940 259270 150198
rect 259886 149940 259914 150198
rect 260530 149940 260558 150198
rect 261128 150090 261156 151370
rect 261772 150226 261800 153002
rect 262140 151814 262168 155654
rect 262416 154465 262444 159200
rect 263244 159174 263364 159200
rect 262864 155440 262916 155446
rect 262864 155382 262916 155388
rect 262876 155106 262904 155382
rect 262772 155100 262824 155106
rect 262772 155042 262824 155048
rect 262864 155100 262916 155106
rect 262864 155042 262916 155048
rect 262402 154456 262458 154465
rect 262402 154391 262458 154400
rect 262784 151978 262812 155042
rect 262680 151972 262732 151978
rect 262680 151914 262732 151920
rect 262772 151972 262824 151978
rect 262772 151914 262824 151920
rect 262692 151858 262720 151914
rect 262692 151842 262904 151858
rect 262692 151836 262916 151842
rect 262692 151830 262864 151836
rect 262140 151786 262444 151814
rect 262416 150226 262444 151786
rect 262864 151778 262916 151784
rect 263048 151564 263100 151570
rect 263048 151506 263100 151512
rect 261772 150198 261846 150226
rect 262416 150198 262490 150226
rect 261128 150062 261202 150090
rect 261174 149940 261202 150062
rect 261818 149940 261846 150198
rect 262462 149940 262490 150198
rect 263060 150090 263088 151506
rect 263520 151298 263548 159310
rect 264058 159200 264114 160400
rect 264886 159200 264942 160400
rect 265714 159200 265770 160400
rect 266542 159200 266598 160400
rect 267370 159200 267426 160400
rect 268198 159200 268254 160400
rect 269118 159200 269174 160400
rect 269946 159200 270002 160400
rect 270774 159200 270830 160400
rect 271602 159200 271658 160400
rect 272430 159200 272486 160400
rect 273258 159200 273314 160400
rect 274086 159200 274142 160400
rect 274914 159200 274970 160400
rect 275834 159200 275890 160400
rect 276662 159200 276718 160400
rect 277490 159200 277546 160400
rect 278318 159200 278374 160400
rect 279146 159200 279202 160400
rect 279974 159200 280030 160400
rect 280802 159200 280858 160400
rect 281630 159200 281686 160400
rect 282550 159200 282606 160400
rect 283378 159200 283434 160400
rect 284206 159200 284262 160400
rect 285034 159200 285090 160400
rect 285862 159200 285918 160400
rect 286690 159200 286746 160400
rect 287518 159200 287574 160400
rect 288346 159200 288402 160400
rect 289266 159200 289322 160400
rect 290094 159200 290150 160400
rect 290922 159200 290978 160400
rect 291750 159202 291806 160400
rect 291856 159310 292160 159338
rect 291856 159202 291884 159310
rect 291750 159200 291884 159202
rect 264072 155718 264100 159200
rect 264060 155712 264112 155718
rect 264060 155654 264112 155660
rect 264900 155446 264928 159200
rect 265164 156256 265216 156262
rect 265164 156198 265216 156204
rect 264888 155440 264940 155446
rect 264888 155382 264940 155388
rect 263690 155136 263746 155145
rect 263690 155071 263746 155080
rect 263704 154698 263732 155071
rect 263600 154692 263652 154698
rect 263600 154634 263652 154640
rect 263692 154692 263744 154698
rect 263692 154634 263744 154640
rect 264520 154692 264572 154698
rect 264520 154634 264572 154640
rect 263612 153066 263640 154634
rect 263692 153400 263744 153406
rect 263692 153342 263744 153348
rect 263600 153060 263652 153066
rect 263600 153002 263652 153008
rect 263508 151292 263560 151298
rect 263508 151234 263560 151240
rect 263704 150226 263732 153342
rect 264532 153202 264560 154634
rect 264428 153196 264480 153202
rect 264428 153138 264480 153144
rect 264520 153196 264572 153202
rect 264520 153138 264572 153144
rect 264440 150226 264468 153138
rect 264978 152688 265034 152697
rect 264978 152623 265034 152632
rect 263704 150198 263778 150226
rect 263060 150062 263134 150090
rect 263106 149940 263134 150062
rect 263750 149940 263778 150198
rect 264394 150198 264468 150226
rect 264992 150226 265020 152623
rect 264992 150198 265066 150226
rect 265176 150210 265204 156198
rect 265728 154329 265756 159200
rect 266452 155440 266504 155446
rect 266452 155382 266504 155388
rect 265714 154320 265770 154329
rect 265714 154255 265770 154264
rect 266464 152697 266492 155382
rect 266556 154698 266584 159200
rect 266728 155712 266780 155718
rect 266728 155654 266780 155660
rect 266544 154692 266596 154698
rect 266544 154634 266596 154640
rect 266740 152998 266768 155654
rect 267384 155446 267412 159200
rect 268108 156324 268160 156330
rect 268108 156266 268160 156272
rect 267372 155440 267424 155446
rect 267372 155382 267424 155388
rect 266912 153128 266964 153134
rect 266912 153070 266964 153076
rect 266728 152992 266780 152998
rect 266728 152934 266780 152940
rect 266450 152688 266506 152697
rect 266450 152623 266506 152632
rect 265624 151768 265676 151774
rect 265624 151710 265676 151716
rect 264394 149940 264422 150198
rect 265038 149940 265066 150198
rect 265164 150204 265216 150210
rect 265164 150146 265216 150152
rect 265636 150090 265664 151710
rect 266924 150226 266952 153070
rect 267556 151972 267608 151978
rect 267556 151914 267608 151920
rect 267568 150226 267596 151914
rect 268120 151814 268148 156266
rect 268212 155718 268240 159200
rect 268200 155712 268252 155718
rect 268200 155654 268252 155660
rect 269028 155100 269080 155106
rect 269028 155042 269080 155048
rect 269040 151978 269068 155042
rect 269132 153542 269160 159200
rect 269960 155106 269988 159200
rect 270788 155922 270816 159200
rect 270224 155916 270276 155922
rect 270224 155858 270276 155864
rect 270776 155916 270828 155922
rect 270776 155858 270828 155864
rect 269948 155100 270000 155106
rect 269948 155042 270000 155048
rect 269120 153536 269172 153542
rect 269120 153478 269172 153484
rect 270236 153105 270264 155858
rect 271512 154624 271564 154630
rect 271512 154566 271564 154572
rect 271616 154578 271644 159200
rect 270222 153096 270278 153105
rect 270222 153031 270278 153040
rect 269486 152824 269542 152833
rect 269486 152759 269542 152768
rect 269028 151972 269080 151978
rect 269028 151914 269080 151920
rect 268120 151786 268240 151814
rect 268212 150226 268240 151786
rect 268844 151700 268896 151706
rect 268844 151642 268896 151648
rect 266314 150204 266366 150210
rect 266924 150198 266998 150226
rect 267568 150198 267642 150226
rect 268212 150198 268286 150226
rect 266314 150146 266366 150152
rect 265636 150062 265710 150090
rect 265682 149940 265710 150062
rect 266326 149940 266354 150146
rect 266970 149940 266998 150198
rect 267614 149940 267642 150198
rect 268258 149940 268286 150198
rect 268856 150090 268884 151642
rect 269500 150226 269528 152759
rect 271524 151842 271552 154566
rect 271616 154550 271920 154578
rect 271892 153134 271920 154550
rect 272444 153406 272472 159200
rect 272536 155638 272840 155666
rect 272536 155582 272564 155638
rect 272524 155576 272576 155582
rect 272524 155518 272576 155524
rect 272708 155576 272760 155582
rect 272708 155518 272760 155524
rect 272524 155440 272576 155446
rect 272720 155428 272748 155518
rect 272812 155446 272840 155638
rect 272576 155400 272748 155428
rect 272800 155440 272852 155446
rect 272524 155382 272576 155388
rect 272800 155382 272852 155388
rect 273272 155174 273300 159200
rect 273350 155680 273406 155689
rect 273350 155615 273406 155624
rect 272616 155168 272668 155174
rect 272616 155110 272668 155116
rect 273260 155168 273312 155174
rect 273260 155110 273312 155116
rect 272628 154698 272656 155110
rect 272616 154692 272668 154698
rect 272616 154634 272668 154640
rect 273258 153912 273314 153921
rect 273258 153847 273314 153856
rect 272432 153400 272484 153406
rect 272432 153342 272484 153348
rect 271880 153128 271932 153134
rect 271880 153070 271932 153076
rect 272706 153096 272762 153105
rect 272064 153060 272116 153066
rect 272706 153031 272762 153040
rect 272064 153002 272116 153008
rect 270132 151836 270184 151842
rect 270132 151778 270184 151784
rect 271512 151836 271564 151842
rect 271512 151778 271564 151784
rect 270144 150226 270172 151778
rect 270776 151632 270828 151638
rect 270776 151574 270828 151580
rect 269500 150198 269574 150226
rect 270144 150198 270218 150226
rect 268856 150062 268930 150090
rect 268902 149940 268930 150062
rect 269546 149940 269574 150198
rect 270190 149940 270218 150198
rect 270788 150090 270816 151574
rect 271420 151020 271472 151026
rect 271420 150962 271472 150968
rect 271432 150090 271460 150962
rect 272076 150226 272104 153002
rect 272720 150226 272748 153031
rect 273272 150226 273300 153847
rect 273364 151881 273392 155615
rect 274100 155446 274128 159200
rect 274928 155689 274956 159200
rect 274914 155680 274970 155689
rect 274914 155615 274970 155624
rect 273996 155440 274048 155446
rect 273996 155382 274048 155388
rect 274088 155440 274140 155446
rect 274088 155382 274140 155388
rect 274008 152538 274036 155382
rect 275742 154048 275798 154057
rect 275742 153983 275798 153992
rect 274008 152510 274772 152538
rect 274548 152448 274600 152454
rect 274548 152390 274600 152396
rect 274640 152448 274692 152454
rect 274640 152390 274692 152396
rect 273350 151872 273406 151881
rect 273350 151807 273406 151816
rect 273904 150952 273956 150958
rect 273904 150894 273956 150900
rect 272076 150198 272150 150226
rect 272720 150198 272794 150226
rect 273272 150198 273346 150226
rect 270788 150062 270862 150090
rect 271432 150062 271506 150090
rect 270834 149940 270862 150062
rect 271478 149940 271506 150062
rect 272122 149940 272150 150198
rect 272766 149940 272794 150198
rect 273318 149940 273346 150198
rect 273916 150090 273944 150894
rect 274560 150226 274588 152390
rect 274652 151842 274680 152390
rect 274744 151842 274772 152510
rect 275192 152312 275244 152318
rect 275192 152254 275244 152260
rect 274640 151836 274692 151842
rect 274640 151778 274692 151784
rect 274732 151836 274784 151842
rect 274732 151778 274784 151784
rect 275204 150226 275232 152254
rect 275756 151814 275784 153983
rect 275848 153921 275876 159200
rect 276478 154184 276534 154193
rect 276478 154119 276534 154128
rect 275834 153912 275890 153921
rect 275834 153847 275890 153856
rect 275756 151786 275876 151814
rect 275848 150226 275876 151786
rect 276492 150226 276520 154119
rect 276676 153134 276704 159200
rect 277216 155916 277268 155922
rect 277216 155858 277268 155864
rect 276664 153128 276716 153134
rect 276664 153070 276716 153076
rect 277228 151978 277256 155858
rect 277504 155854 277532 159200
rect 277492 155848 277544 155854
rect 277492 155790 277544 155796
rect 278332 152833 278360 159200
rect 278688 154692 278740 154698
rect 278688 154634 278740 154640
rect 278700 154057 278728 154634
rect 278686 154048 278742 154057
rect 278686 153983 278742 153992
rect 279160 153610 279188 159200
rect 279514 155408 279570 155417
rect 279514 155343 279570 155352
rect 278412 153604 278464 153610
rect 278412 153546 278464 153552
rect 279148 153604 279200 153610
rect 279148 153546 279200 153552
rect 278318 152824 278374 152833
rect 278318 152759 278374 152768
rect 277124 151972 277176 151978
rect 277124 151914 277176 151920
rect 277216 151972 277268 151978
rect 277216 151914 277268 151920
rect 277136 150226 277164 151914
rect 277766 151872 277822 151881
rect 277766 151807 277822 151816
rect 277780 150226 277808 151807
rect 278424 150226 278452 153546
rect 279528 152318 279556 155343
rect 279988 155038 280016 159200
rect 279884 155032 279936 155038
rect 279882 155000 279884 155009
rect 279976 155032 280028 155038
rect 279936 155000 279938 155009
rect 279976 154974 280028 154980
rect 279882 154935 279938 154944
rect 280816 154698 280844 159200
rect 281644 155922 281672 159200
rect 281632 155916 281684 155922
rect 281632 155858 281684 155864
rect 282460 155848 282512 155854
rect 282460 155790 282512 155796
rect 282092 155168 282144 155174
rect 282092 155110 282144 155116
rect 282184 155168 282236 155174
rect 282184 155110 282236 155116
rect 282104 154766 282132 155110
rect 282196 154834 282224 155110
rect 282184 154828 282236 154834
rect 282184 154770 282236 154776
rect 281448 154760 281500 154766
rect 281448 154702 281500 154708
rect 282092 154760 282144 154766
rect 282092 154702 282144 154708
rect 280804 154692 280856 154698
rect 280804 154634 280856 154640
rect 280988 153944 281040 153950
rect 280988 153886 281040 153892
rect 279516 152312 279568 152318
rect 279516 152254 279568 152260
rect 280344 152244 280396 152250
rect 280344 152186 280396 152192
rect 279700 152176 279752 152182
rect 279700 152118 279752 152124
rect 279056 150884 279108 150890
rect 279056 150826 279108 150832
rect 274560 150198 274634 150226
rect 275204 150198 275278 150226
rect 275848 150198 275922 150226
rect 276492 150198 276566 150226
rect 277136 150198 277210 150226
rect 277780 150198 277854 150226
rect 278424 150198 278498 150226
rect 273916 150062 273990 150090
rect 273962 149940 273990 150062
rect 274606 149940 274634 150198
rect 275250 149940 275278 150198
rect 275894 149940 275922 150198
rect 276538 149940 276566 150198
rect 277182 149940 277210 150198
rect 277826 149940 277854 150198
rect 278470 149940 278498 150198
rect 279068 150090 279096 150826
rect 279712 150226 279740 152118
rect 280356 150226 280384 152186
rect 281000 150226 281028 153886
rect 281460 152250 281488 154702
rect 281632 153332 281684 153338
rect 281632 153274 281684 153280
rect 281448 152244 281500 152250
rect 281448 152186 281500 152192
rect 281644 150226 281672 153274
rect 282276 152448 282328 152454
rect 282276 152390 282328 152396
rect 282288 150226 282316 152390
rect 282472 152182 282500 155790
rect 282564 153950 282592 159200
rect 283012 155984 283064 155990
rect 283012 155926 283064 155932
rect 282918 155000 282974 155009
rect 282918 154935 282974 154944
rect 282552 153944 282604 153950
rect 282552 153886 282604 153892
rect 282932 152454 282960 154935
rect 283024 153338 283052 155926
rect 283288 155848 283340 155854
rect 283288 155790 283340 155796
rect 283300 155174 283328 155790
rect 283392 155174 283420 159200
rect 284116 156664 284168 156670
rect 284116 156606 284168 156612
rect 283288 155168 283340 155174
rect 283288 155110 283340 155116
rect 283380 155168 283432 155174
rect 283380 155110 283432 155116
rect 283012 153332 283064 153338
rect 283012 153274 283064 153280
rect 283564 153264 283616 153270
rect 283564 153206 283616 153212
rect 282920 152448 282972 152454
rect 282920 152390 282972 152396
rect 282920 152312 282972 152318
rect 282920 152254 282972 152260
rect 282460 152176 282512 152182
rect 282460 152118 282512 152124
rect 279712 150198 279786 150226
rect 280356 150198 280430 150226
rect 281000 150198 281074 150226
rect 281644 150198 281718 150226
rect 282288 150198 282362 150226
rect 279068 150062 279142 150090
rect 279114 149940 279142 150062
rect 279758 149940 279786 150198
rect 280402 149940 280430 150198
rect 281046 149940 281074 150198
rect 281690 149940 281718 150198
rect 282334 149940 282362 150198
rect 282932 150090 282960 152254
rect 283576 150090 283604 153206
rect 284128 150226 284156 156606
rect 284220 155258 284248 159200
rect 284220 155230 284432 155258
rect 284300 155168 284352 155174
rect 284300 155110 284352 155116
rect 284312 153270 284340 155110
rect 284300 153264 284352 153270
rect 284300 153206 284352 153212
rect 284404 152250 284432 155230
rect 285048 154834 285076 159200
rect 285876 157334 285904 159200
rect 285876 157306 286272 157334
rect 285036 154828 285088 154834
rect 285036 154770 285088 154776
rect 286244 153882 286272 157306
rect 286704 155174 286732 159200
rect 286784 156732 286836 156738
rect 286784 156674 286836 156680
rect 286692 155168 286744 155174
rect 286692 155110 286744 155116
rect 286140 153876 286192 153882
rect 286140 153818 286192 153824
rect 286232 153876 286284 153882
rect 286232 153818 286284 153824
rect 285494 152416 285550 152425
rect 285494 152351 285550 152360
rect 284392 152244 284444 152250
rect 284392 152186 284444 152192
rect 284852 152108 284904 152114
rect 284852 152050 284904 152056
rect 284128 150198 284294 150226
rect 282932 150062 283006 150090
rect 283576 150062 283650 150090
rect 282978 149940 283006 150062
rect 283622 149940 283650 150062
rect 284266 149940 284294 150198
rect 284864 150090 284892 152050
rect 285508 150090 285536 152351
rect 286152 150090 286180 153818
rect 286796 150090 286824 156674
rect 287532 155854 287560 159200
rect 287336 155848 287388 155854
rect 287336 155790 287388 155796
rect 287520 155848 287572 155854
rect 287520 155790 287572 155796
rect 287060 154828 287112 154834
rect 287060 154770 287112 154776
rect 286968 154080 287020 154086
rect 286968 154022 287020 154028
rect 286980 153338 287008 154022
rect 286876 153332 286928 153338
rect 286876 153274 286928 153280
rect 286968 153332 287020 153338
rect 286968 153274 287020 153280
rect 286888 153241 286916 153274
rect 286874 153232 286930 153241
rect 286874 153167 286930 153176
rect 287072 152425 287100 154770
rect 287152 154216 287204 154222
rect 287152 154158 287204 154164
rect 287164 154086 287192 154158
rect 287152 154080 287204 154086
rect 287152 154022 287204 154028
rect 287058 152416 287114 152425
rect 287058 152351 287114 152360
rect 287348 152114 287376 155790
rect 288360 155038 288388 159200
rect 287704 155032 287756 155038
rect 287704 154974 287756 154980
rect 288348 155032 288400 155038
rect 288348 154974 288400 154980
rect 287520 154828 287572 154834
rect 287520 154770 287572 154776
rect 287532 154630 287560 154770
rect 287716 154698 287744 154974
rect 287704 154692 287756 154698
rect 287704 154634 287756 154640
rect 287520 154624 287572 154630
rect 287520 154566 287572 154572
rect 287796 154216 287848 154222
rect 287624 154164 287796 154170
rect 287624 154158 287848 154164
rect 287624 154154 287836 154158
rect 287612 154148 287836 154154
rect 287664 154142 287836 154148
rect 287612 154090 287664 154096
rect 289280 154018 289308 159200
rect 288716 154012 288768 154018
rect 288716 153954 288768 153960
rect 289268 154012 289320 154018
rect 289268 153954 289320 153960
rect 287426 152552 287482 152561
rect 287426 152487 287482 152496
rect 287336 152108 287388 152114
rect 287336 152050 287388 152056
rect 287440 150090 287468 152487
rect 288072 152448 288124 152454
rect 288072 152390 288124 152396
rect 288164 152448 288216 152454
rect 288164 152390 288216 152396
rect 288084 150090 288112 152390
rect 288176 152250 288204 152390
rect 288164 152244 288216 152250
rect 288164 152186 288216 152192
rect 288728 150090 288756 153954
rect 290108 152114 290136 159200
rect 290936 152250 290964 159200
rect 291764 159174 291884 159200
rect 291936 156868 291988 156874
rect 291936 156810 291988 156816
rect 291200 154828 291252 154834
rect 291200 154770 291252 154776
rect 291212 154154 291240 154770
rect 291200 154148 291252 154154
rect 291200 154090 291252 154096
rect 291292 153332 291344 153338
rect 291292 153274 291344 153280
rect 290924 152244 290976 152250
rect 290924 152186 290976 152192
rect 290004 152108 290056 152114
rect 290004 152050 290056 152056
rect 290096 152108 290148 152114
rect 290096 152050 290148 152056
rect 290016 151994 290044 152050
rect 290648 152040 290700 152046
rect 290016 151966 290136 151994
rect 290648 151982 290700 151988
rect 290108 151910 290136 151966
rect 290004 151904 290056 151910
rect 290004 151846 290056 151852
rect 290096 151904 290148 151910
rect 290096 151846 290148 151852
rect 289360 151088 289412 151094
rect 289360 151030 289412 151036
rect 289372 150090 289400 151030
rect 290016 150090 290044 151846
rect 290660 150090 290688 151982
rect 291304 150090 291332 153274
rect 291476 153264 291528 153270
rect 291474 153232 291476 153241
rect 291528 153232 291530 153241
rect 291474 153167 291530 153176
rect 291948 150090 291976 156810
rect 292132 154834 292160 159310
rect 292578 159200 292634 160400
rect 293406 159200 293462 160400
rect 294234 159200 294290 160400
rect 295154 159200 295210 160400
rect 295982 159200 296038 160400
rect 296810 159200 296866 160400
rect 297638 159200 297694 160400
rect 298466 159200 298522 160400
rect 299294 159200 299350 160400
rect 300122 159200 300178 160400
rect 300950 159200 301006 160400
rect 301870 159200 301926 160400
rect 302698 159200 302754 160400
rect 303526 159200 303582 160400
rect 304354 159200 304410 160400
rect 305182 159200 305238 160400
rect 306010 159200 306066 160400
rect 306838 159200 306894 160400
rect 307666 159200 307722 160400
rect 308586 159200 308642 160400
rect 309414 159200 309470 160400
rect 310242 159200 310298 160400
rect 311070 159202 311126 160400
rect 311176 159310 311572 159338
rect 311176 159202 311204 159310
rect 311070 159200 311204 159202
rect 292592 157334 292620 159200
rect 292592 157306 292988 157334
rect 292212 155984 292264 155990
rect 292212 155926 292264 155932
rect 292120 154828 292172 154834
rect 292120 154770 292172 154776
rect 292224 154630 292252 155926
rect 292580 155644 292632 155650
rect 292580 155586 292632 155592
rect 292592 155174 292620 155586
rect 292304 155168 292356 155174
rect 292304 155110 292356 155116
rect 292580 155168 292632 155174
rect 292580 155110 292632 155116
rect 292212 154624 292264 154630
rect 292212 154566 292264 154572
rect 292316 154442 292344 155110
rect 292394 155000 292450 155009
rect 292394 154935 292396 154944
rect 292448 154935 292450 154944
rect 292396 154906 292448 154912
rect 292488 154624 292540 154630
rect 292488 154566 292540 154572
rect 292500 154442 292528 154566
rect 292316 154414 292528 154442
rect 292684 154414 292896 154442
rect 292684 154358 292712 154414
rect 292672 154352 292724 154358
rect 292672 154294 292724 154300
rect 292304 154284 292356 154290
rect 292304 154226 292356 154232
rect 292316 154193 292344 154226
rect 292488 154216 292540 154222
rect 292302 154184 292358 154193
rect 292868 154193 292896 154414
rect 292960 154222 292988 157306
rect 293222 155272 293278 155281
rect 293222 155207 293278 155216
rect 293132 154828 293184 154834
rect 293132 154770 293184 154776
rect 292948 154216 293000 154222
rect 292488 154158 292540 154164
rect 292670 154184 292726 154193
rect 292302 154119 292358 154128
rect 292396 154080 292448 154086
rect 292396 154022 292448 154028
rect 292408 150142 292436 154022
rect 292500 150210 292528 154158
rect 292670 154119 292726 154128
rect 292854 154184 292910 154193
rect 292948 154158 293000 154164
rect 292854 154119 292910 154128
rect 292684 154086 292712 154119
rect 292672 154080 292724 154086
rect 292672 154022 292724 154028
rect 292764 152312 292816 152318
rect 292764 152254 292816 152260
rect 292776 152046 292804 152254
rect 293144 152250 293172 154770
rect 293132 152244 293184 152250
rect 293132 152186 293184 152192
rect 292764 152040 292816 152046
rect 292764 151982 292816 151988
rect 292580 151836 292632 151842
rect 292580 151778 292632 151784
rect 292488 150204 292540 150210
rect 292488 150146 292540 150152
rect 292396 150136 292448 150142
rect 284864 150062 284938 150090
rect 285508 150062 285582 150090
rect 286152 150062 286226 150090
rect 286796 150062 286870 150090
rect 287440 150062 287514 150090
rect 288084 150062 288158 150090
rect 288728 150062 288802 150090
rect 289372 150062 289446 150090
rect 290016 150062 290090 150090
rect 290660 150062 290734 150090
rect 291304 150062 291378 150090
rect 291948 150062 292022 150090
rect 292396 150078 292448 150084
rect 292592 150090 292620 151778
rect 293236 150090 293264 155207
rect 293420 154902 293448 159200
rect 294052 155304 294104 155310
rect 294052 155246 294104 155252
rect 293958 155000 294014 155009
rect 294064 154970 294092 155246
rect 294248 155242 294276 159200
rect 295168 155281 295196 159200
rect 295800 155984 295852 155990
rect 295800 155926 295852 155932
rect 295812 155854 295840 155926
rect 295708 155848 295760 155854
rect 295708 155790 295760 155796
rect 295800 155848 295852 155854
rect 295800 155790 295852 155796
rect 295154 155272 295210 155281
rect 294236 155236 294288 155242
rect 295154 155207 295210 155216
rect 294236 155178 294288 155184
rect 295720 155174 295748 155790
rect 295892 155644 295944 155650
rect 295892 155586 295944 155592
rect 295616 155168 295668 155174
rect 295616 155110 295668 155116
rect 295708 155168 295760 155174
rect 295904 155156 295932 155586
rect 295708 155110 295760 155116
rect 295812 155128 295932 155156
rect 295628 155020 295656 155110
rect 295812 155020 295840 155128
rect 295628 154992 295840 155020
rect 293958 154935 294014 154944
rect 294052 154964 294104 154970
rect 293408 154896 293460 154902
rect 293408 154838 293460 154844
rect 293972 151842 294000 154935
rect 294052 154906 294104 154912
rect 294328 154828 294380 154834
rect 294328 154770 294380 154776
rect 294340 154714 294368 154770
rect 294696 154760 294748 154766
rect 294340 154708 294696 154714
rect 294340 154702 294748 154708
rect 294340 154686 294736 154702
rect 295996 154290 296024 159200
rect 295984 154284 296036 154290
rect 295984 154226 296036 154232
rect 296444 154080 296496 154086
rect 296444 154022 296496 154028
rect 294510 153776 294566 153785
rect 294510 153711 294566 153720
rect 293960 151836 294012 151842
rect 293960 151778 294012 151784
rect 293914 150204 293966 150210
rect 293914 150146 293966 150152
rect 292592 150062 292666 150090
rect 293236 150062 293310 150090
rect 284910 149940 284938 150062
rect 285554 149940 285582 150062
rect 286198 149940 286226 150062
rect 286842 149940 286870 150062
rect 287486 149940 287514 150062
rect 288130 149940 288158 150062
rect 288774 149940 288802 150062
rect 289418 149940 289446 150062
rect 290062 149940 290090 150062
rect 290706 149940 290734 150062
rect 291350 149940 291378 150062
rect 291994 149940 292022 150062
rect 292638 149940 292666 150062
rect 293282 149940 293310 150062
rect 293926 149940 293954 150146
rect 294524 150090 294552 153711
rect 295800 152516 295852 152522
rect 295800 152458 295852 152464
rect 295064 152244 295116 152250
rect 295064 152186 295116 152192
rect 295524 152244 295576 152250
rect 295524 152186 295576 152192
rect 295076 152130 295104 152186
rect 295536 152130 295564 152186
rect 295076 152102 295288 152130
rect 295352 152114 295564 152130
rect 295260 152046 295288 152102
rect 295340 152108 295564 152114
rect 295392 152102 295564 152108
rect 295340 152050 295392 152056
rect 295156 152040 295208 152046
rect 295156 151982 295208 151988
rect 295248 152040 295300 152046
rect 295248 151982 295300 151988
rect 295168 150090 295196 151982
rect 295812 150090 295840 152458
rect 296456 150090 296484 154022
rect 296824 152046 296852 159200
rect 297652 157334 297680 159200
rect 297652 157306 297864 157334
rect 297088 156800 297140 156806
rect 297088 156742 297140 156748
rect 296812 152040 296864 152046
rect 296812 151982 296864 151988
rect 297100 150090 297128 156742
rect 297364 154148 297416 154154
rect 297364 154090 297416 154096
rect 297272 154080 297324 154086
rect 297272 154022 297324 154028
rect 297284 153474 297312 154022
rect 297376 153474 297404 154090
rect 297272 153468 297324 153474
rect 297272 153410 297324 153416
rect 297364 153468 297416 153474
rect 297364 153410 297416 153416
rect 297836 151910 297864 157306
rect 297732 151904 297784 151910
rect 297732 151846 297784 151852
rect 297824 151904 297876 151910
rect 297824 151846 297876 151852
rect 297744 150090 297772 151846
rect 298480 151842 298508 159200
rect 299308 154086 299336 159200
rect 299446 155922 299612 155938
rect 299434 155916 299624 155922
rect 299486 155910 299572 155916
rect 299434 155858 299486 155864
rect 299572 155858 299624 155864
rect 299492 155786 299612 155802
rect 299480 155780 299624 155786
rect 299532 155774 299572 155780
rect 299480 155722 299532 155728
rect 299572 155722 299624 155728
rect 300136 155650 300164 159200
rect 299664 155644 299716 155650
rect 300124 155644 300176 155650
rect 299716 155604 299980 155632
rect 299664 155586 299716 155592
rect 299572 155576 299624 155582
rect 299624 155524 299888 155530
rect 299572 155518 299888 155524
rect 299584 155502 299888 155518
rect 299664 155440 299716 155446
rect 299570 155408 299626 155417
rect 299756 155440 299808 155446
rect 299716 155388 299756 155394
rect 299664 155382 299808 155388
rect 299676 155366 299796 155382
rect 299860 155378 299888 155502
rect 299848 155372 299900 155378
rect 299570 155343 299572 155352
rect 299624 155343 299626 155352
rect 299572 155314 299624 155320
rect 299848 155314 299900 155320
rect 299480 155304 299532 155310
rect 299532 155252 299704 155258
rect 299480 155246 299704 155252
rect 299492 155230 299704 155246
rect 299400 155106 299520 155122
rect 299388 155100 299520 155106
rect 299440 155094 299520 155100
rect 299388 155042 299440 155048
rect 299492 154494 299520 155094
rect 299676 154873 299704 155230
rect 299662 154864 299718 154873
rect 299662 154799 299718 154808
rect 299952 154574 299980 155604
rect 300124 155586 300176 155592
rect 300964 155242 300992 159200
rect 300860 155236 300912 155242
rect 300860 155178 300912 155184
rect 300952 155236 301004 155242
rect 300952 155178 301004 155184
rect 300872 155106 300900 155178
rect 300860 155100 300912 155106
rect 300860 155042 300912 155048
rect 301884 154766 301912 159200
rect 302240 156936 302292 156942
rect 302240 156878 302292 156884
rect 301044 154760 301096 154766
rect 301044 154702 301096 154708
rect 301872 154760 301924 154766
rect 301872 154702 301924 154708
rect 299584 154546 299980 154574
rect 299480 154488 299532 154494
rect 299480 154430 299532 154436
rect 299296 154080 299348 154086
rect 299296 154022 299348 154028
rect 299584 152522 299612 154546
rect 299662 154184 299718 154193
rect 299662 154119 299718 154128
rect 299572 152516 299624 152522
rect 299572 152458 299624 152464
rect 298376 151836 298428 151842
rect 298376 151778 298428 151784
rect 298468 151836 298520 151842
rect 298468 151778 298520 151784
rect 298388 150090 298416 151778
rect 299066 150136 299118 150142
rect 294524 150062 294598 150090
rect 295168 150062 295242 150090
rect 295812 150062 295886 150090
rect 296456 150062 296530 150090
rect 297100 150062 297174 150090
rect 297744 150062 297818 150090
rect 298388 150062 298462 150090
rect 299066 150078 299118 150084
rect 299676 150090 299704 154119
rect 301056 152930 301084 154702
rect 301596 154148 301648 154154
rect 301596 154090 301648 154096
rect 300952 152924 301004 152930
rect 300952 152866 301004 152872
rect 301044 152924 301096 152930
rect 301044 152866 301096 152872
rect 300308 152720 300360 152726
rect 300308 152662 300360 152668
rect 300320 150090 300348 152662
rect 300964 150090 300992 152866
rect 301608 150090 301636 154090
rect 302252 150090 302280 156878
rect 302712 154222 302740 159200
rect 303540 157334 303568 159200
rect 303448 157306 303568 157334
rect 302792 155644 302844 155650
rect 302792 155586 302844 155592
rect 302884 155644 302936 155650
rect 302884 155586 302936 155592
rect 302804 155310 302832 155586
rect 302792 155304 302844 155310
rect 302792 155246 302844 155252
rect 302896 155242 302924 155586
rect 302884 155236 302936 155242
rect 302884 155178 302936 155184
rect 302700 154216 302752 154222
rect 302700 154158 302752 154164
rect 303448 152590 303476 157306
rect 304368 155242 304396 159200
rect 304724 157004 304776 157010
rect 304724 156946 304776 156952
rect 304356 155236 304408 155242
rect 304356 155178 304408 155184
rect 303526 154864 303582 154873
rect 303526 154799 303582 154808
rect 302516 152584 302568 152590
rect 302516 152526 302568 152532
rect 303436 152584 303488 152590
rect 303436 152526 303488 152532
rect 302528 151910 302556 152526
rect 302884 152516 302936 152522
rect 302884 152458 302936 152464
rect 302516 151904 302568 151910
rect 302516 151846 302568 151852
rect 302896 150090 302924 152458
rect 303540 150090 303568 154799
rect 304080 154352 304132 154358
rect 304080 154294 304132 154300
rect 304092 150090 304120 154294
rect 304736 150090 304764 156946
rect 305000 152652 305052 152658
rect 305052 152612 305132 152640
rect 305000 152594 305052 152600
rect 305104 150226 305132 152612
rect 305196 152590 305224 159200
rect 306024 154358 306052 159200
rect 306852 155582 306880 159200
rect 306840 155576 306892 155582
rect 306840 155518 306892 155524
rect 307116 155304 307168 155310
rect 307116 155246 307168 155252
rect 306380 155236 306432 155242
rect 306380 155178 306432 155184
rect 306932 155236 306984 155242
rect 306932 155178 306984 155184
rect 306012 154352 306064 154358
rect 306012 154294 306064 154300
rect 305184 152584 305236 152590
rect 305184 152526 305236 152532
rect 306012 152380 306064 152386
rect 306012 152322 306064 152328
rect 305104 150198 305454 150226
rect 294570 149940 294598 150062
rect 295214 149940 295242 150062
rect 295858 149940 295886 150062
rect 296502 149940 296530 150062
rect 297146 149940 297174 150062
rect 297790 149940 297818 150062
rect 298434 149940 298462 150062
rect 299078 149940 299106 150078
rect 299676 150062 299750 150090
rect 300320 150062 300394 150090
rect 300964 150062 301038 150090
rect 301608 150062 301682 150090
rect 302252 150062 302326 150090
rect 302896 150062 302970 150090
rect 303540 150062 303614 150090
rect 304092 150062 304166 150090
rect 304736 150062 304810 150090
rect 299722 149940 299750 150062
rect 300366 149940 300394 150062
rect 301010 149940 301038 150062
rect 301654 149940 301682 150062
rect 302298 149940 302326 150062
rect 302942 149940 302970 150062
rect 303586 149940 303614 150062
rect 304138 149940 304166 150062
rect 304782 149940 304810 150062
rect 305426 149940 305454 150198
rect 306024 150090 306052 152322
rect 306392 151842 306420 155178
rect 306944 154970 306972 155178
rect 306932 154964 306984 154970
rect 306932 154906 306984 154912
rect 306932 154828 306984 154834
rect 306932 154770 306984 154776
rect 306944 154562 306972 154770
rect 307128 154766 307156 155246
rect 307680 155242 307708 159200
rect 308600 155310 308628 159200
rect 309138 155408 309194 155417
rect 309138 155343 309194 155352
rect 308496 155304 308548 155310
rect 308496 155246 308548 155252
rect 308588 155304 308640 155310
rect 308588 155246 308640 155252
rect 307668 155236 307720 155242
rect 307668 155178 307720 155184
rect 307208 154964 307260 154970
rect 307208 154906 307260 154912
rect 307024 154760 307076 154766
rect 307024 154702 307076 154708
rect 307116 154760 307168 154766
rect 307116 154702 307168 154708
rect 307036 154578 307064 154702
rect 307220 154578 307248 154906
rect 306932 154556 306984 154562
rect 307036 154550 307248 154578
rect 306932 154498 306984 154504
rect 307116 154488 307168 154494
rect 307116 154430 307168 154436
rect 306656 154420 306708 154426
rect 306656 154362 306708 154368
rect 306932 154420 306984 154426
rect 306932 154362 306984 154368
rect 306380 151836 306432 151842
rect 306380 151778 306432 151784
rect 306668 150090 306696 154362
rect 306944 154306 306972 154362
rect 306944 154278 307064 154306
rect 307036 153814 307064 154278
rect 306932 153808 306984 153814
rect 306932 153750 306984 153756
rect 307024 153808 307076 153814
rect 307024 153750 307076 153756
rect 306944 153626 306972 153750
rect 307128 153626 307156 154430
rect 306944 153598 307156 153626
rect 307944 152924 307996 152930
rect 307944 152866 307996 152872
rect 307300 151156 307352 151162
rect 307300 151098 307352 151104
rect 307312 150090 307340 151098
rect 307956 150090 307984 152866
rect 308508 150226 308536 155246
rect 309152 152930 309180 155343
rect 309428 154426 309456 159200
rect 309876 157072 309928 157078
rect 309876 157014 309928 157020
rect 309232 154420 309284 154426
rect 309232 154362 309284 154368
rect 309416 154420 309468 154426
rect 309416 154362 309468 154368
rect 309140 152924 309192 152930
rect 309140 152866 309192 152872
rect 308508 150198 308674 150226
rect 306024 150062 306098 150090
rect 306668 150062 306742 150090
rect 307312 150062 307386 150090
rect 307956 150062 308030 150090
rect 306070 149940 306098 150062
rect 306714 149940 306742 150062
rect 307358 149940 307386 150062
rect 308002 149940 308030 150062
rect 308646 149940 308674 150198
rect 309244 150090 309272 154362
rect 309888 150090 309916 157014
rect 310256 154834 310284 159200
rect 311084 159174 311204 159200
rect 310610 155544 310666 155553
rect 310610 155479 310666 155488
rect 310244 154828 310296 154834
rect 310244 154770 310296 154776
rect 310520 152720 310572 152726
rect 310520 152662 310572 152668
rect 310532 150226 310560 152662
rect 310624 152386 310652 155479
rect 311438 155000 311494 155009
rect 311438 154935 311494 154944
rect 311452 154698 311480 154935
rect 311440 154692 311492 154698
rect 311440 154634 311492 154640
rect 311440 154488 311492 154494
rect 311440 154430 311492 154436
rect 311164 152788 311216 152794
rect 311164 152730 311216 152736
rect 310612 152380 310664 152386
rect 310612 152322 310664 152328
rect 310532 150198 310606 150226
rect 309244 150062 309318 150090
rect 309888 150062 309962 150090
rect 309290 149940 309318 150062
rect 309934 149940 309962 150062
rect 310578 149940 310606 150198
rect 311176 150090 311204 152730
rect 311452 150226 311480 154430
rect 311544 152794 311572 159310
rect 311898 159200 311954 160400
rect 312726 159200 312782 160400
rect 313554 159200 313610 160400
rect 314382 159200 314438 160400
rect 315302 159200 315358 160400
rect 316130 159202 316186 160400
rect 316236 159310 316540 159338
rect 316236 159202 316264 159310
rect 316130 159200 316264 159202
rect 311912 157334 311940 159200
rect 311912 157306 312032 157334
rect 311624 155780 311676 155786
rect 311624 155722 311676 155728
rect 311636 154748 311664 155722
rect 311898 155544 311954 155553
rect 311716 155508 311768 155514
rect 311716 155450 311768 155456
rect 311808 155508 311860 155514
rect 311898 155479 311954 155488
rect 311808 155450 311860 155456
rect 311728 155417 311756 155450
rect 311714 155408 311770 155417
rect 311714 155343 311770 155352
rect 311820 155009 311848 155450
rect 311912 155378 311940 155479
rect 312004 155378 312032 157306
rect 312084 155712 312136 155718
rect 312084 155654 312136 155660
rect 312096 155417 312124 155654
rect 312082 155408 312138 155417
rect 311900 155372 311952 155378
rect 311900 155314 311952 155320
rect 311992 155372 312044 155378
rect 312082 155343 312138 155352
rect 311992 155314 312044 155320
rect 311806 155000 311862 155009
rect 311806 154935 311862 154944
rect 311808 154760 311860 154766
rect 311636 154720 311808 154748
rect 311808 154702 311860 154708
rect 312740 154494 312768 159200
rect 313188 155372 313240 155378
rect 313188 155314 313240 155320
rect 312728 154488 312780 154494
rect 312728 154430 312780 154436
rect 312266 154048 312322 154057
rect 312266 153983 312322 153992
rect 311716 153740 311768 153746
rect 311716 153682 311768 153688
rect 311808 153740 311860 153746
rect 311808 153682 311860 153688
rect 311728 153377 311756 153682
rect 311714 153368 311770 153377
rect 311714 153303 311770 153312
rect 311820 153270 311848 153682
rect 311898 153368 311954 153377
rect 311898 153303 311954 153312
rect 311912 153270 311940 153303
rect 311808 153264 311860 153270
rect 311808 153206 311860 153212
rect 311900 153264 311952 153270
rect 311900 153206 311952 153212
rect 311532 152788 311584 152794
rect 311532 152730 311584 152736
rect 312280 150226 312308 153983
rect 312360 153740 312412 153746
rect 312728 153740 312780 153746
rect 312360 153682 312412 153688
rect 312556 153700 312728 153728
rect 312372 153649 312400 153682
rect 312358 153640 312414 153649
rect 312358 153575 312414 153584
rect 312360 153536 312412 153542
rect 312556 153490 312584 153700
rect 312728 153682 312780 153688
rect 312910 153640 312966 153649
rect 312910 153575 312966 153584
rect 312412 153484 312584 153490
rect 312360 153478 312584 153484
rect 312372 153462 312584 153478
rect 312924 153406 312952 153575
rect 312912 153400 312964 153406
rect 312912 153342 312964 153348
rect 313200 152930 313228 155314
rect 313568 154766 313596 159200
rect 314396 155378 314424 159200
rect 315316 155514 315344 159200
rect 316144 159174 316264 159200
rect 315948 155712 316000 155718
rect 315948 155654 316000 155660
rect 314568 155508 314620 155514
rect 314568 155450 314620 155456
rect 315304 155508 315356 155514
rect 315304 155450 315356 155456
rect 314384 155372 314436 155378
rect 314384 155314 314436 155320
rect 313464 154760 313516 154766
rect 313464 154702 313516 154708
rect 313556 154760 313608 154766
rect 313556 154702 313608 154708
rect 313096 152924 313148 152930
rect 313096 152866 313148 152872
rect 313188 152924 313240 152930
rect 313188 152866 313240 152872
rect 311452 150198 311894 150226
rect 312280 150198 312538 150226
rect 311176 150062 311250 150090
rect 311222 149940 311250 150062
rect 311866 149940 311894 150198
rect 312510 149940 312538 150198
rect 313108 150090 313136 152866
rect 313476 152658 313504 154702
rect 314580 153270 314608 155450
rect 314384 153264 314436 153270
rect 314384 153206 314436 153212
rect 314568 153264 314620 153270
rect 314568 153206 314620 153212
rect 313832 152924 313884 152930
rect 313832 152866 313884 152872
rect 313464 152652 313516 152658
rect 313464 152594 313516 152600
rect 313844 152386 313872 152866
rect 313740 152380 313792 152386
rect 313740 152322 313792 152328
rect 313832 152380 313884 152386
rect 313832 152322 313884 152328
rect 313752 150090 313780 152322
rect 314396 150090 314424 153206
rect 315960 153202 315988 155654
rect 316512 154562 316540 159310
rect 316958 159200 317014 160400
rect 317786 159200 317842 160400
rect 318614 159200 318670 160400
rect 319442 159200 319498 160400
rect 320270 159200 320326 160400
rect 321098 159200 321154 160400
rect 322018 159200 322074 160400
rect 322846 159200 322902 160400
rect 323674 159200 323730 160400
rect 324502 159200 324558 160400
rect 325330 159200 325386 160400
rect 326158 159200 326214 160400
rect 326986 159200 327042 160400
rect 327906 159200 327962 160400
rect 328734 159200 328790 160400
rect 329562 159200 329618 160400
rect 330390 159202 330446 160400
rect 330496 159310 330800 159338
rect 330496 159202 330524 159310
rect 330390 159200 330524 159202
rect 316972 157334 317000 159200
rect 316972 157306 317092 157334
rect 316592 155712 316644 155718
rect 316592 155654 316644 155660
rect 316604 154630 316632 155654
rect 316774 155544 316830 155553
rect 316774 155479 316830 155488
rect 316788 155446 316816 155479
rect 316684 155440 316736 155446
rect 316684 155382 316736 155388
rect 316776 155440 316828 155446
rect 316776 155382 316828 155388
rect 316696 154630 316724 155382
rect 316592 154624 316644 154630
rect 316592 154566 316644 154572
rect 316684 154624 316736 154630
rect 316684 154566 316736 154572
rect 316408 154556 316460 154562
rect 316408 154498 316460 154504
rect 316500 154556 316552 154562
rect 316500 154498 316552 154504
rect 316420 153678 316448 154498
rect 316316 153672 316368 153678
rect 316316 153614 316368 153620
rect 316408 153672 316460 153678
rect 316408 153614 316460 153620
rect 316328 153270 316356 153614
rect 316224 153264 316276 153270
rect 316222 153232 316224 153241
rect 316316 153264 316368 153270
rect 316276 153232 316278 153241
rect 315672 153196 315724 153202
rect 315672 153138 315724 153144
rect 315948 153196 316000 153202
rect 316316 153206 316368 153212
rect 316960 153264 317012 153270
rect 316960 153206 317012 153212
rect 316222 153167 316278 153176
rect 315948 153138 316000 153144
rect 315028 151224 315080 151230
rect 315028 151166 315080 151172
rect 315040 150090 315068 151166
rect 315684 150090 315712 153138
rect 316684 152924 316736 152930
rect 316684 152866 316736 152872
rect 316316 152856 316368 152862
rect 316316 152798 316368 152804
rect 316328 150090 316356 152798
rect 316592 151972 316644 151978
rect 316592 151914 316644 151920
rect 316604 151774 316632 151914
rect 316696 151842 316724 152866
rect 316684 151836 316736 151842
rect 316684 151778 316736 151784
rect 316592 151768 316644 151774
rect 316592 151710 316644 151716
rect 316972 150090 317000 153206
rect 317064 152862 317092 157306
rect 317800 153406 317828 159200
rect 317604 153400 317656 153406
rect 317604 153342 317656 153348
rect 317788 153400 317840 153406
rect 317788 153342 317840 153348
rect 317144 153264 317196 153270
rect 317142 153232 317144 153241
rect 317196 153232 317198 153241
rect 317142 153167 317198 153176
rect 317052 152856 317104 152862
rect 317052 152798 317104 152804
rect 317616 150090 317644 153342
rect 318628 153202 318656 159200
rect 319456 153406 319484 159200
rect 320284 155718 320312 159200
rect 321112 156466 321140 159200
rect 321100 156460 321152 156466
rect 321100 156402 321152 156408
rect 321376 155984 321428 155990
rect 321376 155926 321428 155932
rect 321560 155984 321612 155990
rect 321560 155926 321612 155932
rect 321388 155786 321416 155926
rect 321376 155780 321428 155786
rect 321376 155722 321428 155728
rect 321468 155780 321520 155786
rect 321468 155722 321520 155728
rect 320180 155712 320232 155718
rect 320180 155654 320232 155660
rect 320272 155712 320324 155718
rect 321480 155666 321508 155722
rect 320272 155654 320324 155660
rect 319534 154456 319590 154465
rect 319534 154391 319590 154400
rect 319352 153400 319404 153406
rect 319352 153342 319404 153348
rect 319444 153400 319496 153406
rect 319444 153342 319496 153348
rect 318248 153196 318300 153202
rect 318248 153138 318300 153144
rect 318616 153196 318668 153202
rect 318616 153138 318668 153144
rect 318260 150090 318288 153138
rect 318892 152652 318944 152658
rect 318892 152594 318944 152600
rect 318984 152652 319036 152658
rect 318984 152594 319036 152600
rect 318904 150090 318932 152594
rect 318996 152386 319024 152594
rect 319364 152386 319392 153342
rect 318984 152380 319036 152386
rect 318984 152322 319036 152328
rect 319352 152380 319404 152386
rect 319352 152322 319404 152328
rect 319548 150090 319576 154391
rect 320192 153785 320220 155654
rect 321388 155638 321508 155666
rect 321388 155514 321416 155638
rect 321376 155508 321428 155514
rect 321376 155450 321428 155456
rect 321468 155508 321520 155514
rect 321468 155450 321520 155456
rect 320272 155440 320324 155446
rect 320272 155382 320324 155388
rect 320178 153776 320234 153785
rect 320178 153711 320234 153720
rect 320284 153105 320312 155382
rect 321480 155122 321508 155450
rect 321388 155094 321508 155122
rect 321388 154902 321416 155094
rect 321376 154896 321428 154902
rect 321376 154838 321428 154844
rect 320270 153096 320326 153105
rect 320270 153031 320326 153040
rect 321572 152998 321600 155926
rect 321928 155032 321980 155038
rect 321834 155000 321890 155009
rect 321928 154974 321980 154980
rect 321834 154935 321836 154944
rect 321888 154935 321890 154944
rect 321836 154906 321888 154912
rect 321940 154902 321968 154974
rect 321928 154896 321980 154902
rect 321928 154838 321980 154844
rect 322032 154698 322060 159200
rect 322112 155032 322164 155038
rect 322112 154974 322164 154980
rect 322202 155000 322258 155009
rect 322020 154692 322072 154698
rect 322020 154634 322072 154640
rect 321836 154624 321888 154630
rect 321888 154584 321968 154612
rect 321836 154566 321888 154572
rect 321940 154578 321968 154584
rect 322124 154578 322152 154974
rect 322202 154935 322204 154944
rect 322256 154935 322258 154944
rect 322204 154906 322256 154912
rect 321940 154550 322152 154578
rect 322110 154320 322166 154329
rect 322110 154255 322166 154264
rect 320824 152992 320876 152998
rect 320824 152934 320876 152940
rect 321560 152992 321612 152998
rect 321560 152934 321612 152940
rect 320180 151292 320232 151298
rect 320180 151234 320232 151240
rect 320192 150090 320220 151234
rect 320836 150090 320864 152934
rect 321466 152688 321522 152697
rect 321466 152623 321522 152632
rect 321480 150226 321508 152623
rect 321480 150198 321554 150226
rect 313108 150062 313182 150090
rect 313752 150062 313826 150090
rect 314396 150062 314470 150090
rect 315040 150062 315114 150090
rect 315684 150062 315758 150090
rect 316328 150062 316402 150090
rect 316972 150062 317046 150090
rect 317616 150062 317690 150090
rect 318260 150062 318334 150090
rect 318904 150062 318978 150090
rect 319548 150062 319622 150090
rect 320192 150062 320266 150090
rect 320836 150062 320910 150090
rect 313154 149940 313182 150062
rect 313798 149940 313826 150062
rect 314442 149940 314470 150062
rect 315086 149940 315114 150062
rect 315730 149940 315758 150062
rect 316374 149940 316402 150062
rect 317018 149940 317046 150062
rect 317662 149940 317690 150062
rect 318306 149940 318334 150062
rect 318950 149940 318978 150062
rect 319594 149940 319622 150062
rect 320238 149940 320266 150062
rect 320882 149940 320910 150062
rect 321526 149940 321554 150198
rect 322124 150090 322152 154255
rect 322860 153542 322888 159200
rect 322756 153536 322808 153542
rect 322756 153478 322808 153484
rect 322848 153536 322900 153542
rect 322848 153478 322900 153484
rect 322768 150090 322796 153478
rect 323398 153096 323454 153105
rect 323398 153031 323454 153040
rect 323412 150090 323440 153031
rect 323688 151978 323716 159200
rect 324516 155990 324544 159200
rect 324504 155984 324556 155990
rect 324504 155926 324556 155932
rect 325240 155440 325292 155446
rect 325240 155382 325292 155388
rect 324688 153740 324740 153746
rect 324688 153682 324740 153688
rect 324044 152992 324096 152998
rect 324044 152934 324096 152940
rect 323676 151972 323728 151978
rect 323676 151914 323728 151920
rect 324056 150090 324084 152934
rect 324700 150090 324728 153682
rect 325252 153513 325280 155382
rect 325344 154442 325372 159200
rect 326172 157334 326200 159200
rect 326172 157306 326752 157334
rect 326620 155984 326672 155990
rect 326620 155926 326672 155932
rect 326160 155916 326212 155922
rect 326160 155858 326212 155864
rect 325424 155576 325476 155582
rect 325424 155518 325476 155524
rect 325436 155446 325464 155518
rect 325424 155440 325476 155446
rect 325424 155382 325476 155388
rect 325976 155032 326028 155038
rect 325976 154974 326028 154980
rect 325344 154414 325740 154442
rect 325332 153808 325384 153814
rect 325332 153750 325384 153756
rect 325238 153504 325294 153513
rect 325238 153439 325294 153448
rect 325344 150090 325372 153750
rect 325712 152998 325740 154414
rect 325700 152992 325752 152998
rect 325700 152934 325752 152940
rect 325988 151960 326016 154974
rect 326172 154630 326200 155858
rect 326436 155848 326488 155854
rect 326436 155790 326488 155796
rect 326344 155712 326396 155718
rect 326344 155654 326396 155660
rect 326356 155038 326384 155654
rect 326448 155174 326476 155790
rect 326528 155712 326580 155718
rect 326528 155654 326580 155660
rect 326436 155168 326488 155174
rect 326436 155110 326488 155116
rect 326344 155032 326396 155038
rect 326344 154974 326396 154980
rect 326540 154902 326568 155654
rect 326632 155582 326660 155926
rect 326620 155576 326672 155582
rect 326620 155518 326672 155524
rect 326528 154896 326580 154902
rect 326528 154838 326580 154844
rect 326620 154896 326672 154902
rect 326620 154838 326672 154844
rect 326632 154698 326660 154838
rect 326620 154692 326672 154698
rect 326620 154634 326672 154640
rect 326068 154624 326120 154630
rect 326066 154592 326068 154601
rect 326160 154624 326212 154630
rect 326120 154592 326122 154601
rect 326160 154566 326212 154572
rect 326066 154527 326122 154536
rect 326252 153944 326304 153950
rect 326080 153892 326252 153898
rect 326080 153886 326304 153892
rect 326080 153882 326292 153886
rect 326068 153876 326292 153882
rect 326120 153870 326292 153876
rect 326436 153876 326488 153882
rect 326068 153818 326120 153824
rect 326436 153818 326488 153824
rect 326344 153740 326396 153746
rect 326344 153682 326396 153688
rect 326356 153406 326384 153682
rect 326344 153400 326396 153406
rect 326344 153342 326396 153348
rect 326448 153338 326476 153818
rect 326528 153808 326580 153814
rect 326528 153750 326580 153756
rect 326620 153808 326672 153814
rect 326620 153750 326672 153756
rect 326540 153338 326568 153750
rect 326632 153542 326660 153750
rect 326620 153536 326672 153542
rect 326620 153478 326672 153484
rect 326724 153406 326752 157306
rect 327000 155174 327028 159200
rect 327264 156460 327316 156466
rect 327264 156402 327316 156408
rect 327276 155514 327304 156402
rect 327264 155508 327316 155514
rect 327264 155450 327316 155456
rect 326988 155168 327040 155174
rect 326988 155110 327040 155116
rect 327920 154698 327948 159200
rect 328748 155582 328776 159200
rect 329194 155680 329250 155689
rect 329194 155615 329250 155624
rect 328644 155576 328696 155582
rect 328644 155518 328696 155524
rect 328736 155576 328788 155582
rect 328736 155518 328788 155524
rect 327908 154692 327960 154698
rect 327908 154634 327960 154640
rect 327630 154592 327686 154601
rect 327630 154527 327686 154536
rect 327538 153504 327594 153513
rect 327264 153468 327316 153474
rect 327644 153474 327672 154527
rect 327908 153672 327960 153678
rect 327908 153614 327960 153620
rect 327538 153439 327594 153448
rect 327632 153468 327684 153474
rect 327264 153410 327316 153416
rect 326712 153400 326764 153406
rect 326712 153342 326764 153348
rect 326436 153332 326488 153338
rect 326436 153274 326488 153280
rect 326528 153332 326580 153338
rect 326528 153274 326580 153280
rect 326620 153060 326672 153066
rect 326620 153002 326672 153008
rect 325988 151932 326108 151960
rect 326080 151842 326108 151932
rect 325976 151836 326028 151842
rect 325976 151778 326028 151784
rect 326068 151836 326120 151842
rect 326068 151778 326120 151784
rect 325988 150090 326016 151778
rect 326632 150090 326660 153002
rect 326804 152992 326856 152998
rect 326804 152934 326856 152940
rect 326816 151978 326844 152934
rect 326804 151972 326856 151978
rect 326804 151914 326856 151920
rect 327276 150090 327304 153410
rect 327552 153406 327580 153439
rect 327632 153410 327684 153416
rect 327540 153400 327592 153406
rect 327540 153342 327592 153348
rect 327920 150090 327948 153614
rect 328656 153241 328684 155518
rect 328642 153232 328698 153241
rect 328642 153167 328698 153176
rect 328552 151836 328604 151842
rect 328552 151778 328604 151784
rect 328564 150090 328592 151778
rect 329208 150090 329236 155615
rect 329576 153678 329604 159200
rect 330404 159174 330524 159200
rect 329838 153912 329894 153921
rect 329838 153847 329894 153856
rect 329564 153672 329616 153678
rect 329564 153614 329616 153620
rect 329852 150090 329880 153847
rect 330772 153134 330800 159310
rect 331218 159200 331274 160400
rect 332046 159200 332102 160400
rect 332874 159200 332930 160400
rect 333702 159200 333758 160400
rect 334622 159200 334678 160400
rect 335450 159200 335506 160400
rect 336278 159200 336334 160400
rect 337106 159200 337162 160400
rect 337934 159200 337990 160400
rect 338762 159200 338818 160400
rect 339590 159200 339646 160400
rect 340418 159200 340474 160400
rect 341338 159200 341394 160400
rect 342166 159200 342222 160400
rect 342994 159200 343050 160400
rect 343822 159200 343878 160400
rect 344650 159200 344706 160400
rect 345478 159200 345534 160400
rect 346306 159200 346362 160400
rect 347134 159200 347190 160400
rect 348054 159200 348110 160400
rect 348882 159200 348938 160400
rect 349710 159200 349766 160400
rect 350538 159200 350594 160400
rect 351366 159200 351422 160400
rect 352194 159200 352250 160400
rect 353022 159200 353078 160400
rect 353850 159200 353906 160400
rect 354770 159200 354826 160400
rect 355598 159200 355654 160400
rect 356426 159200 356482 160400
rect 357254 159200 357310 160400
rect 358082 159200 358138 160400
rect 358910 159200 358966 160400
rect 359738 159200 359794 160400
rect 360658 159200 360714 160400
rect 361486 159200 361542 160400
rect 362314 159200 362370 160400
rect 363142 159200 363198 160400
rect 363970 159200 364026 160400
rect 364798 159200 364854 160400
rect 365626 159200 365682 160400
rect 366454 159200 366510 160400
rect 367374 159200 367430 160400
rect 368202 159200 368258 160400
rect 369030 159200 369086 160400
rect 369858 159200 369914 160400
rect 370686 159200 370742 160400
rect 371514 159200 371570 160400
rect 372342 159200 372398 160400
rect 373170 159200 373226 160400
rect 374090 159200 374146 160400
rect 374918 159200 374974 160400
rect 375746 159200 375802 160400
rect 376574 159200 376630 160400
rect 377402 159200 377458 160400
rect 378230 159200 378286 160400
rect 379058 159200 379114 160400
rect 379886 159200 379942 160400
rect 380806 159200 380862 160400
rect 381634 159200 381690 160400
rect 382462 159200 382518 160400
rect 383290 159200 383346 160400
rect 384118 159200 384174 160400
rect 384946 159200 385002 160400
rect 385774 159200 385830 160400
rect 386602 159200 386658 160400
rect 387522 159200 387578 160400
rect 388350 159200 388406 160400
rect 389178 159200 389234 160400
rect 390006 159200 390062 160400
rect 390834 159200 390890 160400
rect 391662 159200 391718 160400
rect 392490 159200 392546 160400
rect 393410 159200 393466 160400
rect 394238 159200 394294 160400
rect 395066 159200 395122 160400
rect 395894 159200 395950 160400
rect 396722 159200 396778 160400
rect 397550 159200 397606 160400
rect 398378 159200 398434 160400
rect 399206 159200 399262 160400
rect 400126 159200 400182 160400
rect 400954 159200 401010 160400
rect 401782 159200 401838 160400
rect 402610 159200 402666 160400
rect 403438 159200 403494 160400
rect 404266 159200 404322 160400
rect 405094 159200 405150 160400
rect 405922 159200 405978 160400
rect 406842 159200 406898 160400
rect 407670 159200 407726 160400
rect 408498 159200 408554 160400
rect 409326 159200 409382 160400
rect 410154 159200 410210 160400
rect 410982 159200 411038 160400
rect 411810 159200 411866 160400
rect 412638 159200 412694 160400
rect 413558 159200 413614 160400
rect 414386 159200 414442 160400
rect 415214 159200 415270 160400
rect 416042 159200 416098 160400
rect 416870 159200 416926 160400
rect 417698 159200 417754 160400
rect 418526 159200 418582 160400
rect 419354 159200 419410 160400
rect 420274 159200 420330 160400
rect 421102 159200 421158 160400
rect 421930 159200 421986 160400
rect 422758 159200 422814 160400
rect 423586 159200 423642 160400
rect 424414 159200 424470 160400
rect 425242 159200 425298 160400
rect 426162 159200 426218 160400
rect 426990 159200 427046 160400
rect 427818 159200 427874 160400
rect 428646 159200 428702 160400
rect 429474 159200 429530 160400
rect 430302 159200 430358 160400
rect 431130 159200 431186 160400
rect 431958 159200 432014 160400
rect 432878 159200 432934 160400
rect 433706 159200 433762 160400
rect 434534 159200 434590 160400
rect 435362 159200 435418 160400
rect 436190 159200 436246 160400
rect 437018 159200 437074 160400
rect 437846 159200 437902 160400
rect 438674 159200 438730 160400
rect 439594 159200 439650 160400
rect 440422 159200 440478 160400
rect 441250 159200 441306 160400
rect 442078 159200 442134 160400
rect 442906 159200 442962 160400
rect 443734 159200 443790 160400
rect 444562 159200 444618 160400
rect 445390 159200 445446 160400
rect 446310 159200 446366 160400
rect 447138 159200 447194 160400
rect 447966 159200 448022 160400
rect 448794 159200 448850 160400
rect 449622 159200 449678 160400
rect 450450 159200 450506 160400
rect 451278 159200 451334 160400
rect 452106 159200 452162 160400
rect 453026 159200 453082 160400
rect 453854 159200 453910 160400
rect 454682 159200 454738 160400
rect 455510 159200 455566 160400
rect 456338 159200 456394 160400
rect 457166 159200 457222 160400
rect 457994 159200 458050 160400
rect 458914 159200 458970 160400
rect 459742 159200 459798 160400
rect 460570 159200 460626 160400
rect 461398 159200 461454 160400
rect 462226 159200 462282 160400
rect 463054 159200 463110 160400
rect 463882 159200 463938 160400
rect 464710 159200 464766 160400
rect 465630 159200 465686 160400
rect 466458 159200 466514 160400
rect 467286 159200 467342 160400
rect 468114 159200 468170 160400
rect 468942 159200 468998 160400
rect 469770 159200 469826 160400
rect 470598 159200 470654 160400
rect 471426 159200 471482 160400
rect 472346 159200 472402 160400
rect 473174 159200 473230 160400
rect 474002 159200 474058 160400
rect 474830 159200 474886 160400
rect 475658 159200 475714 160400
rect 476486 159200 476542 160400
rect 477314 159200 477370 160400
rect 478142 159200 478198 160400
rect 479062 159200 479118 160400
rect 479890 159200 479946 160400
rect 480718 159200 480774 160400
rect 481546 159200 481602 160400
rect 482374 159200 482430 160400
rect 483202 159200 483258 160400
rect 484030 159200 484086 160400
rect 484858 159200 484914 160400
rect 485778 159200 485834 160400
rect 486606 159200 486662 160400
rect 487434 159200 487490 160400
rect 488262 159200 488318 160400
rect 489090 159200 489146 160400
rect 489918 159200 489974 160400
rect 490746 159200 490802 160400
rect 491666 159200 491722 160400
rect 492494 159200 492550 160400
rect 493322 159200 493378 160400
rect 494150 159200 494206 160400
rect 494978 159200 495034 160400
rect 495806 159200 495862 160400
rect 496634 159200 496690 160400
rect 497462 159200 497518 160400
rect 498382 159200 498438 160400
rect 499210 159200 499266 160400
rect 500038 159200 500094 160400
rect 500866 159200 500922 160400
rect 501694 159200 501750 160400
rect 502522 159200 502578 160400
rect 503350 159200 503406 160400
rect 504178 159202 504234 160400
rect 504284 159310 504496 159338
rect 504284 159202 504312 159310
rect 504178 159200 504312 159202
rect 331232 157334 331260 159200
rect 331232 157306 331352 157334
rect 331324 155446 331352 157306
rect 331784 155786 331996 155802
rect 331772 155780 332008 155786
rect 331824 155774 331956 155780
rect 331772 155722 331824 155728
rect 331956 155722 332008 155728
rect 332060 155718 332088 159200
rect 332048 155712 332100 155718
rect 332048 155654 332100 155660
rect 331220 155440 331272 155446
rect 331220 155382 331272 155388
rect 331312 155440 331364 155446
rect 331312 155382 331364 155388
rect 331232 154329 331260 155382
rect 332508 154624 332560 154630
rect 332508 154566 332560 154572
rect 331218 154320 331274 154329
rect 331218 154255 331274 154264
rect 332416 153604 332468 153610
rect 332416 153546 332468 153552
rect 331404 153400 331456 153406
rect 331456 153348 331628 153354
rect 331404 153342 331628 153348
rect 331416 153338 331628 153342
rect 331416 153332 331640 153338
rect 331416 153326 331588 153332
rect 331588 153274 331640 153280
rect 330484 153128 330536 153134
rect 330484 153070 330536 153076
rect 330760 153128 330812 153134
rect 330760 153070 330812 153076
rect 330496 150090 330524 153070
rect 331770 152824 331826 152833
rect 331770 152759 331826 152768
rect 331128 152176 331180 152182
rect 331128 152118 331180 152124
rect 331140 150090 331168 152118
rect 331784 150090 331812 152759
rect 332428 150090 332456 153546
rect 332520 151858 332548 154566
rect 332888 153610 332916 159200
rect 333716 157334 333744 159200
rect 333716 157306 333836 157334
rect 333612 156052 333664 156058
rect 333612 155994 333664 156000
rect 332876 153604 332928 153610
rect 332876 153546 332928 153552
rect 333060 153264 333112 153270
rect 332782 153232 332838 153241
rect 333060 153206 333112 153212
rect 332782 153167 332838 153176
rect 332796 151978 332824 153167
rect 332784 151972 332836 151978
rect 332784 151914 332836 151920
rect 332520 151842 332732 151858
rect 332520 151836 332744 151842
rect 332520 151830 332692 151836
rect 332692 151778 332744 151784
rect 333072 150090 333100 153206
rect 333624 150226 333652 155994
rect 333808 155854 333836 157306
rect 333796 155848 333848 155854
rect 333796 155790 333848 155796
rect 333980 155712 334032 155718
rect 333980 155654 334032 155660
rect 333992 152182 334020 155654
rect 334636 154630 334664 159200
rect 335268 155916 335320 155922
rect 335268 155858 335320 155864
rect 334624 154624 334676 154630
rect 334624 154566 334676 154572
rect 335280 153406 335308 155858
rect 335464 155718 335492 159200
rect 336004 156052 336056 156058
rect 336004 155994 336056 156000
rect 335452 155712 335504 155718
rect 335452 155654 335504 155660
rect 335912 155440 335964 155446
rect 335912 155382 335964 155388
rect 335924 154986 335952 155382
rect 336016 155106 336044 155994
rect 336188 155848 336240 155854
rect 336188 155790 336240 155796
rect 336200 155582 336228 155790
rect 336096 155576 336148 155582
rect 336096 155518 336148 155524
rect 336188 155576 336240 155582
rect 336188 155518 336240 155524
rect 336108 155446 336136 155518
rect 336096 155440 336148 155446
rect 336096 155382 336148 155388
rect 336004 155100 336056 155106
rect 336004 155042 336056 155048
rect 336096 155100 336148 155106
rect 336096 155042 336148 155048
rect 336108 154986 336136 155042
rect 335924 154958 336136 154986
rect 336186 154320 336242 154329
rect 336096 154284 336148 154290
rect 336186 154255 336188 154264
rect 336096 154226 336148 154232
rect 336240 154255 336242 154264
rect 336188 154226 336240 154232
rect 336108 154154 336136 154226
rect 336004 154148 336056 154154
rect 336004 154090 336056 154096
rect 336096 154148 336148 154154
rect 336096 154090 336148 154096
rect 336016 154018 336044 154090
rect 335912 154012 335964 154018
rect 335912 153954 335964 153960
rect 336004 154012 336056 154018
rect 336004 153954 336056 153960
rect 335544 153876 335596 153882
rect 335544 153818 335596 153824
rect 334900 153400 334952 153406
rect 334900 153342 334952 153348
rect 335268 153400 335320 153406
rect 335268 153342 335320 153348
rect 333980 152176 334032 152182
rect 333980 152118 334032 152124
rect 334348 151836 334400 151842
rect 334348 151778 334400 151784
rect 333624 150198 333790 150226
rect 322124 150062 322198 150090
rect 322768 150062 322842 150090
rect 323412 150062 323486 150090
rect 324056 150062 324130 150090
rect 324700 150062 324774 150090
rect 325344 150062 325418 150090
rect 325988 150062 326062 150090
rect 326632 150062 326706 150090
rect 327276 150062 327350 150090
rect 327920 150062 327994 150090
rect 328564 150062 328638 150090
rect 329208 150062 329282 150090
rect 329852 150062 329926 150090
rect 330496 150062 330570 150090
rect 331140 150062 331214 150090
rect 331784 150062 331858 150090
rect 332428 150062 332502 150090
rect 333072 150062 333146 150090
rect 322170 149940 322198 150062
rect 322814 149940 322842 150062
rect 323458 149940 323486 150062
rect 324102 149940 324130 150062
rect 324746 149940 324774 150062
rect 325390 149940 325418 150062
rect 326034 149940 326062 150062
rect 326678 149940 326706 150062
rect 327322 149940 327350 150062
rect 327966 149940 327994 150062
rect 328610 149940 328638 150062
rect 329254 149940 329282 150062
rect 329898 149940 329926 150062
rect 330542 149940 330570 150062
rect 331186 149940 331214 150062
rect 331830 149940 331858 150062
rect 332474 149940 332502 150062
rect 333118 149940 333146 150062
rect 333762 149940 333790 150198
rect 334360 150090 334388 151778
rect 334912 150090 334940 153342
rect 335556 150090 335584 153818
rect 335924 153270 335952 153954
rect 336292 153950 336320 159200
rect 336280 153944 336332 153950
rect 336280 153886 336332 153892
rect 337120 153406 337148 159200
rect 337948 155854 337976 159200
rect 337844 155848 337896 155854
rect 337844 155790 337896 155796
rect 337936 155848 337988 155854
rect 337936 155790 337988 155796
rect 337476 153876 337528 153882
rect 337476 153818 337528 153824
rect 337016 153400 337068 153406
rect 337014 153368 337016 153377
rect 337108 153400 337160 153406
rect 337068 153368 337070 153377
rect 337108 153342 337160 153348
rect 337014 153303 337070 153312
rect 335912 153264 335964 153270
rect 335912 153206 335964 153212
rect 336188 152448 336240 152454
rect 336188 152390 336240 152396
rect 336830 152416 336886 152425
rect 336200 150090 336228 152390
rect 336830 152351 336886 152360
rect 336844 150090 336872 152351
rect 337488 150090 337516 153818
rect 337856 151842 337884 155790
rect 338118 153776 338174 153785
rect 338118 153711 338174 153720
rect 337844 151836 337896 151842
rect 337844 151778 337896 151784
rect 338132 150090 338160 153711
rect 338776 152454 338804 159200
rect 339604 153882 339632 159200
rect 340234 154864 340290 154873
rect 340234 154799 340290 154808
rect 340328 154828 340380 154834
rect 340248 154766 340276 154799
rect 340328 154770 340380 154776
rect 340236 154760 340288 154766
rect 340340 154737 340368 154770
rect 340236 154702 340288 154708
rect 340326 154728 340382 154737
rect 340326 154663 340382 154672
rect 340432 154290 340460 159200
rect 340788 155848 340840 155854
rect 340788 155790 340840 155796
rect 340510 155000 340566 155009
rect 340510 154935 340512 154944
rect 340564 154935 340566 154944
rect 340512 154906 340564 154912
rect 340144 154284 340196 154290
rect 340144 154226 340196 154232
rect 340420 154284 340472 154290
rect 340420 154226 340472 154232
rect 339592 153876 339644 153882
rect 339592 153818 339644 153824
rect 339406 153368 339462 153377
rect 339406 153303 339462 153312
rect 338764 152448 338816 152454
rect 338764 152390 338816 152396
rect 338764 151836 338816 151842
rect 338764 151778 338816 151784
rect 338776 150090 338804 151778
rect 339420 150090 339448 153303
rect 340156 153270 340184 154226
rect 340052 153264 340104 153270
rect 340052 153206 340104 153212
rect 340144 153264 340196 153270
rect 340144 153206 340196 153212
rect 340064 150090 340092 153206
rect 340800 152250 340828 155790
rect 340972 155644 341024 155650
rect 340972 155586 341024 155592
rect 341064 155644 341116 155650
rect 341064 155586 341116 155592
rect 340984 154952 341012 155586
rect 341076 155310 341104 155586
rect 341064 155304 341116 155310
rect 341064 155246 341116 155252
rect 341248 155236 341300 155242
rect 341248 155178 341300 155184
rect 341156 155100 341208 155106
rect 341156 155042 341208 155048
rect 341064 154964 341116 154970
rect 340984 154924 341064 154952
rect 341064 154906 341116 154912
rect 340878 154864 340934 154873
rect 340878 154799 340934 154808
rect 340892 154766 340920 154799
rect 340880 154760 340932 154766
rect 340880 154702 340932 154708
rect 341168 154698 341196 155042
rect 341260 155009 341288 155178
rect 341352 155106 341380 159200
rect 342180 155854 342208 159200
rect 342168 155848 342220 155854
rect 342168 155790 342220 155796
rect 342166 155272 342222 155281
rect 342166 155207 342222 155216
rect 341340 155100 341392 155106
rect 341340 155042 341392 155048
rect 342076 155100 342128 155106
rect 342076 155042 342128 155048
rect 341246 155000 341302 155009
rect 341246 154935 341302 154944
rect 341156 154692 341208 154698
rect 341156 154634 341208 154640
rect 341340 152312 341392 152318
rect 341340 152254 341392 152260
rect 340696 152244 340748 152250
rect 340696 152186 340748 152192
rect 340788 152244 340840 152250
rect 340788 152186 340840 152192
rect 340708 150090 340736 152186
rect 341352 150090 341380 152254
rect 342088 152114 342116 155042
rect 342180 152318 342208 155207
rect 342810 154728 342866 154737
rect 342810 154663 342866 154672
rect 342718 154320 342774 154329
rect 342718 154255 342774 154264
rect 342732 154222 342760 154255
rect 342824 154222 342852 154663
rect 342720 154216 342772 154222
rect 342720 154158 342772 154164
rect 342812 154216 342864 154222
rect 342812 154158 342864 154164
rect 343008 154018 343036 159200
rect 343836 155106 343864 159200
rect 344664 155922 344692 159200
rect 343916 155916 343968 155922
rect 343916 155858 343968 155864
rect 344652 155916 344704 155922
rect 344652 155858 344704 155864
rect 343824 155100 343876 155106
rect 343824 155042 343876 155048
rect 342628 154012 342680 154018
rect 342628 153954 342680 153960
rect 342996 154012 343048 154018
rect 342996 153954 343048 153960
rect 342168 152312 342220 152318
rect 342168 152254 342220 152260
rect 341984 152108 342036 152114
rect 341984 152050 342036 152056
rect 342076 152108 342128 152114
rect 342076 152050 342128 152056
rect 341996 150090 342024 152050
rect 342640 150090 342668 153954
rect 342904 153400 342956 153406
rect 342902 153368 342904 153377
rect 342956 153368 342958 153377
rect 342902 153303 342958 153312
rect 343272 153332 343324 153338
rect 343272 153274 343324 153280
rect 343284 150090 343312 153274
rect 343928 150090 343956 155858
rect 344928 155236 344980 155242
rect 344928 155178 344980 155184
rect 344560 152312 344612 152318
rect 344560 152254 344612 152260
rect 344652 152312 344704 152318
rect 344652 152254 344704 152260
rect 344572 150090 344600 152254
rect 344664 152114 344692 152254
rect 344652 152108 344704 152114
rect 344652 152050 344704 152056
rect 344940 151910 344968 155178
rect 345204 154148 345256 154154
rect 345204 154090 345256 154096
rect 344928 151904 344980 151910
rect 344928 151846 344980 151852
rect 345216 150090 345244 154090
rect 345388 153400 345440 153406
rect 345386 153368 345388 153377
rect 345440 153368 345442 153377
rect 345386 153303 345442 153312
rect 345492 152114 345520 159200
rect 345754 154320 345810 154329
rect 345664 154284 345716 154290
rect 345754 154255 345756 154264
rect 345664 154226 345716 154232
rect 345808 154255 345810 154264
rect 345756 154226 345808 154232
rect 345676 153474 345704 154226
rect 346320 154154 346348 159200
rect 346308 154148 346360 154154
rect 346308 154090 346360 154096
rect 345664 153468 345716 153474
rect 345664 153410 345716 153416
rect 346492 152516 346544 152522
rect 346492 152458 346544 152464
rect 345480 152108 345532 152114
rect 345480 152050 345532 152056
rect 345848 152040 345900 152046
rect 345848 151982 345900 151988
rect 345860 150090 345888 151982
rect 346504 150090 346532 152458
rect 347148 152114 347176 159200
rect 347780 154080 347832 154086
rect 347780 154022 347832 154028
rect 347136 152108 347188 152114
rect 347136 152050 347188 152056
rect 347228 152040 347280 152046
rect 347228 151982 347280 151988
rect 347240 151842 347268 151982
rect 347136 151836 347188 151842
rect 347136 151778 347188 151784
rect 347228 151836 347280 151842
rect 347228 151778 347280 151784
rect 347148 150090 347176 151778
rect 347792 150090 347820 154022
rect 348068 152046 348096 159200
rect 348896 155990 348924 159200
rect 348884 155984 348936 155990
rect 348884 155926 348936 155932
rect 348792 155304 348844 155310
rect 348792 155246 348844 155252
rect 348804 155145 348832 155246
rect 348790 155136 348846 155145
rect 348790 155071 348846 155080
rect 348792 154964 348844 154970
rect 348792 154906 348844 154912
rect 348516 154216 348568 154222
rect 348516 154158 348568 154164
rect 348528 153338 348556 154158
rect 348424 153332 348476 153338
rect 348424 153274 348476 153280
rect 348516 153332 348568 153338
rect 348516 153274 348568 153280
rect 348056 152040 348108 152046
rect 348056 151982 348108 151988
rect 348436 150090 348464 153274
rect 348804 150226 348832 154906
rect 349724 154086 349752 159200
rect 349896 155644 349948 155650
rect 349896 155586 349948 155592
rect 349908 155281 349936 155586
rect 349894 155272 349950 155281
rect 349894 155207 349950 155216
rect 350356 154284 350408 154290
rect 350356 154226 350408 154232
rect 349712 154080 349764 154086
rect 349712 154022 349764 154028
rect 349712 151904 349764 151910
rect 349712 151846 349764 151852
rect 348804 150198 349154 150226
rect 334360 150062 334434 150090
rect 334912 150062 334986 150090
rect 335556 150062 335630 150090
rect 336200 150062 336274 150090
rect 336844 150062 336918 150090
rect 337488 150062 337562 150090
rect 338132 150062 338206 150090
rect 338776 150062 338850 150090
rect 339420 150062 339494 150090
rect 340064 150062 340138 150090
rect 340708 150062 340782 150090
rect 341352 150062 341426 150090
rect 341996 150062 342070 150090
rect 342640 150062 342714 150090
rect 343284 150062 343358 150090
rect 343928 150062 344002 150090
rect 344572 150062 344646 150090
rect 345216 150062 345290 150090
rect 345860 150062 345934 150090
rect 346504 150062 346578 150090
rect 347148 150062 347222 150090
rect 347792 150062 347866 150090
rect 348436 150062 348510 150090
rect 334406 149940 334434 150062
rect 334958 149940 334986 150062
rect 335602 149940 335630 150062
rect 336246 149940 336274 150062
rect 336890 149940 336918 150062
rect 337534 149940 337562 150062
rect 338178 149940 338206 150062
rect 338822 149940 338850 150062
rect 339466 149940 339494 150062
rect 340110 149940 340138 150062
rect 340754 149940 340782 150062
rect 341398 149940 341426 150062
rect 342042 149940 342070 150062
rect 342686 149940 342714 150062
rect 343330 149940 343358 150062
rect 343974 149940 344002 150062
rect 344618 149940 344646 150062
rect 345262 149940 345290 150062
rect 345906 149940 345934 150062
rect 346550 149940 346578 150062
rect 347194 149940 347222 150062
rect 347838 149940 347866 150062
rect 348482 149940 348510 150062
rect 349126 149940 349154 150198
rect 349724 150090 349752 151846
rect 350368 150090 350396 154226
rect 350552 152522 350580 159200
rect 351380 157334 351408 159200
rect 351380 157306 351868 157334
rect 351288 155786 351776 155802
rect 351276 155780 351776 155786
rect 351328 155774 351776 155780
rect 351276 155722 351328 155728
rect 351748 155514 351776 155774
rect 351644 155508 351696 155514
rect 351644 155450 351696 155456
rect 351736 155508 351788 155514
rect 351736 155450 351788 155456
rect 351276 155304 351328 155310
rect 351276 155246 351328 155252
rect 351288 155174 351316 155246
rect 351276 155168 351328 155174
rect 351276 155110 351328 155116
rect 351656 154902 351684 155450
rect 351840 155174 351868 157306
rect 351828 155168 351880 155174
rect 351828 155110 351880 155116
rect 351644 154896 351696 154902
rect 351644 154838 351696 154844
rect 351828 154760 351880 154766
rect 351828 154702 351880 154708
rect 351840 154222 351868 154702
rect 351828 154216 351880 154222
rect 351828 154158 351880 154164
rect 350724 153808 350776 153814
rect 350776 153756 350948 153762
rect 350724 153750 350948 153756
rect 350736 153746 350948 153750
rect 350736 153740 350960 153746
rect 350736 153734 350908 153740
rect 350908 153682 350960 153688
rect 351644 152924 351696 152930
rect 351644 152866 351696 152872
rect 351000 152720 351052 152726
rect 351000 152662 351052 152668
rect 350540 152516 350592 152522
rect 350540 152458 350592 152464
rect 351012 150090 351040 152662
rect 351656 150090 351684 152866
rect 352208 152726 352236 159200
rect 353036 157334 353064 159200
rect 353036 157306 353156 157334
rect 352840 154352 352892 154358
rect 352840 154294 352892 154300
rect 352196 152720 352248 152726
rect 352196 152662 352248 152668
rect 352288 152584 352340 152590
rect 352288 152526 352340 152532
rect 352300 150090 352328 152526
rect 352852 150226 352880 154294
rect 353128 154222 353156 157306
rect 353864 154766 353892 159200
rect 354586 155272 354642 155281
rect 354586 155207 354642 155216
rect 354218 155136 354274 155145
rect 354218 155071 354274 155080
rect 353852 154760 353904 154766
rect 353852 154702 353904 154708
rect 353116 154216 353168 154222
rect 353116 154158 353168 154164
rect 353576 153264 353628 153270
rect 353576 153206 353628 153212
rect 352852 150198 353018 150226
rect 349724 150062 349798 150090
rect 350368 150062 350442 150090
rect 351012 150062 351086 150090
rect 351656 150062 351730 150090
rect 352300 150062 352374 150090
rect 349770 149940 349798 150062
rect 350414 149940 350442 150062
rect 351058 149940 351086 150062
rect 351702 149940 351730 150062
rect 352346 149940 352374 150062
rect 352990 149940 353018 150198
rect 353588 150090 353616 153206
rect 354232 150090 354260 155071
rect 354600 151858 354628 155207
rect 354784 152930 354812 159200
rect 355232 155780 355284 155786
rect 355232 155722 355284 155728
rect 355244 155514 355272 155722
rect 355232 155508 355284 155514
rect 355232 155450 355284 155456
rect 355324 155508 355376 155514
rect 355324 155450 355376 155456
rect 355232 155032 355284 155038
rect 355232 154974 355284 154980
rect 355244 153270 355272 154974
rect 355336 154970 355364 155450
rect 355416 155304 355468 155310
rect 355416 155246 355468 155252
rect 355428 155038 355456 155246
rect 355612 155242 355640 159200
rect 355600 155236 355652 155242
rect 355600 155178 355652 155184
rect 355416 155032 355468 155038
rect 355416 154974 355468 154980
rect 355324 154964 355376 154970
rect 355324 154906 355376 154912
rect 355508 154420 355560 154426
rect 355508 154362 355560 154368
rect 355324 154284 355376 154290
rect 355324 154226 355376 154232
rect 355336 153746 355364 154226
rect 355324 153740 355376 153746
rect 355324 153682 355376 153688
rect 355232 153264 355284 153270
rect 355232 153206 355284 153212
rect 354772 152924 354824 152930
rect 354772 152866 354824 152872
rect 355232 152516 355284 152522
rect 355232 152458 355284 152464
rect 355244 152114 355272 152458
rect 355232 152108 355284 152114
rect 355232 152050 355284 152056
rect 355324 152108 355376 152114
rect 355324 152050 355376 152056
rect 354600 151830 354904 151858
rect 355336 151842 355364 152050
rect 354876 150226 354904 151830
rect 355324 151836 355376 151842
rect 355324 151778 355376 151784
rect 354876 150198 354950 150226
rect 353588 150062 353662 150090
rect 354232 150062 354306 150090
rect 353634 149940 353662 150062
rect 354278 149940 354306 150062
rect 354922 149940 354950 150198
rect 355520 150090 355548 154362
rect 356152 153332 356204 153338
rect 356152 153274 356204 153280
rect 356164 150090 356192 153274
rect 356440 153270 356468 159200
rect 356520 155984 356572 155990
rect 356520 155926 356572 155932
rect 356532 155650 356560 155926
rect 356520 155644 356572 155650
rect 356520 155586 356572 155592
rect 357268 154970 357296 159200
rect 358096 155786 358124 159200
rect 357992 155780 358044 155786
rect 357992 155722 358044 155728
rect 358084 155780 358136 155786
rect 358084 155722 358136 155728
rect 357440 155032 357492 155038
rect 357440 154974 357492 154980
rect 357256 154964 357308 154970
rect 357256 154906 357308 154912
rect 357452 153746 357480 154974
rect 357440 153740 357492 153746
rect 357440 153682 357492 153688
rect 356428 153264 356480 153270
rect 356428 153206 356480 153212
rect 356796 152788 356848 152794
rect 356796 152730 356848 152736
rect 356888 152788 356940 152794
rect 356888 152730 356940 152736
rect 356808 150090 356836 152730
rect 356900 152590 356928 152730
rect 358004 152658 358032 155722
rect 358452 155304 358504 155310
rect 358452 155246 358504 155252
rect 358084 154488 358136 154494
rect 358084 154430 358136 154436
rect 357440 152652 357492 152658
rect 357440 152594 357492 152600
rect 357992 152652 358044 152658
rect 357992 152594 358044 152600
rect 356888 152584 356940 152590
rect 356888 152526 356940 152532
rect 357452 150090 357480 152594
rect 358096 150090 358124 154430
rect 358464 154426 358492 155246
rect 358452 154420 358504 154426
rect 358452 154362 358504 154368
rect 358728 154352 358780 154358
rect 358728 154294 358780 154300
rect 358740 150090 358768 154294
rect 358924 151842 358952 159200
rect 359372 154420 359424 154426
rect 359372 154362 359424 154368
rect 358912 151836 358964 151842
rect 358912 151778 358964 151784
rect 359384 150090 359412 154362
rect 359752 154358 359780 159200
rect 360672 157334 360700 159200
rect 360672 157306 360792 157334
rect 360660 154556 360712 154562
rect 360660 154498 360712 154504
rect 359740 154352 359792 154358
rect 359740 154294 359792 154300
rect 360016 152652 360068 152658
rect 360016 152594 360068 152600
rect 360028 150090 360056 152594
rect 360672 150090 360700 154498
rect 360764 152794 360792 157306
rect 361304 152856 361356 152862
rect 361304 152798 361356 152804
rect 360752 152788 360804 152794
rect 360752 152730 360804 152736
rect 361316 150090 361344 152798
rect 361500 152658 361528 159200
rect 362328 155378 362356 159200
rect 362684 155508 362736 155514
rect 362684 155450 362736 155456
rect 362316 155372 362368 155378
rect 362316 155314 362368 155320
rect 362592 153196 362644 153202
rect 362592 153138 362644 153144
rect 361488 152652 361540 152658
rect 361488 152594 361540 152600
rect 361948 152380 362000 152386
rect 361948 152322 362000 152328
rect 361960 150090 361988 152322
rect 362604 150090 362632 153138
rect 362696 152386 362724 155450
rect 363156 154494 363184 159200
rect 363984 154834 364012 159200
rect 364812 155786 364840 159200
rect 364708 155780 364760 155786
rect 364708 155722 364760 155728
rect 364800 155780 364852 155786
rect 364800 155722 364852 155728
rect 364720 155310 364748 155722
rect 365352 155712 365404 155718
rect 365088 155650 365300 155666
rect 365352 155654 365404 155660
rect 365076 155644 365312 155650
rect 365128 155638 365260 155644
rect 365076 155586 365128 155592
rect 365260 155586 365312 155592
rect 365364 155582 365392 155654
rect 364984 155576 365036 155582
rect 364984 155518 365036 155524
rect 365352 155576 365404 155582
rect 365352 155518 365404 155524
rect 364708 155304 364760 155310
rect 364708 155246 364760 155252
rect 364996 154902 365024 155518
rect 364248 154896 364300 154902
rect 364248 154838 364300 154844
rect 364984 154896 365036 154902
rect 364984 154838 365036 154844
rect 363880 154828 363932 154834
rect 363880 154770 363932 154776
rect 363972 154828 364024 154834
rect 363972 154770 364024 154776
rect 363892 154562 363920 154770
rect 363880 154556 363932 154562
rect 363880 154498 363932 154504
rect 363144 154488 363196 154494
rect 363144 154430 363196 154436
rect 363236 153808 363288 153814
rect 363236 153750 363288 153756
rect 362684 152380 362736 152386
rect 362684 152322 362736 152328
rect 363248 150090 363276 153750
rect 363880 153332 363932 153338
rect 363880 153274 363932 153280
rect 363892 150090 363920 153274
rect 364260 153218 364288 154838
rect 364892 153536 364944 153542
rect 364892 153478 364944 153484
rect 364904 153338 364932 153478
rect 364996 153474 365208 153490
rect 364984 153468 365220 153474
rect 365036 153462 365168 153468
rect 364984 153410 365036 153416
rect 365168 153410 365220 153416
rect 364892 153332 364944 153338
rect 364892 153274 364944 153280
rect 364260 153190 364564 153218
rect 365640 153202 365668 159200
rect 366468 154426 366496 159200
rect 367388 154698 367416 159200
rect 367100 154692 367152 154698
rect 367100 154634 367152 154640
rect 367376 154692 367428 154698
rect 367376 154634 367428 154640
rect 366456 154420 366508 154426
rect 366456 154362 366508 154368
rect 365720 154284 365772 154290
rect 365720 154226 365772 154232
rect 364536 150226 364564 153190
rect 365628 153196 365680 153202
rect 365628 153138 365680 153144
rect 365168 152380 365220 152386
rect 365168 152322 365220 152328
rect 364536 150198 364610 150226
rect 355520 150062 355594 150090
rect 356164 150062 356238 150090
rect 356808 150062 356882 150090
rect 357452 150062 357526 150090
rect 358096 150062 358170 150090
rect 358740 150062 358814 150090
rect 359384 150062 359458 150090
rect 360028 150062 360102 150090
rect 360672 150062 360746 150090
rect 361316 150062 361390 150090
rect 361960 150062 362034 150090
rect 362604 150062 362678 150090
rect 363248 150062 363322 150090
rect 363892 150062 363966 150090
rect 355566 149940 355594 150062
rect 356210 149940 356238 150062
rect 356854 149940 356882 150062
rect 357498 149940 357526 150062
rect 358142 149940 358170 150062
rect 358786 149940 358814 150062
rect 359430 149940 359458 150062
rect 360074 149940 360102 150062
rect 360718 149940 360746 150062
rect 361362 149940 361390 150062
rect 362006 149940 362034 150062
rect 362650 149940 362678 150062
rect 363294 149940 363322 150062
rect 363938 149940 363966 150062
rect 364582 149940 364610 150198
rect 365180 150090 365208 152322
rect 365732 150090 365760 154226
rect 367112 153814 367140 154634
rect 367100 153808 367152 153814
rect 367100 153750 367152 153756
rect 367652 153060 367704 153066
rect 367652 153002 367704 153008
rect 366364 152992 366416 152998
rect 366364 152934 366416 152940
rect 366376 150090 366404 152934
rect 367008 151972 367060 151978
rect 367008 151914 367060 151920
rect 367020 150090 367048 151914
rect 367664 150090 367692 153002
rect 368216 152862 368244 159200
rect 369044 155514 369072 159200
rect 369032 155508 369084 155514
rect 369032 155450 369084 155456
rect 368480 154624 368532 154630
rect 368480 154566 368532 154572
rect 368492 153406 368520 154566
rect 369872 154562 369900 159200
rect 370228 155440 370280 155446
rect 370228 155382 370280 155388
rect 369584 154556 369636 154562
rect 369584 154498 369636 154504
rect 369860 154556 369912 154562
rect 369860 154498 369912 154504
rect 368940 153740 368992 153746
rect 368940 153682 368992 153688
rect 368480 153400 368532 153406
rect 368480 153342 368532 153348
rect 368296 153332 368348 153338
rect 368296 153274 368348 153280
rect 368204 152856 368256 152862
rect 368204 152798 368256 152804
rect 368308 150090 368336 153274
rect 368952 150090 368980 153682
rect 369596 150090 369624 154498
rect 370240 150226 370268 155382
rect 370700 153066 370728 159200
rect 371528 155038 371556 159200
rect 371516 155032 371568 155038
rect 371516 154974 371568 154980
rect 372160 153808 372212 153814
rect 372160 153750 372212 153756
rect 370872 153672 370924 153678
rect 370872 153614 370924 153620
rect 370688 153060 370740 153066
rect 370688 153002 370740 153008
rect 370884 150226 370912 153614
rect 371516 153128 371568 153134
rect 371516 153070 371568 153076
rect 371528 150226 371556 153070
rect 372172 150226 372200 153750
rect 372356 152998 372384 159200
rect 373184 153814 373212 159200
rect 374000 154896 374052 154902
rect 374000 154838 374052 154844
rect 373172 153808 373224 153814
rect 373172 153750 373224 153756
rect 373448 153604 373500 153610
rect 373448 153546 373500 153552
rect 372344 152992 372396 152998
rect 372344 152934 372396 152940
rect 372804 152176 372856 152182
rect 372804 152118 372856 152124
rect 372816 150226 372844 152118
rect 373460 150226 373488 153546
rect 374012 151814 374040 154838
rect 374104 154630 374132 159200
rect 374932 154902 374960 159200
rect 375472 155576 375524 155582
rect 375472 155518 375524 155524
rect 374920 154896 374972 154902
rect 374920 154838 374972 154844
rect 374092 154624 374144 154630
rect 374092 154566 374144 154572
rect 374736 153400 374788 153406
rect 374736 153342 374788 153348
rect 374012 151786 374132 151814
rect 374104 150226 374132 151786
rect 374748 150226 374776 153342
rect 375484 150226 375512 155518
rect 375760 155446 375788 159200
rect 375748 155440 375800 155446
rect 375748 155382 375800 155388
rect 376588 153950 376616 159200
rect 377220 155100 377272 155106
rect 377220 155042 377272 155048
rect 376024 153944 376076 153950
rect 376024 153886 376076 153892
rect 376576 153944 376628 153950
rect 376576 153886 376628 153892
rect 370240 150198 370314 150226
rect 370884 150198 370958 150226
rect 371528 150198 371602 150226
rect 372172 150198 372246 150226
rect 372816 150198 372890 150226
rect 373460 150198 373534 150226
rect 374104 150198 374178 150226
rect 374748 150198 374822 150226
rect 365180 150062 365254 150090
rect 365732 150062 365806 150090
rect 366376 150062 366450 150090
rect 367020 150062 367094 150090
rect 367664 150062 367738 150090
rect 368308 150062 368382 150090
rect 368952 150062 369026 150090
rect 369596 150062 369670 150090
rect 365226 149940 365254 150062
rect 365778 149940 365806 150062
rect 366422 149940 366450 150062
rect 367066 149940 367094 150062
rect 367710 149940 367738 150062
rect 368354 149940 368382 150062
rect 368998 149940 369026 150062
rect 369642 149940 369670 150062
rect 370286 149940 370314 150198
rect 370930 149940 370958 150198
rect 371574 149940 371602 150198
rect 372218 149940 372246 150198
rect 372862 149940 372890 150198
rect 373506 149940 373534 150198
rect 374150 149940 374178 150198
rect 374794 149940 374822 150198
rect 375438 150198 375512 150226
rect 376036 150226 376064 153886
rect 376668 153536 376720 153542
rect 376668 153478 376720 153484
rect 376680 150226 376708 153478
rect 377232 152386 377260 155042
rect 377416 153134 377444 159200
rect 377404 153128 377456 153134
rect 377404 153070 377456 153076
rect 378244 152454 378272 159200
rect 379072 155582 379100 159200
rect 379060 155576 379112 155582
rect 379060 155518 379112 155524
rect 379900 153882 379928 159200
rect 380532 155848 380584 155854
rect 380532 155790 380584 155796
rect 378600 153876 378652 153882
rect 378600 153818 378652 153824
rect 379888 153876 379940 153882
rect 379888 153818 379940 153824
rect 377956 152448 378008 152454
rect 377956 152390 378008 152396
rect 378232 152448 378284 152454
rect 378232 152390 378284 152396
rect 377220 152380 377272 152386
rect 377220 152322 377272 152328
rect 377312 152244 377364 152250
rect 377312 152186 377364 152192
rect 377324 150226 377352 152186
rect 377968 150226 377996 152390
rect 378612 150226 378640 153818
rect 379244 153468 379296 153474
rect 379244 153410 379296 153416
rect 379256 150226 379284 153410
rect 379888 152312 379940 152318
rect 379888 152254 379940 152260
rect 379900 150226 379928 152254
rect 380544 150226 380572 155790
rect 380820 155106 380848 159200
rect 381648 155854 381676 159200
rect 382372 155916 382424 155922
rect 382372 155858 382424 155864
rect 381636 155848 381688 155854
rect 381636 155790 381688 155796
rect 380808 155100 380860 155106
rect 380808 155042 380860 155048
rect 380992 154964 381044 154970
rect 380992 154906 381044 154912
rect 380900 154760 380952 154766
rect 380900 154702 380952 154708
rect 380912 152250 380940 154702
rect 381004 152318 381032 154906
rect 381176 154012 381228 154018
rect 381176 153954 381228 153960
rect 380992 152312 381044 152318
rect 380992 152254 381044 152260
rect 380900 152244 380952 152250
rect 380900 152186 380952 152192
rect 381188 150226 381216 153954
rect 381820 152380 381872 152386
rect 381820 152322 381872 152328
rect 381832 150226 381860 152322
rect 382384 151814 382412 155858
rect 382476 155718 382504 159200
rect 382464 155712 382516 155718
rect 382464 155654 382516 155660
rect 383304 154018 383332 159200
rect 383752 154148 383804 154154
rect 383752 154090 383804 154096
rect 383292 154012 383344 154018
rect 383292 153954 383344 153960
rect 383108 152108 383160 152114
rect 383108 152050 383160 152056
rect 382384 151786 382504 151814
rect 382476 150226 382504 151786
rect 383120 150226 383148 152050
rect 383764 150226 383792 154090
rect 384132 152386 384160 159200
rect 384580 155780 384632 155786
rect 384580 155722 384632 155728
rect 384592 155106 384620 155722
rect 384488 155100 384540 155106
rect 384488 155042 384540 155048
rect 384580 155100 384632 155106
rect 384580 155042 384632 155048
rect 384500 154986 384528 155042
rect 384500 154970 384712 154986
rect 384500 154964 384724 154970
rect 384500 154958 384672 154964
rect 384672 154906 384724 154912
rect 384960 152522 384988 159200
rect 385592 155644 385644 155650
rect 385592 155586 385644 155592
rect 384396 152516 384448 152522
rect 384396 152458 384448 152464
rect 384948 152516 385000 152522
rect 384948 152458 385000 152464
rect 384120 152380 384172 152386
rect 384120 152322 384172 152328
rect 384408 150226 384436 152458
rect 385040 152040 385092 152046
rect 385040 151982 385092 151988
rect 385052 150226 385080 151982
rect 385604 151814 385632 155586
rect 385788 154766 385816 159200
rect 386236 154828 386288 154834
rect 386236 154770 386288 154776
rect 385684 154760 385736 154766
rect 385684 154702 385736 154708
rect 385776 154760 385828 154766
rect 385776 154702 385828 154708
rect 385696 152046 385724 154702
rect 385684 152040 385736 152046
rect 385684 151982 385736 151988
rect 386248 151978 386276 154770
rect 386616 154154 386644 159200
rect 387536 154698 387564 159200
rect 388364 155786 388392 159200
rect 388352 155780 388404 155786
rect 388352 155722 388404 155728
rect 387616 155168 387668 155174
rect 387616 155110 387668 155116
rect 387524 154692 387576 154698
rect 387524 154634 387576 154640
rect 386604 154148 386656 154154
rect 386604 154090 386656 154096
rect 386328 154080 386380 154086
rect 386328 154022 386380 154028
rect 386236 151972 386288 151978
rect 386236 151914 386288 151920
rect 385604 151786 385724 151814
rect 385696 150226 385724 151786
rect 386340 150226 386368 154022
rect 386972 152720 387024 152726
rect 386972 152662 387024 152668
rect 386984 150226 387012 152662
rect 387628 150226 387656 155110
rect 388536 154964 388588 154970
rect 388536 154906 388588 154912
rect 388444 154624 388496 154630
rect 388444 154566 388496 154572
rect 388260 152584 388312 152590
rect 388260 152526 388312 152532
rect 388272 150226 388300 152526
rect 388456 152114 388484 154566
rect 388548 152182 388576 154906
rect 388904 154216 388956 154222
rect 388904 154158 388956 154164
rect 388536 152176 388588 152182
rect 388536 152118 388588 152124
rect 388444 152108 388496 152114
rect 388444 152050 388496 152056
rect 388916 150226 388944 154158
rect 389192 152726 389220 159200
rect 390020 154086 390048 159200
rect 390744 155236 390796 155242
rect 390744 155178 390796 155184
rect 390008 154080 390060 154086
rect 390008 154022 390060 154028
rect 390192 152924 390244 152930
rect 390192 152866 390244 152872
rect 389180 152720 389232 152726
rect 389180 152662 389232 152668
rect 389548 152244 389600 152250
rect 389548 152186 389600 152192
rect 389560 150226 389588 152186
rect 390204 150226 390232 152866
rect 390756 151814 390784 155178
rect 390848 154630 390876 159200
rect 391676 155174 391704 159200
rect 392400 155304 392452 155310
rect 392400 155246 392452 155252
rect 391664 155168 391716 155174
rect 391664 155110 391716 155116
rect 390928 154692 390980 154698
rect 390928 154634 390980 154640
rect 390836 154624 390888 154630
rect 390836 154566 390888 154572
rect 390940 152250 390968 154634
rect 392308 154624 392360 154630
rect 392308 154566 392360 154572
rect 391480 153264 391532 153270
rect 391480 153206 391532 153212
rect 390928 152244 390980 152250
rect 390928 152186 390980 152192
rect 390756 151786 390876 151814
rect 390848 150226 390876 151786
rect 391492 150226 391520 153206
rect 392320 152318 392348 154566
rect 392124 152312 392176 152318
rect 392124 152254 392176 152260
rect 392308 152312 392360 152318
rect 392308 152254 392360 152260
rect 392136 150226 392164 152254
rect 392412 151814 392440 155246
rect 392504 154970 392532 159200
rect 392492 154964 392544 154970
rect 392492 154906 392544 154912
rect 393424 154290 393452 159200
rect 394056 154352 394108 154358
rect 394056 154294 394108 154300
rect 393412 154284 393464 154290
rect 393412 154226 393464 154232
rect 393412 151904 393464 151910
rect 393412 151846 393464 151852
rect 392412 151786 392808 151814
rect 392780 150226 392808 151786
rect 393424 150226 393452 151846
rect 394068 150226 394096 154294
rect 394252 152930 394280 159200
rect 394884 155372 394936 155378
rect 394884 155314 394936 155320
rect 394240 152924 394292 152930
rect 394240 152866 394292 152872
rect 394700 152788 394752 152794
rect 394700 152730 394752 152736
rect 394712 150226 394740 152730
rect 376036 150198 376110 150226
rect 376680 150198 376754 150226
rect 377324 150198 377398 150226
rect 377968 150198 378042 150226
rect 378612 150198 378686 150226
rect 379256 150198 379330 150226
rect 379900 150198 379974 150226
rect 380544 150198 380618 150226
rect 381188 150198 381262 150226
rect 381832 150198 381906 150226
rect 382476 150198 382550 150226
rect 383120 150198 383194 150226
rect 383764 150198 383838 150226
rect 384408 150198 384482 150226
rect 385052 150198 385126 150226
rect 385696 150198 385770 150226
rect 386340 150198 386414 150226
rect 386984 150198 387058 150226
rect 387628 150198 387702 150226
rect 388272 150198 388346 150226
rect 388916 150198 388990 150226
rect 389560 150198 389634 150226
rect 390204 150198 390278 150226
rect 390848 150198 390922 150226
rect 391492 150198 391566 150226
rect 392136 150198 392210 150226
rect 392780 150198 392854 150226
rect 393424 150198 393498 150226
rect 394068 150198 394142 150226
rect 394712 150198 394786 150226
rect 394896 150210 394924 155314
rect 395080 155310 395108 159200
rect 395068 155304 395120 155310
rect 395068 155246 395120 155252
rect 395436 155100 395488 155106
rect 395436 155042 395488 155048
rect 395448 152658 395476 155042
rect 395344 152652 395396 152658
rect 395344 152594 395396 152600
rect 395436 152652 395488 152658
rect 395436 152594 395488 152600
rect 395356 150226 395384 152594
rect 395908 152590 395936 159200
rect 396448 155032 396500 155038
rect 396448 154974 396500 154980
rect 395896 152584 395948 152590
rect 395896 152526 395948 152532
rect 396460 151910 396488 154974
rect 396540 154488 396592 154494
rect 396540 154430 396592 154436
rect 396448 151904 396500 151910
rect 396448 151846 396500 151852
rect 396552 150226 396580 154430
rect 396736 154222 396764 159200
rect 396724 154216 396776 154222
rect 396724 154158 396776 154164
rect 397564 152794 397592 159200
rect 398392 155650 398420 159200
rect 398840 155848 398892 155854
rect 398840 155790 398892 155796
rect 398380 155644 398432 155650
rect 398380 155586 398432 155592
rect 398104 154896 398156 154902
rect 398104 154838 398156 154844
rect 397552 152788 397604 152794
rect 397552 152730 397604 152736
rect 397828 152652 397880 152658
rect 397828 152594 397880 152600
rect 397184 151972 397236 151978
rect 397184 151914 397236 151920
rect 397196 150226 397224 151914
rect 397840 150226 397868 152594
rect 398116 151978 398144 154838
rect 398472 153196 398524 153202
rect 398472 153138 398524 153144
rect 398104 151972 398156 151978
rect 398104 151914 398156 151920
rect 398484 150226 398512 153138
rect 398852 151842 398880 155790
rect 399220 155786 399248 159200
rect 399208 155780 399260 155786
rect 399208 155722 399260 155728
rect 399116 154420 399168 154426
rect 399116 154362 399168 154368
rect 398840 151836 398892 151842
rect 398840 151778 398892 151784
rect 399128 150226 399156 154362
rect 400140 154358 400168 159200
rect 400968 154426 400996 159200
rect 401796 155854 401824 159200
rect 402244 155916 402296 155922
rect 402244 155858 402296 155864
rect 401784 155848 401836 155854
rect 401784 155790 401836 155796
rect 401048 155508 401100 155514
rect 401048 155450 401100 155456
rect 400956 154420 401008 154426
rect 400956 154362 401008 154368
rect 400128 154352 400180 154358
rect 400128 154294 400180 154300
rect 400404 152856 400456 152862
rect 400404 152798 400456 152804
rect 399760 152040 399812 152046
rect 399760 151982 399812 151988
rect 399772 150226 399800 151982
rect 400416 150226 400444 152798
rect 401060 150226 401088 155450
rect 401692 154556 401744 154562
rect 401692 154498 401744 154504
rect 401704 150226 401732 154498
rect 402256 151842 402284 155858
rect 402336 153060 402388 153066
rect 402336 153002 402388 153008
rect 402244 151836 402296 151842
rect 402244 151778 402296 151784
rect 402348 150226 402376 153002
rect 402624 152658 402652 159200
rect 403452 154494 403480 159200
rect 404280 155242 404308 159200
rect 405108 155718 405136 159200
rect 405096 155712 405148 155718
rect 405096 155654 405148 155660
rect 404912 155644 404964 155650
rect 404912 155586 404964 155592
rect 404924 155530 404952 155586
rect 404924 155502 405044 155530
rect 405936 155514 405964 159200
rect 404268 155236 404320 155242
rect 404268 155178 404320 155184
rect 404176 155168 404228 155174
rect 404176 155110 404228 155116
rect 403440 154488 403492 154494
rect 403440 154430 403492 154436
rect 404188 153202 404216 155110
rect 404268 153808 404320 153814
rect 404268 153750 404320 153756
rect 404176 153196 404228 153202
rect 404176 153138 404228 153144
rect 403624 152992 403676 152998
rect 403624 152934 403676 152940
rect 402612 152652 402664 152658
rect 402612 152594 402664 152600
rect 402980 151904 403032 151910
rect 402980 151846 403032 151852
rect 402992 150226 403020 151846
rect 403636 150226 403664 152934
rect 404280 150226 404308 153750
rect 405016 152114 405044 155502
rect 405924 155508 405976 155514
rect 405924 155450 405976 155456
rect 406200 155440 406252 155446
rect 406200 155382 406252 155388
rect 405648 155304 405700 155310
rect 405648 155246 405700 155252
rect 404912 152108 404964 152114
rect 404912 152050 404964 152056
rect 405004 152108 405056 152114
rect 405004 152050 405056 152056
rect 404924 150226 404952 152050
rect 405660 151978 405688 155246
rect 405556 151972 405608 151978
rect 405556 151914 405608 151920
rect 405648 151972 405700 151978
rect 405648 151914 405700 151920
rect 405568 150226 405596 151914
rect 406212 150226 406240 155382
rect 406856 155378 406884 159200
rect 407304 155848 407356 155854
rect 407304 155790 407356 155796
rect 406844 155372 406896 155378
rect 406844 155314 406896 155320
rect 406844 153944 406896 153950
rect 406844 153886 406896 153892
rect 406856 150226 406884 153886
rect 407316 152046 407344 155790
rect 407684 153950 407712 159200
rect 408512 155106 408540 159200
rect 408868 155712 408920 155718
rect 408868 155654 408920 155660
rect 408776 155576 408828 155582
rect 408776 155518 408828 155524
rect 408500 155100 408552 155106
rect 408500 155042 408552 155048
rect 407672 153944 407724 153950
rect 407672 153886 407724 153892
rect 407488 153128 407540 153134
rect 407488 153070 407540 153076
rect 407304 152040 407356 152046
rect 407304 151982 407356 151988
rect 407500 150226 407528 153070
rect 408132 152448 408184 152454
rect 408132 152390 408184 152396
rect 408144 150226 408172 152390
rect 408788 150226 408816 155518
rect 408880 152454 408908 155654
rect 409340 152862 409368 159200
rect 410168 155582 410196 159200
rect 410156 155576 410208 155582
rect 410156 155518 410208 155524
rect 409420 153876 409472 153882
rect 409420 153818 409472 153824
rect 409328 152856 409380 152862
rect 409328 152798 409380 152804
rect 408868 152448 408920 152454
rect 408868 152390 408920 152396
rect 409432 150226 409460 153818
rect 410996 152998 411024 159200
rect 411824 155922 411852 159200
rect 411812 155916 411864 155922
rect 411812 155858 411864 155864
rect 412652 155650 412680 159200
rect 411352 155644 411404 155650
rect 411352 155586 411404 155592
rect 412640 155644 412692 155650
rect 412640 155586 412692 155592
rect 410984 152992 411036 152998
rect 410984 152934 411036 152940
rect 410064 152176 410116 152182
rect 410064 152118 410116 152124
rect 410076 150226 410104 152118
rect 410708 151836 410760 151842
rect 410708 151778 410760 151784
rect 410720 150226 410748 151778
rect 411364 150226 411392 155586
rect 413572 155446 413600 159200
rect 413928 155916 413980 155922
rect 413928 155858 413980 155864
rect 413560 155440 413612 155446
rect 413560 155382 413612 155388
rect 411720 155100 411772 155106
rect 411720 155042 411772 155048
rect 411732 152182 411760 155042
rect 413192 154760 413244 154766
rect 413192 154702 413244 154708
rect 411996 154012 412048 154018
rect 411996 153954 412048 153960
rect 411720 152176 411772 152182
rect 411720 152118 411772 152124
rect 412008 150226 412036 153954
rect 413100 152516 413152 152522
rect 413100 152458 413152 152464
rect 412640 152380 412692 152386
rect 412640 152322 412692 152328
rect 412652 150226 412680 152322
rect 413112 150498 413140 152458
rect 413204 151814 413232 154702
rect 413940 153066 413968 155858
rect 414400 153134 414428 159200
rect 414572 154148 414624 154154
rect 414572 154090 414624 154096
rect 414388 153128 414440 153134
rect 414388 153070 414440 153076
rect 413928 153060 413980 153066
rect 413928 153002 413980 153008
rect 413204 151786 413968 151814
rect 413112 150470 413324 150498
rect 413296 150226 413324 150470
rect 413940 150226 413968 151786
rect 414584 150226 414612 154090
rect 415228 152522 415256 159200
rect 416056 155174 416084 159200
rect 416688 155780 416740 155786
rect 416688 155722 416740 155728
rect 416044 155168 416096 155174
rect 416044 155110 416096 155116
rect 415492 154964 415544 154970
rect 415492 154906 415544 154912
rect 415216 152516 415268 152522
rect 415216 152458 415268 152464
rect 415504 152386 415532 154906
rect 416504 152720 416556 152726
rect 416504 152662 416556 152668
rect 415492 152380 415544 152386
rect 415492 152322 415544 152328
rect 415216 152244 415268 152250
rect 415216 152186 415268 152192
rect 415228 150226 415256 152186
rect 415860 151904 415912 151910
rect 415860 151846 415912 151852
rect 415872 150226 415900 151846
rect 416516 150226 416544 152662
rect 416700 151842 416728 155722
rect 416884 153882 416912 159200
rect 417424 155576 417476 155582
rect 417424 155518 417476 155524
rect 417436 154154 417464 155518
rect 417424 154148 417476 154154
rect 417424 154090 417476 154096
rect 417148 154080 417200 154086
rect 417148 154022 417200 154028
rect 416872 153876 416924 153882
rect 416872 153818 416924 153824
rect 416688 151836 416740 151842
rect 416688 151778 416740 151784
rect 417160 150226 417188 154022
rect 417712 152726 417740 159200
rect 418540 153202 418568 159200
rect 419368 155854 419396 159200
rect 419356 155848 419408 155854
rect 419356 155790 419408 155796
rect 420184 155644 420236 155650
rect 420184 155586 420236 155592
rect 419172 155508 419224 155514
rect 419172 155450 419224 155456
rect 418436 153196 418488 153202
rect 418436 153138 418488 153144
rect 418528 153196 418580 153202
rect 418528 153138 418580 153144
rect 417700 152720 417752 152726
rect 417700 152662 417752 152668
rect 417792 152312 417844 152318
rect 417792 152254 417844 152260
rect 417804 150226 417832 152254
rect 418448 150226 418476 153138
rect 419184 152386 419212 155450
rect 419724 154284 419776 154290
rect 419724 154226 419776 154232
rect 419080 152380 419132 152386
rect 419080 152322 419132 152328
rect 419172 152380 419224 152386
rect 419172 152322 419224 152328
rect 419092 150226 419120 152322
rect 419736 150226 419764 154226
rect 420196 151910 420224 155586
rect 420288 155310 420316 159200
rect 421116 155582 421144 159200
rect 421104 155576 421156 155582
rect 421104 155518 421156 155524
rect 420276 155304 420328 155310
rect 420276 155246 420328 155252
rect 421944 152930 421972 159200
rect 422772 155378 422800 159200
rect 423220 155848 423272 155854
rect 423220 155790 423272 155796
rect 422668 155372 422720 155378
rect 422668 155314 422720 155320
rect 422760 155372 422812 155378
rect 422760 155314 422812 155320
rect 422680 155174 422708 155314
rect 422576 155168 422628 155174
rect 422576 155110 422628 155116
rect 422668 155168 422720 155174
rect 422668 155110 422720 155116
rect 422300 154216 422352 154222
rect 422300 154158 422352 154164
rect 420368 152924 420420 152930
rect 420368 152866 420420 152872
rect 421932 152924 421984 152930
rect 421932 152866 421984 152872
rect 420184 151904 420236 151910
rect 420184 151846 420236 151852
rect 420380 150226 420408 152866
rect 421656 152584 421708 152590
rect 421656 152526 421708 152532
rect 421012 151972 421064 151978
rect 421012 151914 421064 151920
rect 421024 150226 421052 151914
rect 421668 150226 421696 152526
rect 422312 150226 422340 154158
rect 422588 151978 422616 155110
rect 422944 152788 422996 152794
rect 422944 152730 422996 152736
rect 422576 151972 422628 151978
rect 422576 151914 422628 151920
rect 422956 150226 422984 152730
rect 423232 152250 423260 155790
rect 423600 154018 423628 159200
rect 424428 155786 424456 159200
rect 424416 155780 424468 155786
rect 424416 155722 424468 155728
rect 424968 155372 425020 155378
rect 424968 155314 425020 155320
rect 424876 154352 424928 154358
rect 424876 154294 424928 154300
rect 423588 154012 423640 154018
rect 423588 153954 423640 153960
rect 423220 152244 423272 152250
rect 423220 152186 423272 152192
rect 423588 152108 423640 152114
rect 423588 152050 423640 152056
rect 423600 150226 423628 152050
rect 424232 151836 424284 151842
rect 424232 151778 424284 151784
rect 424244 150226 424272 151778
rect 424888 150226 424916 154294
rect 424980 152794 425008 155314
rect 424968 152788 425020 152794
rect 424968 152730 425020 152736
rect 425256 152250 425284 159200
rect 425520 154420 425572 154426
rect 425520 154362 425572 154368
rect 425244 152244 425296 152250
rect 425244 152186 425296 152192
rect 425532 150226 425560 154362
rect 426176 152590 426204 159200
rect 427004 155514 427032 159200
rect 426992 155508 427044 155514
rect 426992 155450 427044 155456
rect 427728 155236 427780 155242
rect 427728 155178 427780 155184
rect 427360 154488 427412 154494
rect 427360 154430 427412 154436
rect 426808 152652 426860 152658
rect 426808 152594 426860 152600
rect 426164 152584 426216 152590
rect 426164 152526 426216 152532
rect 426164 152040 426216 152046
rect 426164 151982 426216 151988
rect 426176 150226 426204 151982
rect 426820 150226 426848 152594
rect 427372 150226 427400 154430
rect 427740 153898 427768 155178
rect 427832 154086 427860 159200
rect 427820 154080 427872 154086
rect 427820 154022 427872 154028
rect 427740 153870 427860 153898
rect 427832 151814 427860 153870
rect 428660 152538 428688 159200
rect 428660 152510 428780 152538
rect 428752 152454 428780 152510
rect 428648 152448 428700 152454
rect 428648 152390 428700 152396
rect 428740 152448 428792 152454
rect 428740 152390 428792 152396
rect 427832 151786 428044 151814
rect 428016 150226 428044 151786
rect 428660 150226 428688 152390
rect 429488 152386 429516 159200
rect 429936 155168 429988 155174
rect 429936 155110 429988 155116
rect 429292 152380 429344 152386
rect 429292 152322 429344 152328
rect 429476 152380 429528 152386
rect 429476 152322 429528 152328
rect 429304 150226 429332 152322
rect 429948 150226 429976 155110
rect 430316 152658 430344 159200
rect 430580 155576 430632 155582
rect 430580 155518 430632 155524
rect 430592 153950 430620 155518
rect 430488 153944 430540 153950
rect 430488 153886 430540 153892
rect 430580 153944 430632 153950
rect 430580 153886 430632 153892
rect 430500 153762 430528 153886
rect 430500 153734 430712 153762
rect 430580 152856 430632 152862
rect 430580 152798 430632 152804
rect 430304 152652 430356 152658
rect 430304 152594 430356 152600
rect 430592 152046 430620 152798
rect 430580 152040 430632 152046
rect 430580 151982 430632 151988
rect 430684 150226 430712 153734
rect 431144 152862 431172 159200
rect 431972 155582 432000 159200
rect 431960 155576 432012 155582
rect 431960 155518 432012 155524
rect 432512 154148 432564 154154
rect 432512 154090 432564 154096
rect 431132 152856 431184 152862
rect 431132 152798 431184 152804
rect 431224 152312 431276 152318
rect 431224 152254 431276 152260
rect 375438 149940 375466 150198
rect 376082 149940 376110 150198
rect 376726 149940 376754 150198
rect 377370 149940 377398 150198
rect 378014 149940 378042 150198
rect 378658 149940 378686 150198
rect 379302 149940 379330 150198
rect 379946 149940 379974 150198
rect 380590 149940 380618 150198
rect 381234 149940 381262 150198
rect 381878 149940 381906 150198
rect 382522 149940 382550 150198
rect 383166 149940 383194 150198
rect 383810 149940 383838 150198
rect 384454 149940 384482 150198
rect 385098 149940 385126 150198
rect 385742 149940 385770 150198
rect 386386 149940 386414 150198
rect 387030 149940 387058 150198
rect 387674 149940 387702 150198
rect 388318 149940 388346 150198
rect 388962 149940 388990 150198
rect 389606 149940 389634 150198
rect 390250 149940 390278 150198
rect 390894 149940 390922 150198
rect 391538 149940 391566 150198
rect 392182 149940 392210 150198
rect 392826 149940 392854 150198
rect 393470 149940 393498 150198
rect 394114 149940 394142 150198
rect 394758 149940 394786 150198
rect 394884 150204 394936 150210
rect 395356 150198 395430 150226
rect 394884 150146 394936 150152
rect 395402 149940 395430 150198
rect 396034 150204 396086 150210
rect 396552 150198 396626 150226
rect 397196 150198 397270 150226
rect 397840 150198 397914 150226
rect 398484 150198 398558 150226
rect 399128 150198 399202 150226
rect 399772 150198 399846 150226
rect 400416 150198 400490 150226
rect 401060 150198 401134 150226
rect 401704 150198 401778 150226
rect 402348 150198 402422 150226
rect 402992 150198 403066 150226
rect 403636 150198 403710 150226
rect 404280 150198 404354 150226
rect 404924 150198 404998 150226
rect 405568 150198 405642 150226
rect 406212 150198 406286 150226
rect 406856 150198 406930 150226
rect 407500 150198 407574 150226
rect 408144 150198 408218 150226
rect 408788 150198 408862 150226
rect 409432 150198 409506 150226
rect 410076 150198 410150 150226
rect 410720 150198 410794 150226
rect 411364 150198 411438 150226
rect 412008 150198 412082 150226
rect 412652 150198 412726 150226
rect 413296 150198 413370 150226
rect 413940 150198 414014 150226
rect 414584 150198 414658 150226
rect 415228 150198 415302 150226
rect 415872 150198 415946 150226
rect 416516 150198 416590 150226
rect 417160 150198 417234 150226
rect 417804 150198 417878 150226
rect 418448 150198 418522 150226
rect 419092 150198 419166 150226
rect 419736 150198 419810 150226
rect 420380 150198 420454 150226
rect 421024 150198 421098 150226
rect 421668 150198 421742 150226
rect 422312 150198 422386 150226
rect 422956 150198 423030 150226
rect 423600 150198 423674 150226
rect 424244 150198 424318 150226
rect 424888 150198 424962 150226
rect 425532 150198 425606 150226
rect 426176 150198 426250 150226
rect 426820 150198 426894 150226
rect 427372 150198 427446 150226
rect 428016 150198 428090 150226
rect 428660 150198 428734 150226
rect 429304 150198 429378 150226
rect 429948 150198 430022 150226
rect 396034 150146 396086 150152
rect 396046 149940 396074 150146
rect 396598 149940 396626 150198
rect 397242 149940 397270 150198
rect 397886 149940 397914 150198
rect 398530 149940 398558 150198
rect 399174 149940 399202 150198
rect 399818 149940 399846 150198
rect 400462 149940 400490 150198
rect 401106 149940 401134 150198
rect 401750 149940 401778 150198
rect 402394 149940 402422 150198
rect 403038 149940 403066 150198
rect 403682 149940 403710 150198
rect 404326 149940 404354 150198
rect 404970 149940 404998 150198
rect 405614 149940 405642 150198
rect 406258 149940 406286 150198
rect 406902 149940 406930 150198
rect 407546 149940 407574 150198
rect 408190 149940 408218 150198
rect 408834 149940 408862 150198
rect 409478 149940 409506 150198
rect 410122 149940 410150 150198
rect 410766 149940 410794 150198
rect 411410 149940 411438 150198
rect 412054 149940 412082 150198
rect 412698 149940 412726 150198
rect 413342 149940 413370 150198
rect 413986 149940 414014 150198
rect 414630 149940 414658 150198
rect 415274 149940 415302 150198
rect 415918 149940 415946 150198
rect 416562 149940 416590 150198
rect 417206 149940 417234 150198
rect 417850 149940 417878 150198
rect 418494 149940 418522 150198
rect 419138 149940 419166 150198
rect 419782 149940 419810 150198
rect 420426 149940 420454 150198
rect 421070 149940 421098 150198
rect 421714 149940 421742 150198
rect 422358 149940 422386 150198
rect 423002 149940 423030 150198
rect 423646 149940 423674 150198
rect 424290 149940 424318 150198
rect 424934 149940 424962 150198
rect 425578 149940 425606 150198
rect 426222 149940 426250 150198
rect 426866 149940 426894 150198
rect 427418 149940 427446 150198
rect 428062 149940 428090 150198
rect 428706 149940 428734 150198
rect 429350 149940 429378 150198
rect 429994 149940 430022 150198
rect 430638 150198 430712 150226
rect 431236 150226 431264 152254
rect 431776 152040 431828 152046
rect 431776 151982 431828 151988
rect 431788 151814 431816 151982
rect 431788 151786 431908 151814
rect 431880 150226 431908 151786
rect 432524 150226 432552 154090
rect 432892 152425 432920 159200
rect 433720 155718 433748 159200
rect 433708 155712 433760 155718
rect 433708 155654 433760 155660
rect 434548 155242 434576 159200
rect 435376 155650 435404 159200
rect 435364 155644 435416 155650
rect 435364 155586 435416 155592
rect 435088 155440 435140 155446
rect 435088 155382 435140 155388
rect 434536 155236 434588 155242
rect 434536 155178 434588 155184
rect 433800 153060 433852 153066
rect 433800 153002 433852 153008
rect 433156 152992 433208 152998
rect 433156 152934 433208 152940
rect 432878 152416 432934 152425
rect 432878 152351 432934 152360
rect 433168 150226 433196 152934
rect 433812 150226 433840 153002
rect 434444 151904 434496 151910
rect 434444 151846 434496 151852
rect 434456 150226 434484 151846
rect 435100 150226 435128 155382
rect 436204 155106 436232 159200
rect 437032 155378 437060 159200
rect 437480 155780 437532 155786
rect 437480 155722 437532 155728
rect 437020 155372 437072 155378
rect 437020 155314 437072 155320
rect 436192 155100 436244 155106
rect 436192 155042 436244 155048
rect 437492 153270 437520 155722
rect 437860 155174 437888 159200
rect 438688 155446 438716 159200
rect 439608 155786 439636 159200
rect 439596 155780 439648 155786
rect 439596 155722 439648 155728
rect 438676 155440 438728 155446
rect 438676 155382 438728 155388
rect 440240 155304 440292 155310
rect 440240 155246 440292 155252
rect 437848 155168 437900 155174
rect 437848 155110 437900 155116
rect 437664 153876 437716 153882
rect 437664 153818 437716 153824
rect 437480 153264 437532 153270
rect 437480 153206 437532 153212
rect 435732 153128 435784 153134
rect 435732 153070 435784 153076
rect 435744 150226 435772 153070
rect 436376 152516 436428 152522
rect 436376 152458 436428 152464
rect 436388 150226 436416 152458
rect 437020 151972 437072 151978
rect 437020 151914 437072 151920
rect 437032 150226 437060 151914
rect 437676 150226 437704 153818
rect 438952 153196 439004 153202
rect 438952 153138 439004 153144
rect 438308 152720 438360 152726
rect 438308 152662 438360 152668
rect 438320 150226 438348 152662
rect 438964 150226 438992 153138
rect 439596 152176 439648 152182
rect 439596 152118 439648 152124
rect 439608 150226 439636 152118
rect 440252 150226 440280 155246
rect 440436 154970 440464 159200
rect 441264 155038 441292 159200
rect 442092 155854 442120 159200
rect 442080 155848 442132 155854
rect 442080 155790 442132 155796
rect 442920 155310 442948 159200
rect 443748 155922 443776 159200
rect 443736 155916 443788 155922
rect 443736 155858 443788 155864
rect 442908 155304 442960 155310
rect 442908 155246 442960 155252
rect 441252 155032 441304 155038
rect 441252 154974 441304 154980
rect 440424 154964 440476 154970
rect 440424 154906 440476 154912
rect 444576 154834 444604 159200
rect 445208 155576 445260 155582
rect 445208 155518 445260 155524
rect 445116 155508 445168 155514
rect 445116 155450 445168 155456
rect 444564 154828 444616 154834
rect 444564 154770 444616 154776
rect 442816 154012 442868 154018
rect 442816 153954 442868 153960
rect 440884 153944 440936 153950
rect 440884 153886 440936 153892
rect 440896 150226 440924 153886
rect 441528 152924 441580 152930
rect 441528 152866 441580 152872
rect 441540 150226 441568 152866
rect 442172 152788 442224 152794
rect 442172 152730 442224 152736
rect 442184 150226 442212 152730
rect 442828 150226 442856 153954
rect 443460 153264 443512 153270
rect 443460 153206 443512 153212
rect 443472 150226 443500 153206
rect 444748 152584 444800 152590
rect 444748 152526 444800 152532
rect 444104 152312 444156 152318
rect 444104 152254 444156 152260
rect 444116 150226 444144 152254
rect 444760 150226 444788 152526
rect 445128 151814 445156 155450
rect 445220 154698 445248 155518
rect 445404 154766 445432 159200
rect 446324 154902 446352 159200
rect 446404 155644 446456 155650
rect 446404 155586 446456 155592
rect 446416 155446 446444 155586
rect 446404 155440 446456 155446
rect 446404 155382 446456 155388
rect 446312 154896 446364 154902
rect 446312 154838 446364 154844
rect 445392 154760 445444 154766
rect 445392 154702 445444 154708
rect 445208 154692 445260 154698
rect 445208 154634 445260 154640
rect 447152 154630 447180 159200
rect 447980 155514 448008 159200
rect 448612 155712 448664 155718
rect 448612 155654 448664 155660
rect 447968 155508 448020 155514
rect 447968 155450 448020 155456
rect 448520 155236 448572 155242
rect 448520 155178 448572 155184
rect 447232 154692 447284 154698
rect 447232 154634 447284 154640
rect 447140 154624 447192 154630
rect 447140 154566 447192 154572
rect 446036 154080 446088 154086
rect 446036 154022 446088 154028
rect 445128 151786 445432 151814
rect 445404 150226 445432 151786
rect 446048 150226 446076 154022
rect 447244 153134 447272 154634
rect 448532 153202 448560 155178
rect 448520 153196 448572 153202
rect 448520 153138 448572 153144
rect 447232 153128 447284 153134
rect 447232 153070 447284 153076
rect 448624 153066 448652 155654
rect 448808 154698 448836 159200
rect 449636 155582 449664 159200
rect 449624 155576 449676 155582
rect 449624 155518 449676 155524
rect 450464 155446 450492 159200
rect 451292 155530 451320 159200
rect 452120 155650 452148 159200
rect 452844 155712 452896 155718
rect 452844 155654 452896 155660
rect 452108 155644 452160 155650
rect 452108 155586 452160 155592
rect 451292 155502 451504 155530
rect 449992 155440 450044 155446
rect 449992 155382 450044 155388
rect 450452 155440 450504 155446
rect 450452 155382 450504 155388
rect 448796 154692 448848 154698
rect 448796 154634 448848 154640
rect 449256 153128 449308 153134
rect 449256 153070 449308 153076
rect 448612 153060 448664 153066
rect 448612 153002 448664 153008
rect 448612 152856 448664 152862
rect 448612 152798 448664 152804
rect 447968 152652 448020 152658
rect 447968 152594 448020 152600
rect 446680 152448 446732 152454
rect 446680 152390 446732 152396
rect 446692 150226 446720 152390
rect 447324 152380 447376 152386
rect 447324 152322 447376 152328
rect 447336 150226 447364 152322
rect 447980 150226 448008 152594
rect 448624 150226 448652 152798
rect 449268 150226 449296 153070
rect 449898 152416 449954 152425
rect 449898 152351 449954 152360
rect 449912 150226 449940 152351
rect 450004 151910 450032 155382
rect 451280 155372 451332 155378
rect 451280 155314 451332 155320
rect 451292 153202 451320 155314
rect 451476 155106 451504 155502
rect 451372 155100 451424 155106
rect 451372 155042 451424 155048
rect 451464 155100 451516 155106
rect 451464 155042 451516 155048
rect 451188 153196 451240 153202
rect 451188 153138 451240 153144
rect 451280 153196 451332 153202
rect 451280 153138 451332 153144
rect 450636 153060 450688 153066
rect 450636 153002 450688 153008
rect 449992 151904 450044 151910
rect 449992 151846 450044 151852
rect 450648 150226 450676 153002
rect 431236 150198 431310 150226
rect 431880 150198 431954 150226
rect 432524 150198 432598 150226
rect 433168 150198 433242 150226
rect 433812 150198 433886 150226
rect 434456 150198 434530 150226
rect 435100 150198 435174 150226
rect 435744 150198 435818 150226
rect 436388 150198 436462 150226
rect 437032 150198 437106 150226
rect 437676 150198 437750 150226
rect 438320 150198 438394 150226
rect 438964 150198 439038 150226
rect 439608 150198 439682 150226
rect 440252 150198 440326 150226
rect 440896 150198 440970 150226
rect 441540 150198 441614 150226
rect 442184 150198 442258 150226
rect 442828 150198 442902 150226
rect 443472 150198 443546 150226
rect 444116 150198 444190 150226
rect 444760 150198 444834 150226
rect 445404 150198 445478 150226
rect 446048 150198 446122 150226
rect 446692 150198 446766 150226
rect 447336 150198 447410 150226
rect 447980 150198 448054 150226
rect 448624 150198 448698 150226
rect 449268 150198 449342 150226
rect 449912 150198 449986 150226
rect 430638 149940 430666 150198
rect 431282 149940 431310 150198
rect 431926 149940 431954 150198
rect 432570 149940 432598 150198
rect 433214 149940 433242 150198
rect 433858 149940 433886 150198
rect 434502 149940 434530 150198
rect 435146 149940 435174 150198
rect 435790 149940 435818 150198
rect 436434 149940 436462 150198
rect 437078 149940 437106 150198
rect 437722 149940 437750 150198
rect 438366 149940 438394 150198
rect 439010 149940 439038 150198
rect 439654 149940 439682 150198
rect 440298 149940 440326 150198
rect 440942 149940 440970 150198
rect 441586 149940 441614 150198
rect 442230 149940 442258 150198
rect 442874 149940 442902 150198
rect 443518 149940 443546 150198
rect 444162 149940 444190 150198
rect 444806 149940 444834 150198
rect 445450 149940 445478 150198
rect 446094 149940 446122 150198
rect 446738 149940 446766 150198
rect 447382 149940 447410 150198
rect 448026 149940 448054 150198
rect 448670 149940 448698 150198
rect 449314 149940 449342 150198
rect 449958 149940 449986 150198
rect 450602 150198 450676 150226
rect 451200 150226 451228 153138
rect 451200 150198 451274 150226
rect 451384 150210 451412 155042
rect 452856 153134 452884 155654
rect 453040 155394 453068 159200
rect 453868 155718 453896 159200
rect 453856 155712 453908 155718
rect 453856 155654 453908 155660
rect 454696 155446 454724 159200
rect 455052 155780 455104 155786
rect 455052 155722 455104 155728
rect 454592 155440 454644 155446
rect 453040 155378 453160 155394
rect 454592 155382 454644 155388
rect 454684 155440 454736 155446
rect 454684 155382 454736 155388
rect 453040 155372 453172 155378
rect 453040 155366 453120 155372
rect 453120 155314 453172 155320
rect 454604 155242 454632 155382
rect 454592 155236 454644 155242
rect 454592 155178 454644 155184
rect 453212 155168 453264 155174
rect 453212 155110 453264 155116
rect 453120 153196 453172 153202
rect 453120 153138 453172 153144
rect 452844 153128 452896 153134
rect 452844 153070 452896 153076
rect 451832 151904 451884 151910
rect 451832 151846 451884 151852
rect 451844 150226 451872 151846
rect 453132 150226 453160 153138
rect 453224 151814 453252 155110
rect 454408 153128 454460 153134
rect 454408 153070 454460 153076
rect 453224 151786 453804 151814
rect 453776 150226 453804 151786
rect 454420 150226 454448 153070
rect 455064 150226 455092 155722
rect 455524 155038 455552 159200
rect 456352 155786 456380 159200
rect 456984 155848 457036 155854
rect 456984 155790 457036 155796
rect 456340 155780 456392 155786
rect 456340 155722 456392 155728
rect 456800 155304 456852 155310
rect 456800 155246 456852 155252
rect 455420 155032 455472 155038
rect 455420 154974 455472 154980
rect 455512 155032 455564 155038
rect 455512 154974 455564 154980
rect 450602 149940 450630 150198
rect 451246 149940 451274 150198
rect 451372 150204 451424 150210
rect 451844 150198 451918 150226
rect 451372 150146 451424 150152
rect 451890 149940 451918 150198
rect 452522 150204 452574 150210
rect 453132 150198 453206 150226
rect 453776 150198 453850 150226
rect 454420 150198 454494 150226
rect 455064 150198 455138 150226
rect 455432 150210 455460 154974
rect 455696 154964 455748 154970
rect 455696 154906 455748 154912
rect 455708 150226 455736 154906
rect 452522 150146 452574 150152
rect 452534 149940 452562 150146
rect 453178 149940 453206 150198
rect 453822 149940 453850 150198
rect 454466 149940 454494 150198
rect 455110 149940 455138 150198
rect 455420 150204 455472 150210
rect 455708 150198 455782 150226
rect 456812 150210 456840 155246
rect 456996 150226 457024 155790
rect 457180 155038 457208 159200
rect 458008 155174 458036 159200
rect 458272 155916 458324 155922
rect 458272 155858 458324 155864
rect 457996 155168 458048 155174
rect 457996 155110 458048 155116
rect 457168 155032 457220 155038
rect 457168 154974 457220 154980
rect 458180 154624 458232 154630
rect 458180 154566 458232 154572
rect 458192 153202 458220 154566
rect 458180 153196 458232 153202
rect 458180 153138 458232 153144
rect 458284 150226 458312 155858
rect 458928 155854 458956 159200
rect 458916 155848 458968 155854
rect 458916 155790 458968 155796
rect 459652 154896 459704 154902
rect 459652 154838 459704 154844
rect 458364 154828 458416 154834
rect 458364 154770 458416 154776
rect 458376 151814 458404 154770
rect 458732 154760 458784 154766
rect 458732 154702 458784 154708
rect 458744 151814 458772 154702
rect 459560 154692 459612 154698
rect 459560 154634 459612 154640
rect 459572 151910 459600 154634
rect 459560 151904 459612 151910
rect 459560 151846 459612 151852
rect 459664 151814 459692 154838
rect 459756 154630 459784 159200
rect 460584 155922 460612 159200
rect 460572 155916 460624 155922
rect 460572 155858 460624 155864
rect 461412 155666 461440 159200
rect 461412 155638 461532 155666
rect 461400 155508 461452 155514
rect 461400 155450 461452 155456
rect 459744 154624 459796 154630
rect 459744 154566 459796 154572
rect 460756 153196 460808 153202
rect 460756 153138 460808 153144
rect 458376 151786 458680 151814
rect 458744 151786 459508 151814
rect 459664 151786 460152 151814
rect 455420 150146 455472 150152
rect 455754 149940 455782 150198
rect 456386 150204 456438 150210
rect 456386 150146 456438 150152
rect 456800 150204 456852 150210
rect 456996 150198 457070 150226
rect 456800 150146 456852 150152
rect 456398 149940 456426 150146
rect 457042 149940 457070 150198
rect 457674 150204 457726 150210
rect 457674 150146 457726 150152
rect 458238 150198 458312 150226
rect 458652 150226 458680 151786
rect 459480 150226 459508 151786
rect 460124 150226 460152 151786
rect 460768 150226 460796 153138
rect 461412 150226 461440 155450
rect 461504 154766 461532 155638
rect 462240 155310 462268 159200
rect 462688 155576 462740 155582
rect 462688 155518 462740 155524
rect 462228 155304 462280 155310
rect 462228 155246 462280 155252
rect 462320 155236 462372 155242
rect 462320 155178 462372 155184
rect 461492 154760 461544 154766
rect 461492 154702 461544 154708
rect 462044 151904 462096 151910
rect 462044 151846 462096 151852
rect 462056 150226 462084 151846
rect 458652 150198 458910 150226
rect 459480 150198 459554 150226
rect 460124 150198 460198 150226
rect 460768 150198 460842 150226
rect 461412 150198 461486 150226
rect 462056 150198 462130 150226
rect 462332 150210 462360 155178
rect 462700 150226 462728 155518
rect 463068 154834 463096 159200
rect 463896 155650 463924 159200
rect 464344 155780 464396 155786
rect 464344 155722 464396 155728
rect 463884 155644 463936 155650
rect 463884 155586 463936 155592
rect 464356 155514 464384 155722
rect 464724 155582 464752 159200
rect 465540 155712 465592 155718
rect 465540 155654 465592 155660
rect 464620 155576 464672 155582
rect 464620 155518 464672 155524
rect 464712 155576 464764 155582
rect 464712 155518 464764 155524
rect 464344 155508 464396 155514
rect 464344 155450 464396 155456
rect 463700 155100 463752 155106
rect 463700 155042 463752 155048
rect 463056 154828 463108 154834
rect 463056 154770 463108 154776
rect 463712 151814 463740 155042
rect 463712 151786 464016 151814
rect 463988 150226 464016 151786
rect 464632 150226 464660 155518
rect 465080 155372 465132 155378
rect 465080 155314 465132 155320
rect 465092 151814 465120 155314
rect 465552 151814 465580 155654
rect 465644 155378 465672 159200
rect 466472 155854 466500 159200
rect 466460 155848 466512 155854
rect 466460 155790 466512 155796
rect 466368 155440 466420 155446
rect 466368 155382 466420 155388
rect 465632 155372 465684 155378
rect 465632 155314 465684 155320
rect 466380 151814 466408 155382
rect 467300 155242 467328 159200
rect 468128 155718 468156 159200
rect 468116 155712 468168 155718
rect 468116 155654 468168 155660
rect 467748 155508 467800 155514
rect 467748 155450 467800 155456
rect 467288 155236 467340 155242
rect 467288 155178 467340 155184
rect 467012 154964 467064 154970
rect 467012 154906 467064 154912
rect 467024 151814 467052 154906
rect 467760 151814 467788 155450
rect 468956 155446 468984 159200
rect 469784 155786 469812 159200
rect 470508 155916 470560 155922
rect 470508 155858 470560 155864
rect 469312 155780 469364 155786
rect 469312 155722 469364 155728
rect 469772 155780 469824 155786
rect 469772 155722 469824 155728
rect 468944 155440 468996 155446
rect 468944 155382 468996 155388
rect 468024 155168 468076 155174
rect 468024 155110 468076 155116
rect 465092 151786 465304 151814
rect 465552 151786 465948 151814
rect 466380 151786 466592 151814
rect 467024 151786 467236 151814
rect 467760 151786 467880 151814
rect 465276 150226 465304 151786
rect 465920 150226 465948 151786
rect 466564 150226 466592 151786
rect 467208 150226 467236 151786
rect 467852 150226 467880 151786
rect 457686 149940 457714 150146
rect 458238 149940 458266 150198
rect 458882 149940 458910 150198
rect 459526 149940 459554 150198
rect 460170 149940 460198 150198
rect 460814 149940 460842 150198
rect 461458 149940 461486 150198
rect 462102 149940 462130 150198
rect 462320 150204 462372 150210
rect 462700 150198 462774 150226
rect 462320 150146 462372 150152
rect 462746 149940 462774 150198
rect 463378 150204 463430 150210
rect 463988 150198 464062 150226
rect 464632 150198 464706 150226
rect 465276 150198 465350 150226
rect 465920 150198 465994 150226
rect 466564 150198 466638 150226
rect 467208 150198 467282 150226
rect 467852 150198 467926 150226
rect 468036 150210 468064 155110
rect 468484 155032 468536 155038
rect 468484 154974 468536 154980
rect 468496 150226 468524 154974
rect 469324 151814 469352 155722
rect 470520 155394 470548 155858
rect 470612 155530 470640 159200
rect 471440 155922 471468 159200
rect 471428 155916 471480 155922
rect 471428 155858 471480 155864
rect 470612 155502 470732 155530
rect 472360 155514 472388 159200
rect 473084 155848 473136 155854
rect 473084 155790 473136 155796
rect 470520 155366 470640 155394
rect 470416 154624 470468 154630
rect 470416 154566 470468 154572
rect 469324 151786 469812 151814
rect 469784 150226 469812 151786
rect 470428 150226 470456 154566
rect 470612 151814 470640 155366
rect 470704 155106 470732 155502
rect 472348 155508 472400 155514
rect 472348 155450 472400 155456
rect 472348 155304 472400 155310
rect 472348 155246 472400 155252
rect 470692 155100 470744 155106
rect 470692 155042 470744 155048
rect 471980 154828 472032 154834
rect 471980 154770 472032 154776
rect 471704 154760 471756 154766
rect 471704 154702 471756 154708
rect 470612 151786 471100 151814
rect 471072 150226 471100 151786
rect 471716 150226 471744 154702
rect 463378 150146 463430 150152
rect 463390 149940 463418 150146
rect 464034 149940 464062 150198
rect 464678 149940 464706 150198
rect 465322 149940 465350 150198
rect 465966 149940 465994 150198
rect 466610 149940 466638 150198
rect 467254 149940 467282 150198
rect 467898 149940 467926 150198
rect 468024 150204 468076 150210
rect 468496 150198 468570 150226
rect 468024 150146 468076 150152
rect 468542 149940 468570 150198
rect 469174 150204 469226 150210
rect 469784 150198 469858 150226
rect 470428 150198 470502 150226
rect 471072 150198 471146 150226
rect 471716 150198 471790 150226
rect 471992 150210 472020 154770
rect 472360 150226 472388 155246
rect 473096 153202 473124 155790
rect 473188 155310 473216 159200
rect 473636 155712 473688 155718
rect 473636 155654 473688 155660
rect 473360 155644 473412 155650
rect 473360 155586 473412 155592
rect 473176 155304 473228 155310
rect 473176 155246 473228 155252
rect 473084 153196 473136 153202
rect 473084 153138 473136 153144
rect 473372 151814 473400 155586
rect 473648 153134 473676 155654
rect 473912 155576 473964 155582
rect 473912 155518 473964 155524
rect 473636 153128 473688 153134
rect 473636 153070 473688 153076
rect 473924 151814 473952 155518
rect 474016 155038 474044 159200
rect 474740 155780 474792 155786
rect 474740 155722 474792 155728
rect 474004 155032 474056 155038
rect 474004 154974 474056 154980
rect 474752 153066 474780 155722
rect 474844 155650 474872 159200
rect 475672 155718 475700 159200
rect 476500 155922 476528 159200
rect 476120 155916 476172 155922
rect 476120 155858 476172 155864
rect 476488 155916 476540 155922
rect 476488 155858 476540 155864
rect 475660 155712 475712 155718
rect 475660 155654 475712 155660
rect 474832 155644 474884 155650
rect 474832 155586 474884 155592
rect 474924 155372 474976 155378
rect 474924 155314 474976 155320
rect 474740 153060 474792 153066
rect 474740 153002 474792 153008
rect 473372 151786 473676 151814
rect 473924 151786 474320 151814
rect 473648 150226 473676 151786
rect 474292 150226 474320 151786
rect 474936 150226 474964 155314
rect 475568 153196 475620 153202
rect 475568 153138 475620 153144
rect 475580 150226 475608 153138
rect 476132 152794 476160 155858
rect 476212 155236 476264 155242
rect 476212 155178 476264 155184
rect 476120 152788 476172 152794
rect 476120 152730 476172 152736
rect 476224 150226 476252 155178
rect 477328 154698 477356 159200
rect 477592 155508 477644 155514
rect 477592 155450 477644 155456
rect 477500 155440 477552 155446
rect 477500 155382 477552 155388
rect 477408 155100 477460 155106
rect 477408 155042 477460 155048
rect 477316 154692 477368 154698
rect 477316 154634 477368 154640
rect 477420 153202 477448 155042
rect 477408 153196 477460 153202
rect 477408 153138 477460 153144
rect 476948 153128 477000 153134
rect 476948 153070 477000 153076
rect 476960 150226 476988 153070
rect 469174 150146 469226 150152
rect 469186 149940 469214 150146
rect 469830 149940 469858 150198
rect 470474 149940 470502 150198
rect 471118 149940 471146 150198
rect 471762 149940 471790 150198
rect 471980 150204 472032 150210
rect 472360 150198 472434 150226
rect 471980 150146 472032 150152
rect 472406 149940 472434 150198
rect 473038 150204 473090 150210
rect 473648 150198 473722 150226
rect 474292 150198 474366 150226
rect 474936 150198 475010 150226
rect 475580 150198 475654 150226
rect 476224 150198 476298 150226
rect 473038 150146 473090 150152
rect 473050 149940 473078 150146
rect 473694 149940 473722 150198
rect 474338 149940 474366 150198
rect 474982 149940 475010 150198
rect 475626 149940 475654 150198
rect 476270 149940 476298 150198
rect 476914 150198 476988 150226
rect 477512 150226 477540 155382
rect 477604 152522 477632 155450
rect 478156 155446 478184 159200
rect 479076 155786 479104 159200
rect 479064 155780 479116 155786
rect 479064 155722 479116 155728
rect 478144 155440 478196 155446
rect 478144 155382 478196 155388
rect 479904 155310 479932 159200
rect 480732 155854 480760 159200
rect 480720 155848 480772 155854
rect 480720 155790 480772 155796
rect 480720 155712 480772 155718
rect 480720 155654 480772 155660
rect 477684 155304 477736 155310
rect 477684 155246 477736 155252
rect 479892 155304 479944 155310
rect 479892 155246 479944 155252
rect 477592 152516 477644 152522
rect 477592 152458 477644 152464
rect 477696 151910 477724 155246
rect 479524 155032 479576 155038
rect 479524 154974 479576 154980
rect 478788 153196 478840 153202
rect 478788 153138 478840 153144
rect 478144 153060 478196 153066
rect 478144 153002 478196 153008
rect 477684 151904 477736 151910
rect 477684 151846 477736 151852
rect 478156 150226 478184 153002
rect 478800 150226 478828 153138
rect 479432 152788 479484 152794
rect 479432 152730 479484 152736
rect 479444 150226 479472 152730
rect 479536 151978 479564 154974
rect 480732 153066 480760 155654
rect 481560 155650 481588 159200
rect 480812 155644 480864 155650
rect 480812 155586 480864 155592
rect 481548 155644 481600 155650
rect 481548 155586 481600 155592
rect 480824 153202 480852 155586
rect 482388 155514 482416 159200
rect 482928 155916 482980 155922
rect 482928 155858 482980 155864
rect 482376 155508 482428 155514
rect 482376 155450 482428 155456
rect 481732 154692 481784 154698
rect 481732 154634 481784 154640
rect 480812 153196 480864 153202
rect 480812 153138 480864 153144
rect 481744 153134 481772 154634
rect 482008 153196 482060 153202
rect 482008 153138 482060 153144
rect 481732 153128 481784 153134
rect 481732 153070 481784 153076
rect 480720 153060 480772 153066
rect 480720 153002 480772 153008
rect 480076 152516 480128 152522
rect 480076 152458 480128 152464
rect 479524 151972 479576 151978
rect 479524 151914 479576 151920
rect 480088 150226 480116 152458
rect 481364 151972 481416 151978
rect 481364 151914 481416 151920
rect 480720 151904 480772 151910
rect 480720 151846 480772 151852
rect 480732 150226 480760 151846
rect 481376 150226 481404 151914
rect 482020 150226 482048 153138
rect 482652 153060 482704 153066
rect 482652 153002 482704 153008
rect 482664 150226 482692 153002
rect 482940 151814 482968 155858
rect 483216 155582 483244 159200
rect 483204 155576 483256 155582
rect 483204 155518 483256 155524
rect 484044 154834 484072 159200
rect 484308 155440 484360 155446
rect 484308 155382 484360 155388
rect 484032 154828 484084 154834
rect 484032 154770 484084 154776
rect 483940 153128 483992 153134
rect 483940 153070 483992 153076
rect 482940 151786 483336 151814
rect 483308 150226 483336 151786
rect 483952 150226 483980 153070
rect 484320 151814 484348 155382
rect 484872 155174 484900 159200
rect 484952 155780 485004 155786
rect 484952 155722 485004 155728
rect 484860 155168 484912 155174
rect 484860 155110 484912 155116
rect 484964 151814 484992 155722
rect 485688 155304 485740 155310
rect 485688 155246 485740 155252
rect 485700 151814 485728 155246
rect 485792 154766 485820 159200
rect 486332 155848 486384 155854
rect 486332 155790 486384 155796
rect 485872 155576 485924 155582
rect 485872 155518 485924 155524
rect 485780 154760 485832 154766
rect 485780 154702 485832 154708
rect 485884 152726 485912 155518
rect 485872 152720 485924 152726
rect 485872 152662 485924 152668
rect 486344 151814 486372 155790
rect 486620 154630 486648 159200
rect 487068 155644 487120 155650
rect 487068 155586 487120 155592
rect 486608 154624 486660 154630
rect 486608 154566 486660 154572
rect 487080 151814 487108 155586
rect 487448 155310 487476 159200
rect 488276 155922 488304 159200
rect 488264 155916 488316 155922
rect 488264 155858 488316 155864
rect 487712 155508 487764 155514
rect 487712 155450 487764 155456
rect 487436 155304 487488 155310
rect 487436 155246 487488 155252
rect 487724 151814 487752 155450
rect 489104 155174 489132 159200
rect 489932 155378 489960 159200
rect 490380 155916 490432 155922
rect 490380 155858 490432 155864
rect 489920 155372 489972 155378
rect 489920 155314 489972 155320
rect 488448 155168 488500 155174
rect 488448 155110 488500 155116
rect 489092 155168 489144 155174
rect 489092 155110 489144 155116
rect 488460 152862 488488 155110
rect 489000 154828 489052 154834
rect 489000 154770 489052 154776
rect 488908 154760 488960 154766
rect 488908 154702 488960 154708
rect 488540 154624 488592 154630
rect 488540 154566 488592 154572
rect 488448 152856 488500 152862
rect 488448 152798 488500 152804
rect 488448 152720 488500 152726
rect 488448 152662 488500 152668
rect 484320 151786 484624 151814
rect 484964 151786 485268 151814
rect 485700 151786 485912 151814
rect 486344 151786 486556 151814
rect 487080 151786 487200 151814
rect 487724 151786 487844 151814
rect 484596 150226 484624 151786
rect 485240 150226 485268 151786
rect 485884 150226 485912 151786
rect 486528 150226 486556 151786
rect 487172 150226 487200 151786
rect 487816 150226 487844 151786
rect 488460 150226 488488 152662
rect 488552 152046 488580 154566
rect 488540 152040 488592 152046
rect 488540 151982 488592 151988
rect 488920 151910 488948 154702
rect 488908 151904 488960 151910
rect 488908 151846 488960 151852
rect 489012 150226 489040 154770
rect 490392 153202 490420 155858
rect 490760 155582 490788 159200
rect 491680 155650 491708 159200
rect 492508 155718 492536 159200
rect 492496 155712 492548 155718
rect 492496 155654 492548 155660
rect 491668 155644 491720 155650
rect 491668 155586 491720 155592
rect 490748 155576 490800 155582
rect 490748 155518 490800 155524
rect 493232 155372 493284 155378
rect 493232 155314 493284 155320
rect 491208 155304 491260 155310
rect 491208 155246 491260 155252
rect 490380 153196 490432 153202
rect 490380 153138 490432 153144
rect 489644 152856 489696 152862
rect 489644 152798 489696 152804
rect 489656 150226 489684 152798
rect 490932 152040 490984 152046
rect 490932 151982 490984 151988
rect 490288 151904 490340 151910
rect 490288 151846 490340 151852
rect 490300 150226 490328 151846
rect 490944 150226 490972 151982
rect 491220 151814 491248 155246
rect 492588 155168 492640 155174
rect 492588 155110 492640 155116
rect 492220 153196 492272 153202
rect 492220 153138 492272 153144
rect 491220 151786 491616 151814
rect 491588 150226 491616 151786
rect 492232 150226 492260 153138
rect 492600 151814 492628 155110
rect 493244 151814 493272 155314
rect 493336 155242 493364 159200
rect 494164 155582 494192 159200
rect 494612 155644 494664 155650
rect 494612 155586 494664 155592
rect 493968 155576 494020 155582
rect 493968 155518 494020 155524
rect 494152 155576 494204 155582
rect 494152 155518 494204 155524
rect 493324 155236 493376 155242
rect 493324 155178 493376 155184
rect 493980 151814 494008 155518
rect 494624 151814 494652 155586
rect 494992 155310 495020 159200
rect 495348 155712 495400 155718
rect 495348 155654 495400 155660
rect 494980 155304 495032 155310
rect 494980 155246 495032 155252
rect 495360 151814 495388 155654
rect 495820 155378 495848 159200
rect 495808 155372 495860 155378
rect 495808 155314 495860 155320
rect 495808 155236 495860 155242
rect 495808 155178 495860 155184
rect 495820 151814 495848 155178
rect 496648 154766 496676 159200
rect 497476 155582 497504 159200
rect 498396 155854 498424 159200
rect 499224 155922 499252 159200
rect 499212 155916 499264 155922
rect 499212 155858 499264 155864
rect 498384 155848 498436 155854
rect 498384 155790 498436 155796
rect 499580 155848 499632 155854
rect 499580 155790 499632 155796
rect 496728 155576 496780 155582
rect 496728 155518 496780 155524
rect 497464 155576 497516 155582
rect 497464 155518 497516 155524
rect 499304 155576 499356 155582
rect 499304 155518 499356 155524
rect 496636 154760 496688 154766
rect 496636 154702 496688 154708
rect 492600 151786 492904 151814
rect 493244 151786 493548 151814
rect 493980 151786 494192 151814
rect 494624 151786 494836 151814
rect 495360 151786 495480 151814
rect 495820 151786 496124 151814
rect 492876 150226 492904 151786
rect 493520 150226 493548 151786
rect 494164 150226 494192 151786
rect 494808 150226 494836 151786
rect 495452 150226 495480 151786
rect 496096 150226 496124 151786
rect 496740 150226 496768 155518
rect 496912 155372 496964 155378
rect 496912 155314 496964 155320
rect 477512 150198 477586 150226
rect 478156 150198 478230 150226
rect 478800 150198 478874 150226
rect 479444 150198 479518 150226
rect 480088 150198 480162 150226
rect 480732 150198 480806 150226
rect 481376 150198 481450 150226
rect 482020 150198 482094 150226
rect 482664 150198 482738 150226
rect 483308 150198 483382 150226
rect 483952 150198 484026 150226
rect 484596 150198 484670 150226
rect 485240 150198 485314 150226
rect 485884 150198 485958 150226
rect 486528 150198 486602 150226
rect 487172 150198 487246 150226
rect 487816 150198 487890 150226
rect 488460 150198 488534 150226
rect 489012 150198 489086 150226
rect 489656 150198 489730 150226
rect 490300 150198 490374 150226
rect 490944 150198 491018 150226
rect 491588 150198 491662 150226
rect 492232 150198 492306 150226
rect 492876 150198 492950 150226
rect 493520 150198 493594 150226
rect 494164 150198 494238 150226
rect 494808 150198 494882 150226
rect 495452 150198 495526 150226
rect 496096 150198 496170 150226
rect 496740 150198 496814 150226
rect 496924 150210 496952 155314
rect 497372 155304 497424 155310
rect 497372 155246 497424 155252
rect 497384 150226 497412 155246
rect 498200 154760 498252 154766
rect 498200 154702 498252 154708
rect 498212 151814 498240 154702
rect 498212 151786 498700 151814
rect 498672 150226 498700 151786
rect 499316 150226 499344 155518
rect 499592 151814 499620 155790
rect 500052 155514 500080 159200
rect 500592 155916 500644 155922
rect 500592 155858 500644 155864
rect 500040 155508 500092 155514
rect 500040 155450 500092 155456
rect 499592 151786 499988 151814
rect 499960 150226 499988 151786
rect 500604 150226 500632 155858
rect 500880 155530 500908 159200
rect 501708 155582 501736 159200
rect 501696 155576 501748 155582
rect 500880 155502 501000 155530
rect 501696 155518 501748 155524
rect 502432 155576 502484 155582
rect 502432 155518 502484 155524
rect 476914 149940 476942 150198
rect 477558 149940 477586 150198
rect 478202 149940 478230 150198
rect 478846 149940 478874 150198
rect 479490 149940 479518 150198
rect 480134 149940 480162 150198
rect 480778 149940 480806 150198
rect 481422 149940 481450 150198
rect 482066 149940 482094 150198
rect 482710 149940 482738 150198
rect 483354 149940 483382 150198
rect 483998 149940 484026 150198
rect 484642 149940 484670 150198
rect 485286 149940 485314 150198
rect 485930 149940 485958 150198
rect 486574 149940 486602 150198
rect 487218 149940 487246 150198
rect 487862 149940 487890 150198
rect 488506 149940 488534 150198
rect 489058 149940 489086 150198
rect 489702 149940 489730 150198
rect 490346 149940 490374 150198
rect 490990 149940 491018 150198
rect 491634 149940 491662 150198
rect 492278 149940 492306 150198
rect 492922 149940 492950 150198
rect 493566 149940 493594 150198
rect 494210 149940 494238 150198
rect 494854 149940 494882 150198
rect 495498 149940 495526 150198
rect 496142 149940 496170 150198
rect 496786 149940 496814 150198
rect 496912 150204 496964 150210
rect 497384 150198 497458 150226
rect 496912 150146 496964 150152
rect 497430 149940 497458 150198
rect 498062 150204 498114 150210
rect 498672 150198 498746 150226
rect 499316 150198 499390 150226
rect 499960 150198 500034 150226
rect 500604 150198 500678 150226
rect 500972 150210 501000 155502
rect 501236 155508 501288 155514
rect 501236 155450 501288 155456
rect 501248 150226 501276 155450
rect 502444 151814 502472 155518
rect 502536 152930 502564 159200
rect 503364 155242 503392 159200
rect 504192 159174 504312 159200
rect 503352 155236 503404 155242
rect 503352 155178 503404 155184
rect 503812 155236 503864 155242
rect 503812 155178 503864 155184
rect 502524 152924 502576 152930
rect 502524 152866 502576 152872
rect 503168 152924 503220 152930
rect 503168 152866 503220 152872
rect 502444 151786 502564 151814
rect 502536 150226 502564 151786
rect 503180 150226 503208 152866
rect 503824 150226 503852 155178
rect 504468 150226 504496 159310
rect 505098 159200 505154 160400
rect 505926 159200 505982 160400
rect 506492 159310 506704 159338
rect 505112 150226 505140 159200
rect 505940 151814 505968 159200
rect 506492 155530 506520 159310
rect 506676 159202 506704 159310
rect 506754 159202 506810 160400
rect 506676 159200 506810 159202
rect 507582 159200 507638 160400
rect 508410 159200 508466 160400
rect 509238 159200 509294 160400
rect 510066 159200 510122 160400
rect 510894 159200 510950 160400
rect 511814 159200 511870 160400
rect 512642 159200 512698 160400
rect 513470 159200 513526 160400
rect 514298 159200 514354 160400
rect 515126 159200 515182 160400
rect 515954 159200 516010 160400
rect 516782 159200 516838 160400
rect 517610 159200 517666 160400
rect 518530 159200 518586 160400
rect 519358 159200 519414 160400
rect 520186 159200 520242 160400
rect 520922 159216 520978 159225
rect 506676 159174 506796 159200
rect 505848 151786 505968 151814
rect 506400 155502 506520 155530
rect 505848 150226 505876 151786
rect 498062 150146 498114 150152
rect 498074 149940 498102 150146
rect 498718 149940 498746 150198
rect 499362 149940 499390 150198
rect 500006 149940 500034 150198
rect 500650 149940 500678 150198
rect 500960 150204 501012 150210
rect 501248 150198 501322 150226
rect 500960 150146 501012 150152
rect 501294 149940 501322 150198
rect 501926 150204 501978 150210
rect 502536 150198 502610 150226
rect 503180 150198 503254 150226
rect 503824 150198 503898 150226
rect 504468 150198 504542 150226
rect 505112 150198 505186 150226
rect 501926 150146 501978 150152
rect 501938 149940 501966 150146
rect 502582 149940 502610 150198
rect 503226 149940 503254 150198
rect 503870 149940 503898 150198
rect 504514 149940 504542 150198
rect 505158 149940 505186 150198
rect 505802 150198 505876 150226
rect 506400 150226 506428 155502
rect 507596 151978 507624 159200
rect 508424 155582 508452 159200
rect 509056 155916 509108 155922
rect 509056 155858 509108 155864
rect 507768 155576 507820 155582
rect 507768 155518 507820 155524
rect 508412 155576 508464 155582
rect 508412 155518 508464 155524
rect 507032 151972 507084 151978
rect 507032 151914 507084 151920
rect 507584 151972 507636 151978
rect 507584 151914 507636 151920
rect 507044 150226 507072 151914
rect 507780 150226 507808 155518
rect 508412 152244 508464 152250
rect 508412 152186 508464 152192
rect 508424 150226 508452 152186
rect 509068 150226 509096 155858
rect 509252 154574 509280 159200
rect 510080 155922 510108 159200
rect 510068 155916 510120 155922
rect 510068 155858 510120 155864
rect 510528 155576 510580 155582
rect 510528 155518 510580 155524
rect 509700 154828 509752 154834
rect 509700 154770 509752 154776
rect 509160 154546 509280 154574
rect 509160 152250 509188 154546
rect 509148 152244 509200 152250
rect 509148 152186 509200 152192
rect 509712 150226 509740 154770
rect 510540 151814 510568 155518
rect 510908 154834 510936 159200
rect 511828 155582 511856 159200
rect 511816 155576 511868 155582
rect 511816 155518 511868 155524
rect 512276 155576 512328 155582
rect 512276 155518 512328 155524
rect 510988 155236 511040 155242
rect 510988 155178 511040 155184
rect 510896 154828 510948 154834
rect 510896 154770 510948 154776
rect 510356 151786 510568 151814
rect 510356 150226 510384 151786
rect 511000 150226 511028 155178
rect 511632 155032 511684 155038
rect 511632 154974 511684 154980
rect 511644 150226 511672 154974
rect 512288 150226 512316 155518
rect 512656 155242 512684 159200
rect 512920 155304 512972 155310
rect 512920 155246 512972 155252
rect 512644 155236 512696 155242
rect 512644 155178 512696 155184
rect 512932 150226 512960 155246
rect 513484 155038 513512 159200
rect 513564 155644 513616 155650
rect 513564 155586 513616 155592
rect 513472 155032 513524 155038
rect 513472 154974 513524 154980
rect 513576 150226 513604 155586
rect 514312 155582 514340 159200
rect 514300 155576 514352 155582
rect 514300 155518 514352 155524
rect 514852 155576 514904 155582
rect 514852 155518 514904 155524
rect 514208 155508 514260 155514
rect 514208 155450 514260 155456
rect 514220 150226 514248 155450
rect 514864 150226 514892 155518
rect 515140 155310 515168 159200
rect 515496 155712 515548 155718
rect 515496 155654 515548 155660
rect 515128 155304 515180 155310
rect 515128 155246 515180 155252
rect 515508 150226 515536 155654
rect 515968 155650 515996 159200
rect 516048 155916 516100 155922
rect 516048 155858 516100 155864
rect 515956 155644 516008 155650
rect 515956 155586 516008 155592
rect 506400 150198 506474 150226
rect 507044 150198 507118 150226
rect 505802 149940 505830 150198
rect 506446 149940 506474 150198
rect 507090 149940 507118 150198
rect 507734 150198 507808 150226
rect 508378 150198 508452 150226
rect 509022 150198 509096 150226
rect 509666 150198 509740 150226
rect 510310 150198 510384 150226
rect 510954 150198 511028 150226
rect 511598 150198 511672 150226
rect 512242 150198 512316 150226
rect 512886 150198 512960 150226
rect 513530 150198 513604 150226
rect 514174 150198 514248 150226
rect 514818 150198 514892 150226
rect 515462 150198 515536 150226
rect 516060 150226 516088 155858
rect 516796 155514 516824 159200
rect 517336 155780 517388 155786
rect 517336 155722 517388 155728
rect 516784 155508 516836 155514
rect 516784 155450 516836 155456
rect 516784 155236 516836 155242
rect 516784 155178 516836 155184
rect 516796 150226 516824 155178
rect 516060 150198 516134 150226
rect 507734 149940 507762 150198
rect 508378 149940 508406 150198
rect 509022 149940 509050 150198
rect 509666 149940 509694 150198
rect 510310 149940 510338 150198
rect 510954 149940 510982 150198
rect 511598 149940 511626 150198
rect 512242 149940 512270 150198
rect 512886 149940 512914 150198
rect 513530 149940 513558 150198
rect 514174 149940 514202 150198
rect 514818 149940 514846 150198
rect 515462 149940 515490 150198
rect 516106 149940 516134 150198
rect 516750 150198 516824 150226
rect 517348 150226 517376 155722
rect 517624 155582 517652 159200
rect 518544 155718 518572 159200
rect 519372 155922 519400 159200
rect 519542 157720 519598 157729
rect 519542 157655 519598 157664
rect 519360 155916 519412 155922
rect 519360 155858 519412 155864
rect 518532 155712 518584 155718
rect 518532 155654 518584 155660
rect 517612 155576 517664 155582
rect 517612 155518 517664 155524
rect 518072 155372 518124 155378
rect 518072 155314 518124 155320
rect 518084 150226 518112 155314
rect 518808 155304 518860 155310
rect 518808 155246 518860 155252
rect 517348 150198 517422 150226
rect 516750 149940 516778 150198
rect 517394 149940 517422 150198
rect 518038 150198 518112 150226
rect 518038 149940 518066 150198
rect 518820 149954 518848 155246
rect 518696 149926 518848 149954
rect 519556 147937 519584 157655
rect 519634 156224 519690 156233
rect 519634 156159 519690 156168
rect 519542 147928 519598 147937
rect 519542 147863 519598 147872
rect 519648 146577 519676 156159
rect 520200 155242 520228 159200
rect 521014 159200 521070 160400
rect 521842 159200 521898 160400
rect 522670 159200 522726 160400
rect 523498 159200 523554 160400
rect 520922 159151 520978 159160
rect 520188 155236 520240 155242
rect 520188 155178 520240 155184
rect 519726 154728 519782 154737
rect 519726 154663 519782 154672
rect 519634 146568 519690 146577
rect 519634 146503 519690 146512
rect 519740 145217 519768 154663
rect 519818 153232 519874 153241
rect 519818 153167 519874 153176
rect 519726 145208 519782 145217
rect 519726 145143 519782 145152
rect 519832 143857 519860 153167
rect 519910 150240 519966 150249
rect 519910 150175 519966 150184
rect 519818 143848 519874 143857
rect 519818 143783 519874 143792
rect 519924 141137 519952 150175
rect 520936 149297 520964 159151
rect 521028 155786 521056 159200
rect 521016 155780 521068 155786
rect 521016 155722 521068 155728
rect 521856 155378 521884 159200
rect 521844 155372 521896 155378
rect 521844 155314 521896 155320
rect 522684 155310 522712 159200
rect 522672 155304 522724 155310
rect 522672 155246 522724 155252
rect 523512 155242 523540 159200
rect 521844 155236 521896 155242
rect 521844 155178 521896 155184
rect 523500 155236 523552 155242
rect 523500 155178 523552 155184
rect 521014 151736 521070 151745
rect 521014 151671 521070 151680
rect 520922 149288 520978 149297
rect 520922 149223 520978 149232
rect 520922 145888 520978 145897
rect 520922 145823 520978 145832
rect 520278 144392 520334 144401
rect 520278 144327 520334 144336
rect 519910 141128 519966 141137
rect 519910 141063 519966 141072
rect 520292 135697 520320 144327
rect 520738 142896 520794 142905
rect 520738 142831 520794 142840
rect 520278 135688 520334 135697
rect 520278 135623 520334 135632
rect 117226 135552 117282 135561
rect 117226 135487 117282 135496
rect 520752 134337 520780 142831
rect 520936 137057 520964 145823
rect 521028 142497 521056 151671
rect 521106 148744 521162 148753
rect 521106 148679 521162 148688
rect 521014 142488 521070 142497
rect 521014 142423 521070 142432
rect 521014 141400 521070 141409
rect 521014 141335 521070 141344
rect 520922 137048 520978 137057
rect 520922 136983 520978 136992
rect 520738 134328 520794 134337
rect 520738 134263 520794 134272
rect 520278 134056 520334 134065
rect 520278 133991 520334 134000
rect 117134 133648 117190 133657
rect 117134 133583 117190 133592
rect 520186 131064 520242 131073
rect 520186 130999 520242 131008
rect 519910 129568 519966 129577
rect 519910 129503 519966 129512
rect 519542 128072 519598 128081
rect 519542 128007 519598 128016
rect 519266 123584 519322 123593
rect 519266 123519 519322 123528
rect 117042 118280 117098 118289
rect 117042 118215 117098 118224
rect 519280 116657 519308 123519
rect 519556 120737 519584 128007
rect 519726 126576 519782 126585
rect 519726 126511 519782 126520
rect 519542 120728 519598 120737
rect 519542 120663 519598 120672
rect 519740 119377 519768 126511
rect 519818 125080 519874 125089
rect 519818 125015 519874 125024
rect 519726 119368 519782 119377
rect 519726 119303 519782 119312
rect 519832 118017 519860 125015
rect 519924 122097 519952 129503
rect 520200 123457 520228 130999
rect 520292 126177 520320 133991
rect 521028 132977 521056 141335
rect 521120 139777 521148 148679
rect 521198 147384 521254 147393
rect 521198 147319 521254 147328
rect 521106 139768 521162 139777
rect 521106 139703 521162 139712
rect 521212 138417 521240 147319
rect 521290 139904 521346 139913
rect 521290 139839 521346 139848
rect 521198 138408 521254 138417
rect 521198 138343 521254 138352
rect 521198 136912 521254 136921
rect 521198 136847 521254 136856
rect 521106 135416 521162 135425
rect 521106 135351 521162 135360
rect 521014 132968 521070 132977
rect 521014 132903 521070 132912
rect 521014 132560 521070 132569
rect 521014 132495 521070 132504
rect 520278 126168 520334 126177
rect 520278 126103 520334 126112
rect 521028 124817 521056 132495
rect 521120 127537 521148 135351
rect 521212 128897 521240 136847
rect 521304 131617 521332 139839
rect 521382 138408 521438 138417
rect 521382 138343 521438 138352
rect 521290 131608 521346 131617
rect 521290 131543 521346 131552
rect 521396 130257 521424 138343
rect 521382 130248 521438 130257
rect 521382 130183 521438 130192
rect 521198 128888 521254 128897
rect 521198 128823 521254 128832
rect 521106 127528 521162 127537
rect 521106 127463 521162 127472
rect 521014 124808 521070 124817
rect 521014 124743 521070 124752
rect 520186 123448 520242 123457
rect 520186 123383 520242 123392
rect 519910 122088 519966 122097
rect 519910 122023 519966 122032
rect 520094 122088 520150 122097
rect 520094 122023 520150 122032
rect 519910 119232 519966 119241
rect 519910 119167 519966 119176
rect 519818 118008 519874 118017
rect 519818 117943 519874 117952
rect 519726 117736 519782 117745
rect 519726 117671 519782 117680
rect 519266 116648 519322 116657
rect 519266 116583 519322 116592
rect 116950 116376 117006 116385
rect 116950 116311 117006 116320
rect 519266 113248 519322 113257
rect 519266 113183 519322 113192
rect 116858 112568 116914 112577
rect 116858 112503 116914 112512
rect 519280 107137 519308 113183
rect 519740 111217 519768 117671
rect 519818 114744 519874 114753
rect 519818 114679 519874 114688
rect 519726 111208 519782 111217
rect 519726 111143 519782 111152
rect 519634 108760 519690 108769
rect 519634 108695 519690 108704
rect 519266 107128 519322 107137
rect 519266 107063 519322 107072
rect 519082 104408 519138 104417
rect 519082 104343 519138 104352
rect 116766 102912 116822 102921
rect 116766 102847 116822 102856
rect 519096 98977 519124 104343
rect 519648 103057 519676 108695
rect 519832 108497 519860 114679
rect 519924 112577 519952 119167
rect 520002 116240 520058 116249
rect 520002 116175 520058 116184
rect 519910 112568 519966 112577
rect 519910 112503 519966 112512
rect 520016 109857 520044 116175
rect 520108 115297 520136 122023
rect 520186 120728 520242 120737
rect 520186 120663 520242 120672
rect 520094 115288 520150 115297
rect 520094 115223 520150 115232
rect 520200 113937 520228 120663
rect 520186 113928 520242 113937
rect 520186 113863 520242 113872
rect 520094 111752 520150 111761
rect 520094 111687 520150 111696
rect 520002 109848 520058 109857
rect 520002 109783 520058 109792
rect 519818 108488 519874 108497
rect 519818 108423 519874 108432
rect 519726 107400 519782 107409
rect 519726 107335 519782 107344
rect 519634 103048 519690 103057
rect 519634 102983 519690 102992
rect 519740 101697 519768 107335
rect 519910 105904 519966 105913
rect 519910 105839 519966 105848
rect 519726 101688 519782 101697
rect 519726 101623 519782 101632
rect 519924 100337 519952 105839
rect 520108 105777 520136 111687
rect 520186 110256 520242 110265
rect 520186 110191 520242 110200
rect 520094 105768 520150 105777
rect 520094 105703 520150 105712
rect 520200 104553 520228 110191
rect 520186 104544 520242 104553
rect 520186 104479 520242 104488
rect 520094 102912 520150 102921
rect 520094 102847 520150 102856
rect 519910 100328 519966 100337
rect 519910 100263 519966 100272
rect 519450 99920 519506 99929
rect 519450 99855 519506 99864
rect 519082 98968 519138 98977
rect 519082 98903 519138 98912
rect 519464 94897 519492 99855
rect 519818 98424 519874 98433
rect 519818 98359 519874 98368
rect 519542 96928 519598 96937
rect 519542 96863 519598 96872
rect 519450 94888 519506 94897
rect 519450 94823 519506 94832
rect 519082 94072 519138 94081
rect 519082 94007 519138 94016
rect 116582 91352 116638 91361
rect 116582 91287 116638 91296
rect 519096 89457 519124 94007
rect 519266 92576 519322 92585
rect 519266 92511 519322 92520
rect 519082 89448 519138 89457
rect 519082 89383 519138 89392
rect 115940 88324 115992 88330
rect 115940 88266 115992 88272
rect 115952 87553 115980 88266
rect 519280 88097 519308 92511
rect 519556 92177 519584 96863
rect 519726 95432 519782 95441
rect 519726 95367 519782 95376
rect 519542 92168 519598 92177
rect 519542 92103 519598 92112
rect 519450 91080 519506 91089
rect 519450 91015 519506 91024
rect 519266 88088 519322 88097
rect 519266 88023 519322 88032
rect 115938 87544 115994 87553
rect 115938 87479 115994 87488
rect 114282 87272 114338 87281
rect 114282 87207 114338 87216
rect 114192 80028 114244 80034
rect 114192 79970 114244 79976
rect 114296 78674 114324 87207
rect 116400 86964 116452 86970
rect 116400 86906 116452 86912
rect 116412 85649 116440 86906
rect 116398 85640 116454 85649
rect 116398 85575 116454 85584
rect 519464 85377 519492 91015
rect 519740 90817 519768 95367
rect 519832 93537 519860 98359
rect 520108 97617 520136 102847
rect 520186 101416 520242 101425
rect 520186 101351 520242 101360
rect 520094 97608 520150 97617
rect 520094 97543 520150 97552
rect 520200 96257 520228 101351
rect 520186 96248 520242 96257
rect 520186 96183 520242 96192
rect 521856 93854 521884 155178
rect 521672 93826 521884 93854
rect 519818 93528 519874 93537
rect 519818 93463 519874 93472
rect 519726 90808 519782 90817
rect 519726 90743 519782 90752
rect 519910 89584 519966 89593
rect 519910 89519 519966 89528
rect 519726 86592 519782 86601
rect 519726 86527 519782 86536
rect 519450 85368 519506 85377
rect 519450 85303 519506 85312
rect 519082 85096 519138 85105
rect 519082 85031 519138 85040
rect 116584 83972 116636 83978
rect 116584 83914 116636 83920
rect 116596 83745 116624 83914
rect 116582 83736 116638 83745
rect 116582 83671 116638 83680
rect 116308 82816 116360 82822
rect 116308 82758 116360 82764
rect 116320 81841 116348 82758
rect 116306 81832 116362 81841
rect 116306 81767 116362 81776
rect 115940 80028 115992 80034
rect 115940 79970 115992 79976
rect 115952 79937 115980 79970
rect 519096 79937 519124 85031
rect 519740 81297 519768 86527
rect 519924 84017 519952 89519
rect 520002 88088 520058 88097
rect 520002 88023 520058 88032
rect 519910 84008 519966 84017
rect 519910 83943 519966 83952
rect 520016 82657 520044 88023
rect 521566 86728 521622 86737
rect 521672 86714 521700 93826
rect 521622 86686 521700 86714
rect 521566 86663 521622 86672
rect 520094 83600 520150 83609
rect 520094 83535 520150 83544
rect 520002 82648 520058 82657
rect 520002 82583 520058 82592
rect 519726 81288 519782 81297
rect 519726 81223 519782 81232
rect 115938 79928 115994 79937
rect 115938 79863 115994 79872
rect 519082 79928 519138 79937
rect 519082 79863 519138 79872
rect 114284 78668 114336 78674
rect 114284 78610 114336 78616
rect 116216 78668 116268 78674
rect 116216 78610 116268 78616
rect 116228 78033 116256 78610
rect 520108 78577 520136 83535
rect 520186 82104 520242 82113
rect 520186 82039 520242 82048
rect 520094 78568 520150 78577
rect 520094 78503 520150 78512
rect 116214 78024 116270 78033
rect 116214 77959 116270 77968
rect 520200 77217 520228 82039
rect 521106 80744 521162 80753
rect 521106 80679 521162 80688
rect 520554 79248 520610 79257
rect 520554 79183 520610 79192
rect 520186 77208 520242 77217
rect 520186 77143 520242 77152
rect 520568 74633 520596 79183
rect 521014 77752 521070 77761
rect 521014 77687 521070 77696
rect 520554 74624 520610 74633
rect 520554 74559 520610 74568
rect 116674 74080 116730 74089
rect 116674 74015 116730 74024
rect 116582 72176 116638 72185
rect 116582 72111 116638 72120
rect 116596 71806 116624 72111
rect 114192 71800 114244 71806
rect 114192 71742 114244 71748
rect 116584 71800 116636 71806
rect 116584 71742 116636 71748
rect 114100 69080 114152 69086
rect 114100 69022 114152 69028
rect 114008 67652 114060 67658
rect 114008 67594 114060 67600
rect 113916 66292 113968 66298
rect 113916 66234 113968 66240
rect 113364 64728 113416 64734
rect 113364 64670 113416 64676
rect 113376 64569 113404 64670
rect 113362 64560 113418 64569
rect 113362 64495 113418 64504
rect 113824 63572 113876 63578
rect 113824 63514 113876 63520
rect 112444 62144 112496 62150
rect 112444 62086 112496 62092
rect 110326 59392 110382 59401
rect 110326 59327 110382 59336
rect 110340 55214 110368 59327
rect 109696 55186 110368 55214
rect 109406 3632 109462 3641
rect 109406 3567 109462 3576
rect 109420 3233 109448 3567
rect 109498 3496 109554 3505
rect 109498 3431 109554 3440
rect 109406 3224 109462 3233
rect 109406 3159 109462 3168
rect 33046 2680 33102 2689
rect 76194 2680 76250 2689
rect 76038 2638 76194 2666
rect 33046 2615 33102 2624
rect 76194 2615 76250 2624
rect 88890 2680 88946 2689
rect 88890 2615 88946 2624
rect 98274 2680 98330 2689
rect 98274 2615 98330 2624
rect 100298 2680 100354 2689
rect 100298 2615 100354 2624
rect 102138 2680 102194 2689
rect 102138 2615 102194 2624
rect 102322 2680 102378 2689
rect 102322 2615 102378 2624
rect 26054 2136 26110 2145
rect 2700 1358 2728 2108
rect 2688 1352 2740 1358
rect 2688 1294 2740 1300
rect 6012 1290 6040 2108
rect 6000 1284 6052 1290
rect 6000 1226 6052 1232
rect 9324 1222 9352 2108
rect 12636 1601 12664 2108
rect 15948 1737 15976 2108
rect 19352 1873 19380 2108
rect 22678 2094 22968 2122
rect 25990 2094 26054 2122
rect 22940 2009 22968 2094
rect 26054 2071 26110 2080
rect 22926 2000 22982 2009
rect 22926 1935 22982 1944
rect 19338 1864 19394 1873
rect 19338 1799 19394 1808
rect 15934 1728 15990 1737
rect 15934 1663 15990 1672
rect 12622 1592 12678 1601
rect 12622 1527 12678 1536
rect 29288 1426 29316 2108
rect 32692 1494 32720 2108
rect 32680 1488 32732 1494
rect 32680 1430 32732 1436
rect 29276 1420 29328 1426
rect 29276 1362 29328 1368
rect 9312 1216 9364 1222
rect 9312 1158 9364 1164
rect 32784 870 32904 898
rect 32784 800 32812 870
rect 32770 -400 32826 800
rect 32876 762 32904 870
rect 33060 762 33088 2615
rect 36004 1154 36032 2108
rect 35992 1148 36044 1154
rect 35992 1090 36044 1096
rect 39316 1086 39344 2108
rect 39304 1080 39356 1086
rect 39304 1022 39356 1028
rect 42628 1018 42656 2108
rect 42616 1012 42668 1018
rect 42616 954 42668 960
rect 46032 950 46060 2108
rect 46020 944 46072 950
rect 46020 886 46072 892
rect 49344 882 49372 2108
rect 49332 876 49384 882
rect 49332 818 49384 824
rect 52656 814 52684 2108
rect 55968 1465 55996 2108
rect 55954 1456 56010 1465
rect 55954 1391 56010 1400
rect 32876 734 33088 762
rect 52644 808 52696 814
rect 52644 750 52696 756
rect 59372 746 59400 2108
rect 59360 740 59412 746
rect 59360 682 59412 688
rect 62684 678 62712 2108
rect 65996 1766 66024 2108
rect 65984 1760 66036 1766
rect 65984 1702 66036 1708
rect 62672 672 62724 678
rect 62672 614 62724 620
rect 69308 610 69336 2108
rect 72712 1562 72740 2108
rect 72700 1556 72752 1562
rect 72700 1498 72752 1504
rect 69296 604 69348 610
rect 69296 546 69348 552
rect 79336 542 79364 2108
rect 82648 1630 82676 2108
rect 86052 1698 86080 2108
rect 88904 1766 88932 2615
rect 94410 2408 94466 2417
rect 94410 2343 94466 2352
rect 89364 1834 89392 2108
rect 92676 1902 92704 2108
rect 94424 1902 94452 2343
rect 98288 2281 98316 2615
rect 98274 2272 98330 2281
rect 98274 2207 98330 2216
rect 95988 1902 96016 2108
rect 92664 1896 92716 1902
rect 92664 1838 92716 1844
rect 94412 1896 94464 1902
rect 94412 1838 94464 1844
rect 95976 1896 96028 1902
rect 95976 1838 96028 1844
rect 89352 1828 89404 1834
rect 89352 1770 89404 1776
rect 99392 1766 99420 2108
rect 88892 1760 88944 1766
rect 88892 1702 88944 1708
rect 99380 1760 99432 1766
rect 99380 1702 99432 1708
rect 86040 1692 86092 1698
rect 86040 1634 86092 1640
rect 82636 1624 82688 1630
rect 82636 1566 82688 1572
rect 100312 1562 100340 2615
rect 102152 2417 102180 2615
rect 102138 2408 102194 2417
rect 102138 2343 102194 2352
rect 100300 1556 100352 1562
rect 100300 1498 100352 1504
rect 102336 1329 102364 2615
rect 109512 2281 109540 3431
rect 109498 2272 109554 2281
rect 109498 2207 109554 2216
rect 102704 1970 102732 2108
rect 102692 1964 102744 1970
rect 102692 1906 102744 1912
rect 106016 1902 106044 2108
rect 106004 1896 106056 1902
rect 106004 1838 106056 1844
rect 109328 1834 109356 2108
rect 109696 1902 109724 55186
rect 110326 53952 110382 53961
rect 109788 53910 110326 53938
rect 109684 1896 109736 1902
rect 109684 1838 109736 1844
rect 105820 1828 105872 1834
rect 105820 1770 105872 1776
rect 109040 1828 109092 1834
rect 109040 1770 109092 1776
rect 109316 1828 109368 1834
rect 109316 1770 109368 1776
rect 105832 1698 105860 1770
rect 109052 1698 109080 1770
rect 109788 1698 109816 53910
rect 110326 53887 110382 53896
rect 110326 51096 110382 51105
rect 109880 51054 110326 51082
rect 105820 1692 105872 1698
rect 105820 1634 105872 1640
rect 105912 1692 105964 1698
rect 105912 1634 105964 1640
rect 108948 1692 109000 1698
rect 108948 1634 109000 1640
rect 109040 1692 109092 1698
rect 109040 1634 109092 1640
rect 109776 1692 109828 1698
rect 109776 1634 109828 1640
rect 105636 1624 105688 1630
rect 105924 1578 105952 1634
rect 105688 1572 105952 1578
rect 105636 1566 105952 1572
rect 105648 1550 105952 1566
rect 108960 1578 108988 1634
rect 109880 1630 109908 51054
rect 110326 51031 110382 51040
rect 110326 48376 110382 48385
rect 109972 48334 110326 48362
rect 109868 1624 109920 1630
rect 108960 1550 109172 1578
rect 109868 1566 109920 1572
rect 109972 1562 110000 48334
rect 110326 48311 110382 48320
rect 110326 47152 110382 47161
rect 110326 47087 110382 47096
rect 110340 45554 110368 47087
rect 110064 45526 110368 45554
rect 109144 1442 109172 1550
rect 109960 1556 110012 1562
rect 109960 1498 110012 1504
rect 110064 1442 110092 45526
rect 110326 42936 110382 42945
rect 110326 42871 110382 42880
rect 110340 26234 110368 42871
rect 110156 26206 110368 26234
rect 110156 4049 110184 26206
rect 111156 5568 111208 5574
rect 111156 5510 111208 5516
rect 110142 4040 110198 4049
rect 110142 3975 110198 3984
rect 110142 2952 110198 2961
rect 110142 2887 110198 2896
rect 110156 1562 110184 2887
rect 111064 2848 111116 2854
rect 111062 2816 111064 2825
rect 111116 2816 111118 2825
rect 111062 2751 111118 2760
rect 110144 1556 110196 1562
rect 110144 1498 110196 1504
rect 109144 1414 110092 1442
rect 98274 1320 98330 1329
rect 98274 1255 98330 1264
rect 102322 1320 102378 1329
rect 102322 1255 102378 1264
rect 98288 800 98316 1255
rect 111168 1222 111196 5510
rect 111800 4208 111852 4214
rect 111800 4150 111852 4156
rect 111812 1290 111840 4150
rect 112456 1834 112484 62086
rect 112536 44192 112588 44198
rect 112536 44134 112588 44140
rect 112444 1828 112496 1834
rect 112444 1770 112496 1776
rect 111800 1284 111852 1290
rect 111800 1226 111852 1232
rect 111156 1216 111208 1222
rect 111156 1158 111208 1164
rect 79324 536 79376 542
rect 79324 478 79376 484
rect 98274 -400 98330 800
rect 108224 746 108436 762
rect 108212 740 108448 746
rect 108264 734 108396 740
rect 108212 682 108264 688
rect 108396 682 108448 688
rect 112548 406 112576 44134
rect 112628 34536 112680 34542
rect 112628 34478 112680 34484
rect 112640 610 112668 34478
rect 112720 29028 112772 29034
rect 112720 28970 112772 28976
rect 112732 882 112760 28970
rect 112812 24880 112864 24886
rect 112812 24822 112864 24828
rect 112824 1018 112852 24822
rect 112904 22160 112956 22166
rect 112904 22102 112956 22108
rect 112916 1154 112944 22102
rect 113836 7721 113864 63514
rect 113928 19009 113956 66234
rect 114020 30433 114048 67594
rect 114112 41857 114140 69022
rect 114204 53145 114232 71742
rect 116306 70272 116362 70281
rect 116306 70207 116362 70216
rect 116320 69086 116348 70207
rect 116308 69080 116360 69086
rect 116308 69022 116360 69028
rect 116122 68368 116178 68377
rect 116122 68303 116178 68312
rect 116136 67658 116164 68303
rect 116124 67652 116176 67658
rect 116124 67594 116176 67600
rect 116582 66464 116638 66473
rect 116582 66399 116638 66408
rect 116596 66298 116624 66399
rect 116584 66292 116636 66298
rect 116584 66234 116636 66240
rect 116688 64874 116716 74015
rect 521028 73817 521056 77687
rect 521120 75993 521148 80679
rect 521198 76256 521254 76265
rect 521198 76191 521254 76200
rect 521106 75984 521162 75993
rect 521106 75919 521162 75928
rect 521106 74760 521162 74769
rect 521106 74695 521162 74704
rect 521014 73808 521070 73817
rect 521014 73743 521070 73752
rect 521014 73264 521070 73273
rect 521014 73199 521070 73208
rect 520002 71768 520058 71777
rect 520002 71703 520058 71712
rect 519266 70272 519322 70281
rect 519266 70207 519322 70216
rect 519280 66473 519308 70207
rect 520016 67833 520044 71703
rect 521028 69193 521056 73199
rect 521120 70553 521148 74695
rect 521212 71913 521240 76191
rect 521198 71904 521254 71913
rect 521198 71839 521254 71848
rect 521106 70544 521162 70553
rect 521106 70479 521162 70488
rect 521014 69184 521070 69193
rect 521014 69119 521070 69128
rect 520186 68776 520242 68785
rect 520186 68711 520242 68720
rect 520002 67824 520058 67833
rect 520002 67759 520058 67768
rect 519910 67416 519966 67425
rect 519910 67351 519966 67360
rect 519266 66464 519322 66473
rect 519266 66399 519322 66408
rect 519818 65920 519874 65929
rect 519818 65855 519874 65864
rect 116596 64846 116716 64874
rect 116596 64734 116624 64846
rect 116584 64728 116636 64734
rect 116584 64670 116636 64676
rect 116214 64560 116270 64569
rect 116214 64495 116270 64504
rect 116228 63578 116256 64495
rect 519082 64424 519138 64433
rect 519082 64359 519138 64368
rect 116216 63572 116268 63578
rect 116216 63514 116268 63520
rect 116122 62656 116178 62665
rect 116122 62591 116178 62600
rect 116136 62150 116164 62591
rect 116124 62144 116176 62150
rect 116124 62086 116176 62092
rect 519096 61033 519124 64359
rect 519832 62393 519860 65855
rect 519924 63753 519952 67351
rect 520200 65113 520228 68711
rect 520186 65104 520242 65113
rect 520186 65039 520242 65048
rect 519910 63744 519966 63753
rect 519910 63679 519966 63688
rect 520094 62928 520150 62937
rect 520094 62863 520150 62872
rect 519818 62384 519874 62393
rect 519818 62319 519874 62328
rect 519082 61024 519138 61033
rect 519082 60959 519138 60968
rect 519082 59936 519138 59945
rect 519082 59871 519138 59880
rect 116582 58712 116638 58721
rect 116582 58647 116638 58656
rect 114190 53136 114246 53145
rect 114190 53071 114246 53080
rect 116122 45248 116178 45257
rect 116122 45183 116178 45192
rect 116136 44198 116164 45183
rect 116124 44192 116176 44198
rect 116124 44134 116176 44140
rect 114098 41848 114154 41857
rect 114098 41783 114154 41792
rect 115202 39536 115258 39545
rect 115202 39471 115258 39480
rect 114100 33176 114152 33182
rect 114100 33118 114152 33124
rect 114006 30424 114062 30433
rect 114006 30359 114062 30368
rect 114008 23520 114060 23526
rect 114008 23462 114060 23468
rect 113914 19000 113970 19009
rect 113914 18935 113970 18944
rect 113822 7712 113878 7721
rect 113822 7647 113878 7656
rect 112904 1148 112956 1154
rect 112904 1090 112956 1096
rect 114020 1086 114048 23462
rect 114008 1080 114060 1086
rect 114008 1022 114060 1028
rect 112812 1012 112864 1018
rect 112812 954 112864 960
rect 112720 876 112772 882
rect 112720 818 112772 824
rect 114112 746 114140 33118
rect 114100 740 114152 746
rect 114100 682 114152 688
rect 112628 604 112680 610
rect 112628 546 112680 552
rect 115216 474 115244 39471
rect 115938 35728 115994 35737
rect 115938 35663 115994 35672
rect 115952 34542 115980 35663
rect 115940 34536 115992 34542
rect 115940 34478 115992 34484
rect 115938 33824 115994 33833
rect 115938 33759 115994 33768
rect 115952 33182 115980 33759
rect 115940 33176 115992 33182
rect 115940 33118 115992 33124
rect 115294 31784 115350 31793
rect 115294 31719 115350 31728
rect 115308 610 115336 31719
rect 116122 29880 116178 29889
rect 116122 29815 116178 29824
rect 116136 29034 116164 29815
rect 116124 29028 116176 29034
rect 116124 28970 116176 28976
rect 115386 27976 115442 27985
rect 115386 27911 115442 27920
rect 115400 814 115428 27911
rect 116122 26072 116178 26081
rect 116122 26007 116178 26016
rect 116136 24886 116164 26007
rect 116124 24880 116176 24886
rect 116124 24822 116176 24828
rect 115938 24168 115994 24177
rect 115938 24103 115994 24112
rect 115952 23526 115980 24103
rect 115940 23520 115992 23526
rect 115940 23462 115992 23468
rect 116122 22264 116178 22273
rect 116122 22199 116178 22208
rect 116136 22166 116164 22199
rect 116124 22160 116176 22166
rect 116124 22102 116176 22108
rect 116490 14512 116546 14521
rect 116490 14447 116546 14456
rect 116214 12608 116270 12617
rect 116214 12543 116270 12552
rect 116032 11688 116084 11694
rect 116032 11630 116084 11636
rect 115938 6896 115994 6905
rect 115938 6831 115994 6840
rect 115952 5574 115980 6831
rect 115940 5568 115992 5574
rect 115940 5510 115992 5516
rect 116044 5250 116072 11630
rect 116122 10704 116178 10713
rect 116122 10639 116178 10648
rect 115952 5222 116072 5250
rect 115952 1426 115980 5222
rect 116136 5114 116164 10639
rect 116044 5086 116164 5114
rect 116044 1737 116072 5086
rect 116122 4992 116178 5001
rect 116122 4927 116178 4936
rect 116136 4214 116164 4927
rect 116124 4208 116176 4214
rect 116124 4150 116176 4156
rect 116122 3088 116178 3097
rect 116122 3023 116178 3032
rect 116030 1728 116086 1737
rect 116030 1663 116086 1672
rect 115940 1420 115992 1426
rect 115940 1362 115992 1368
rect 116136 1358 116164 3023
rect 116228 1873 116256 12543
rect 116400 11756 116452 11762
rect 116400 11698 116452 11704
rect 116214 1864 116270 1873
rect 116214 1799 116270 1808
rect 116412 1494 116440 11698
rect 116504 2009 116532 14447
rect 116490 2000 116546 2009
rect 116596 1970 116624 58647
rect 519096 56953 519124 59871
rect 520108 59673 520136 62863
rect 520186 61432 520242 61441
rect 520186 61367 520242 61376
rect 520094 59664 520150 59673
rect 520094 59599 520150 59608
rect 520002 58440 520058 58449
rect 520002 58375 520058 58384
rect 519082 56944 519138 56953
rect 519082 56879 519138 56888
rect 519450 56944 519506 56953
rect 519450 56879 519506 56888
rect 116674 56808 116730 56817
rect 116674 56743 116730 56752
rect 116490 1935 116546 1944
rect 116584 1964 116636 1970
rect 116584 1906 116636 1912
rect 116688 1766 116716 56743
rect 519464 54233 519492 56879
rect 520016 55593 520044 58375
rect 520200 58313 520228 61367
rect 520186 58304 520242 58313
rect 520186 58239 520242 58248
rect 520002 55584 520058 55593
rect 520002 55519 520058 55528
rect 519818 55448 519874 55457
rect 519818 55383 519874 55392
rect 519450 54224 519506 54233
rect 519450 54159 519506 54168
rect 116766 53000 116822 53009
rect 116766 52935 116822 52944
rect 116780 3641 116808 52935
rect 519832 52873 519860 55383
rect 520002 54088 520058 54097
rect 520002 54023 520058 54032
rect 519818 52864 519874 52873
rect 519818 52799 519874 52808
rect 520016 51513 520044 54023
rect 520094 52592 520150 52601
rect 520094 52527 520150 52536
rect 520002 51504 520058 51513
rect 520002 51439 520058 51448
rect 520108 50153 520136 52527
rect 520186 51096 520242 51105
rect 520186 51031 520242 51040
rect 520094 50144 520150 50153
rect 520094 50079 520150 50088
rect 520200 48793 520228 51031
rect 521106 49600 521162 49609
rect 521106 49535 521162 49544
rect 520186 48784 520242 48793
rect 520186 48719 520242 48728
rect 520922 48104 520978 48113
rect 520922 48039 520978 48048
rect 520936 46753 520964 48039
rect 521120 47433 521148 49535
rect 521106 47424 521162 47433
rect 521106 47359 521162 47368
rect 520922 46744 520978 46753
rect 520922 46679 520978 46688
rect 521566 46608 521622 46617
rect 521566 46543 521622 46552
rect 521580 45665 521608 46543
rect 521566 45656 521622 45665
rect 521566 45591 521622 45600
rect 521106 45112 521162 45121
rect 521106 45047 521162 45056
rect 521120 44033 521148 45047
rect 521106 44024 521162 44033
rect 521106 43959 521162 43968
rect 520922 43616 520978 43625
rect 520922 43551 520978 43560
rect 520936 42673 520964 43551
rect 520922 42664 520978 42673
rect 520922 42599 520978 42608
rect 521106 42120 521162 42129
rect 521106 42055 521162 42064
rect 116950 41440 117006 41449
rect 116950 41375 117006 41384
rect 116858 20360 116914 20369
rect 116858 20295 116914 20304
rect 116872 11762 116900 20295
rect 116860 11756 116912 11762
rect 116860 11698 116912 11704
rect 116964 6914 116992 41375
rect 521120 41313 521148 42055
rect 521106 41304 521162 41313
rect 521106 41239 521162 41248
rect 521106 40760 521162 40769
rect 521106 40695 521162 40704
rect 521120 39953 521148 40695
rect 521106 39944 521162 39953
rect 521106 39879 521162 39888
rect 521106 39264 521162 39273
rect 521106 39199 521162 39208
rect 521120 37913 521148 39199
rect 521106 37904 521162 37913
rect 521106 37839 521162 37848
rect 117134 37632 117190 37641
rect 117134 37567 117190 37576
rect 117042 18456 117098 18465
rect 117042 18391 117098 18400
rect 117056 11694 117084 18391
rect 117044 11688 117096 11694
rect 117044 11630 117096 11636
rect 117042 8800 117098 8809
rect 117042 8735 117098 8744
rect 116872 6886 116992 6914
rect 116872 3777 116900 6886
rect 116858 3768 116914 3777
rect 116858 3703 116914 3712
rect 116766 3632 116822 3641
rect 116766 3567 116822 3576
rect 116676 1760 116728 1766
rect 116676 1702 116728 1708
rect 117056 1601 117084 8735
rect 117148 3505 117176 37567
rect 520922 30288 520978 30297
rect 520922 30223 520978 30232
rect 520936 29073 520964 30223
rect 520922 29064 520978 29073
rect 520922 28999 520978 29008
rect 521106 28792 521162 28801
rect 521106 28727 521162 28736
rect 521120 27713 521148 28727
rect 521106 27704 521162 27713
rect 521106 27639 521162 27648
rect 521106 27432 521162 27441
rect 521106 27367 521162 27376
rect 521120 26353 521148 27367
rect 521106 26344 521162 26353
rect 521106 26279 521162 26288
rect 520922 25936 520978 25945
rect 520922 25871 520978 25880
rect 520936 24993 520964 25871
rect 520922 24984 520978 24993
rect 520922 24919 520978 24928
rect 519082 24440 519138 24449
rect 519082 24375 519138 24384
rect 519096 23633 519124 24375
rect 519082 23624 519138 23633
rect 519082 23559 519138 23568
rect 521106 22944 521162 22953
rect 521106 22879 521162 22888
rect 521120 22273 521148 22879
rect 521106 22264 521162 22273
rect 521106 22199 521162 22208
rect 117226 16416 117282 16425
rect 117226 16351 117282 16360
rect 117134 3496 117190 3505
rect 117134 3431 117190 3440
rect 117240 2145 117268 16351
rect 521106 10704 521162 10713
rect 521106 10639 521162 10648
rect 521120 9625 521148 10639
rect 521106 9616 521162 9625
rect 521106 9551 521162 9560
rect 520922 9344 520978 9353
rect 520922 9279 520978 9288
rect 520936 8129 520964 9279
rect 520922 8120 520978 8129
rect 520922 8055 520978 8064
rect 520278 7984 520334 7993
rect 520278 7919 520334 7928
rect 520292 6633 520320 7919
rect 520278 6624 520334 6633
rect 520278 6559 520334 6568
rect 521106 6488 521162 6497
rect 521106 6423 521162 6432
rect 521014 5264 521070 5273
rect 521014 5199 521070 5208
rect 521028 3641 521056 5199
rect 521120 5137 521148 6423
rect 521106 5128 521162 5137
rect 521106 5063 521162 5072
rect 521198 3904 521254 3913
rect 521198 3839 521254 3848
rect 521014 3632 521070 3641
rect 521014 3567 521070 3576
rect 521106 2680 521162 2689
rect 521106 2615 521162 2624
rect 143644 2514 143980 2530
rect 443656 2514 443992 2530
rect 143632 2508 143980 2514
rect 143684 2502 143980 2508
rect 425796 2508 425848 2514
rect 143632 2450 143684 2456
rect 425796 2450 425848 2456
rect 443644 2508 443992 2514
rect 443696 2502 443992 2508
rect 443644 2450 443696 2456
rect 117226 2136 117282 2145
rect 117226 2071 117282 2080
rect 193600 2094 193936 2122
rect 243648 2094 243984 2122
rect 293604 2094 293940 2122
rect 343652 2094 343988 2122
rect 393608 2094 393944 2122
rect 117042 1592 117098 1601
rect 117042 1527 117098 1536
rect 163778 1592 163834 1601
rect 193600 1562 193628 2094
rect 229282 1728 229338 1737
rect 229282 1663 229338 1672
rect 163778 1527 163834 1536
rect 193588 1556 193640 1562
rect 116400 1488 116452 1494
rect 116400 1430 116452 1436
rect 116124 1352 116176 1358
rect 116124 1294 116176 1300
rect 115388 808 115440 814
rect 163792 800 163820 1527
rect 193588 1498 193640 1504
rect 229296 800 229324 1663
rect 243648 1601 243676 2094
rect 293604 1737 293632 2094
rect 293590 1728 293646 1737
rect 293590 1663 293646 1672
rect 243634 1592 243690 1601
rect 243634 1527 243690 1536
rect 294786 1456 294842 1465
rect 343652 1426 343680 2094
rect 393608 1465 393636 2094
rect 360290 1456 360346 1465
rect 294786 1391 294788 1400
rect 294840 1391 294842 1400
rect 343640 1420 343692 1426
rect 294788 1362 294840 1368
rect 360290 1391 360346 1400
rect 393594 1456 393650 1465
rect 393594 1391 393650 1400
rect 343640 1362 343692 1368
rect 294800 800 294828 1362
rect 360304 800 360332 1391
rect 425808 800 425836 2450
rect 493612 2094 493948 2122
rect 493612 1426 493640 2094
rect 491300 1420 491352 1426
rect 491300 1362 491352 1368
rect 493600 1420 493652 1426
rect 493600 1362 493652 1368
rect 491312 800 491340 1362
rect 115388 750 115440 756
rect 115296 604 115348 610
rect 115296 546 115348 552
rect 115204 468 115256 474
rect 115204 410 115256 416
rect 112536 400 112588 406
rect 112536 342 112588 348
rect 163778 -400 163834 800
rect 229282 -400 229338 800
rect 294786 -400 294842 800
rect 360290 -400 360346 800
rect 425794 -400 425850 800
rect 491298 -400 491354 800
rect 521120 785 521148 2615
rect 521212 2145 521240 3839
rect 521198 2136 521254 2145
rect 521198 2071 521254 2080
rect 521106 776 521162 785
rect 521106 711 521162 720
<< via2 >>
rect 2870 155080 2926 155136
rect 2042 153720 2098 153776
rect 2686 151816 2742 151872
rect 8298 156032 8354 156088
rect 9586 155216 9642 155272
rect 6182 152360 6238 152416
rect 9494 151408 9550 151464
rect 16302 155488 16358 155544
rect 18786 152496 18842 152552
rect 16394 151952 16450 152008
rect 12990 150592 13046 150648
rect 23018 155624 23074 155680
rect 20534 153856 20590 153912
rect 19614 152632 19670 152688
rect 28906 155896 28962 155952
rect 29734 155760 29790 155816
rect 33966 156576 34022 156632
rect 44822 153992 44878 154048
rect 61658 154128 61714 154184
rect 37002 152088 37058 152144
rect 33598 151544 33654 151600
rect 30194 151136 30250 151192
rect 23294 150864 23350 150920
rect 19798 150728 19854 150784
rect 67546 151000 67602 151056
rect 91834 156712 91890 156768
rect 91098 153040 91154 153096
rect 93582 152768 93638 152824
rect 98642 154264 98698 154320
rect 101954 156848 102010 156904
rect 104438 156984 104494 157040
rect 107750 155388 107752 155408
rect 107752 155388 107804 155408
rect 107804 155388 107806 155408
rect 107750 155352 107806 155388
rect 109038 155388 109040 155408
rect 109040 155388 109092 155408
rect 109092 155388 109094 155408
rect 108670 154400 108726 154456
rect 109038 155352 109094 155388
rect 109130 152904 109186 152960
rect 109038 152224 109094 152280
rect 109866 152088 109922 152144
rect 109682 151816 109738 151872
rect 109222 150456 109278 150512
rect 80610 149640 80666 149696
rect 64694 149504 64750 149560
rect 26974 149368 27030 149424
rect 57886 149368 57942 149424
rect 61474 149368 61530 149424
rect 109774 150728 109830 150784
rect 110878 151408 110934 151464
rect 110970 150864 111026 150920
rect 111338 150592 111394 150648
rect 111154 150456 111210 150512
rect 110326 140800 110382 140856
rect 110326 113192 110382 113248
rect 110326 110608 110382 110664
rect 110326 107616 110382 107672
rect 110326 98096 110382 98152
rect 113178 154844 113180 154864
rect 113180 154844 113232 154864
rect 113232 154844 113234 154864
rect 113178 154808 113234 154844
rect 112902 154672 112958 154728
rect 113454 154672 113510 154728
rect 113638 154672 113694 154728
rect 112442 151544 112498 151600
rect 111706 151272 111762 151328
rect 111706 151136 111762 151192
rect 115938 154808 115994 154864
rect 116214 151952 116270 152008
rect 115846 151136 115902 151192
rect 112902 149504 112958 149560
rect 112718 149368 112774 149424
rect 112534 149232 112590 149288
rect 113822 144200 113878 144256
rect 110326 88304 110382 88360
rect 113914 132776 113970 132832
rect 116122 148996 116124 149016
rect 116124 148996 116176 149016
rect 116176 148996 116178 149016
rect 116122 148960 116178 148996
rect 116030 145152 116086 145208
rect 116122 143248 116178 143304
rect 116122 139440 116178 139496
rect 116122 137536 116178 137592
rect 115938 131688 115994 131744
rect 115938 129784 115994 129840
rect 115202 127880 115258 127936
rect 116122 125976 116178 126032
rect 116122 124108 116124 124128
rect 116124 124108 116176 124128
rect 116176 124108 116178 124128
rect 116122 124072 116178 124108
rect 116122 122168 116178 122224
rect 114006 121352 114062 121408
rect 116122 120128 116178 120184
rect 114098 110064 114154 110120
rect 116122 106800 116178 106856
rect 116122 104796 116124 104816
rect 116124 104796 116176 104816
rect 116176 104796 116178 104816
rect 116122 104760 116178 104796
rect 115938 100952 115994 101008
rect 114190 98640 114246 98696
rect 116398 149640 116454 149696
rect 116858 154692 116914 154728
rect 116858 154672 116860 154692
rect 116860 154672 116912 154692
rect 116912 154672 116914 154692
rect 116582 151408 116638 151464
rect 116582 149096 116638 149152
rect 116490 147056 116546 147112
rect 116214 97144 116270 97200
rect 116122 95240 116178 95296
rect 116122 93336 116178 93392
rect 118790 153584 118846 153640
rect 120446 155352 120502 155408
rect 121090 155080 121146 155136
rect 120446 153720 120502 153776
rect 123666 152360 123722 152416
rect 124954 156032 125010 156088
rect 126242 155216 126298 155272
rect 125598 152224 125654 152280
rect 126334 152224 126390 152280
rect 131118 155896 131174 155952
rect 131026 155488 131082 155544
rect 130750 153040 130806 153096
rect 132958 155252 132960 155272
rect 132960 155252 133012 155272
rect 133012 155252 133014 155272
rect 132958 155216 133014 155252
rect 134522 155624 134578 155680
rect 131118 153040 131174 153096
rect 134614 153856 134670 153912
rect 133970 152632 134026 152688
rect 134522 152632 134578 152688
rect 133234 152496 133290 152552
rect 133326 152360 133382 152416
rect 136914 154808 136970 154864
rect 136546 152632 136602 152688
rect 138018 155760 138074 155816
rect 137374 155252 137376 155272
rect 137376 155252 137428 155272
rect 137428 155252 137430 155272
rect 137374 155216 137430 155252
rect 137558 154844 137560 154864
rect 137560 154844 137612 154864
rect 137612 154844 137614 154864
rect 137558 154808 137614 154844
rect 138938 153720 138994 153776
rect 140594 155216 140650 155272
rect 141054 153040 141110 153096
rect 145194 156576 145250 156632
rect 147310 155488 147366 155544
rect 153198 153992 153254 154048
rect 162858 152904 162914 152960
rect 164238 153856 164294 153912
rect 166078 154128 166134 154184
rect 170586 151000 170642 151056
rect 173438 155796 173440 155816
rect 173440 155796 173492 155816
rect 173492 155796 173494 155816
rect 173438 155760 173494 155796
rect 175830 155796 175832 155816
rect 175832 155796 175884 155816
rect 175884 155796 175886 155816
rect 175830 155760 175886 155796
rect 184662 151408 184718 151464
rect 189170 156712 189226 156768
rect 190826 154672 190882 154728
rect 190458 152768 190514 152824
rect 191838 152632 191894 152688
rect 192022 154672 192078 154728
rect 193218 154264 193274 154320
rect 194322 154128 194378 154184
rect 196806 156848 196862 156904
rect 198830 156984 198886 157040
rect 200118 153856 200174 153912
rect 202050 154400 202106 154456
rect 201866 153856 201922 153912
rect 200210 152768 200266 152824
rect 203982 151272 204038 151328
rect 205270 153992 205326 154048
rect 207754 155624 207810 155680
rect 206098 154128 206154 154184
rect 207202 151136 207258 151192
rect 208674 155352 208730 155408
rect 209778 153584 209834 153640
rect 211894 154964 211950 155000
rect 211894 154944 211896 154964
rect 211896 154944 211948 154964
rect 211948 154944 211950 154964
rect 212538 154964 212594 155000
rect 212538 154944 212540 154964
rect 212540 154944 212592 154964
rect 212592 154944 212594 154964
rect 214470 155352 214526 155408
rect 215482 152360 215538 152416
rect 218058 154264 218114 154320
rect 217874 152360 217930 152416
rect 220726 154264 220782 154320
rect 218702 152496 218758 152552
rect 222566 155488 222622 155544
rect 222750 155488 222806 155544
rect 222566 155080 222622 155136
rect 220818 152496 220874 152552
rect 223578 155488 223634 155544
rect 223578 155216 223634 155272
rect 225142 153720 225198 153776
rect 227902 155216 227958 155272
rect 227810 155080 227866 155136
rect 229650 153720 229706 153776
rect 232042 154964 232098 155000
rect 232042 154944 232044 154964
rect 232044 154944 232096 154964
rect 232096 154944 232098 154964
rect 233238 154944 233294 155000
rect 233514 154264 233570 154320
rect 238574 154828 238630 154864
rect 238574 154808 238576 154828
rect 238576 154808 238628 154828
rect 238628 154808 238630 154828
rect 239034 154828 239090 154864
rect 239034 154808 239036 154828
rect 239036 154808 239088 154828
rect 239088 154808 239090 154828
rect 240414 155488 240470 155544
rect 242990 155488 243046 155544
rect 254766 155488 254822 155544
rect 260562 155080 260618 155136
rect 262402 154400 262458 154456
rect 263690 155080 263746 155136
rect 264978 152632 265034 152688
rect 265714 154264 265770 154320
rect 266450 152632 266506 152688
rect 270222 153040 270278 153096
rect 269486 152768 269542 152824
rect 273350 155624 273406 155680
rect 273258 153856 273314 153912
rect 272706 153040 272762 153096
rect 274914 155624 274970 155680
rect 275742 153992 275798 154048
rect 273350 151816 273406 151872
rect 276478 154128 276534 154184
rect 275834 153856 275890 153912
rect 278686 153992 278742 154048
rect 279514 155352 279570 155408
rect 278318 152768 278374 152824
rect 277766 151816 277822 151872
rect 279882 154980 279884 155000
rect 279884 154980 279936 155000
rect 279936 154980 279938 155000
rect 279882 154944 279938 154980
rect 282918 154944 282974 155000
rect 285494 152360 285550 152416
rect 286874 153176 286930 153232
rect 287058 152360 287114 152416
rect 287426 152496 287482 152552
rect 291474 153212 291476 153232
rect 291476 153212 291528 153232
rect 291528 153212 291530 153232
rect 291474 153176 291530 153212
rect 292394 154964 292450 155000
rect 292394 154944 292396 154964
rect 292396 154944 292448 154964
rect 292448 154944 292450 154964
rect 292302 154128 292358 154184
rect 293222 155216 293278 155272
rect 292670 154128 292726 154184
rect 292854 154128 292910 154184
rect 293958 154944 294014 155000
rect 295154 155216 295210 155272
rect 294510 153720 294566 153776
rect 299570 155372 299626 155408
rect 299570 155352 299572 155372
rect 299572 155352 299624 155372
rect 299624 155352 299626 155372
rect 299662 154808 299718 154864
rect 299662 154128 299718 154184
rect 303526 154808 303582 154864
rect 309138 155352 309194 155408
rect 310610 155488 310666 155544
rect 311438 154944 311494 155000
rect 311898 155488 311954 155544
rect 311714 155352 311770 155408
rect 312082 155352 312138 155408
rect 311806 154944 311862 155000
rect 312266 153992 312322 154048
rect 311714 153312 311770 153368
rect 311898 153312 311954 153368
rect 312358 153584 312414 153640
rect 312910 153584 312966 153640
rect 316774 155488 316830 155544
rect 316222 153212 316224 153232
rect 316224 153212 316276 153232
rect 316276 153212 316278 153232
rect 316222 153176 316278 153212
rect 317142 153212 317144 153232
rect 317144 153212 317196 153232
rect 317196 153212 317198 153232
rect 317142 153176 317198 153212
rect 319534 154400 319590 154456
rect 320178 153720 320234 153776
rect 320270 153040 320326 153096
rect 321834 154964 321890 155000
rect 321834 154944 321836 154964
rect 321836 154944 321888 154964
rect 321888 154944 321890 154964
rect 322202 154964 322258 155000
rect 322202 154944 322204 154964
rect 322204 154944 322256 154964
rect 322256 154944 322258 154964
rect 322110 154264 322166 154320
rect 321466 152632 321522 152688
rect 323398 153040 323454 153096
rect 325238 153448 325294 153504
rect 326066 154572 326068 154592
rect 326068 154572 326120 154592
rect 326120 154572 326122 154592
rect 326066 154536 326122 154572
rect 329194 155624 329250 155680
rect 327630 154536 327686 154592
rect 327538 153448 327594 153504
rect 328642 153176 328698 153232
rect 329838 153856 329894 153912
rect 331218 154264 331274 154320
rect 331770 152768 331826 152824
rect 332782 153176 332838 153232
rect 336186 154284 336242 154320
rect 336186 154264 336188 154284
rect 336188 154264 336240 154284
rect 336240 154264 336242 154284
rect 337014 153348 337016 153368
rect 337016 153348 337068 153368
rect 337068 153348 337070 153368
rect 337014 153312 337070 153348
rect 336830 152360 336886 152416
rect 338118 153720 338174 153776
rect 340234 154808 340290 154864
rect 340326 154672 340382 154728
rect 340510 154964 340566 155000
rect 340510 154944 340512 154964
rect 340512 154944 340564 154964
rect 340564 154944 340566 154964
rect 339406 153312 339462 153368
rect 340878 154808 340934 154864
rect 342166 155216 342222 155272
rect 341246 154944 341302 155000
rect 342810 154672 342866 154728
rect 342718 154264 342774 154320
rect 342902 153348 342904 153368
rect 342904 153348 342956 153368
rect 342956 153348 342958 153368
rect 342902 153312 342958 153348
rect 345386 153348 345388 153368
rect 345388 153348 345440 153368
rect 345440 153348 345442 153368
rect 345386 153312 345442 153348
rect 345754 154284 345810 154320
rect 345754 154264 345756 154284
rect 345756 154264 345808 154284
rect 345808 154264 345810 154284
rect 348790 155080 348846 155136
rect 349894 155216 349950 155272
rect 354586 155216 354642 155272
rect 354218 155080 354274 155136
rect 432878 152360 432934 152416
rect 449898 152360 449954 152416
rect 519542 157664 519598 157720
rect 519634 156168 519690 156224
rect 519542 147872 519598 147928
rect 520922 159160 520978 159216
rect 519726 154672 519782 154728
rect 519634 146512 519690 146568
rect 519818 153176 519874 153232
rect 519726 145152 519782 145208
rect 519910 150184 519966 150240
rect 519818 143792 519874 143848
rect 521014 151680 521070 151736
rect 520922 149232 520978 149288
rect 520922 145832 520978 145888
rect 520278 144336 520334 144392
rect 519910 141072 519966 141128
rect 520738 142840 520794 142896
rect 520278 135632 520334 135688
rect 117226 135496 117282 135552
rect 521106 148688 521162 148744
rect 521014 142432 521070 142488
rect 521014 141344 521070 141400
rect 520922 136992 520978 137048
rect 520738 134272 520794 134328
rect 520278 134000 520334 134056
rect 117134 133592 117190 133648
rect 520186 131008 520242 131064
rect 519910 129512 519966 129568
rect 519542 128016 519598 128072
rect 519266 123528 519322 123584
rect 117042 118224 117098 118280
rect 519726 126520 519782 126576
rect 519542 120672 519598 120728
rect 519818 125024 519874 125080
rect 519726 119312 519782 119368
rect 521198 147328 521254 147384
rect 521106 139712 521162 139768
rect 521290 139848 521346 139904
rect 521198 138352 521254 138408
rect 521198 136856 521254 136912
rect 521106 135360 521162 135416
rect 521014 132912 521070 132968
rect 521014 132504 521070 132560
rect 520278 126112 520334 126168
rect 521382 138352 521438 138408
rect 521290 131552 521346 131608
rect 521382 130192 521438 130248
rect 521198 128832 521254 128888
rect 521106 127472 521162 127528
rect 521014 124752 521070 124808
rect 520186 123392 520242 123448
rect 519910 122032 519966 122088
rect 520094 122032 520150 122088
rect 519910 119176 519966 119232
rect 519818 117952 519874 118008
rect 519726 117680 519782 117736
rect 519266 116592 519322 116648
rect 116950 116320 117006 116376
rect 519266 113192 519322 113248
rect 116858 112512 116914 112568
rect 519818 114688 519874 114744
rect 519726 111152 519782 111208
rect 519634 108704 519690 108760
rect 519266 107072 519322 107128
rect 519082 104352 519138 104408
rect 116766 102856 116822 102912
rect 520002 116184 520058 116240
rect 519910 112512 519966 112568
rect 520186 120672 520242 120728
rect 520094 115232 520150 115288
rect 520186 113872 520242 113928
rect 520094 111696 520150 111752
rect 520002 109792 520058 109848
rect 519818 108432 519874 108488
rect 519726 107344 519782 107400
rect 519634 102992 519690 103048
rect 519910 105848 519966 105904
rect 519726 101632 519782 101688
rect 520186 110200 520242 110256
rect 520094 105712 520150 105768
rect 520186 104488 520242 104544
rect 520094 102856 520150 102912
rect 519910 100272 519966 100328
rect 519450 99864 519506 99920
rect 519082 98912 519138 98968
rect 519818 98368 519874 98424
rect 519542 96872 519598 96928
rect 519450 94832 519506 94888
rect 519082 94016 519138 94072
rect 116582 91296 116638 91352
rect 519266 92520 519322 92576
rect 519082 89392 519138 89448
rect 519726 95376 519782 95432
rect 519542 92112 519598 92168
rect 519450 91024 519506 91080
rect 519266 88032 519322 88088
rect 115938 87488 115994 87544
rect 114282 87216 114338 87272
rect 116398 85584 116454 85640
rect 520186 101360 520242 101416
rect 520094 97552 520150 97608
rect 520186 96192 520242 96248
rect 519818 93472 519874 93528
rect 519726 90752 519782 90808
rect 519910 89528 519966 89584
rect 519726 86536 519782 86592
rect 519450 85312 519506 85368
rect 519082 85040 519138 85096
rect 116582 83680 116638 83736
rect 116306 81776 116362 81832
rect 520002 88032 520058 88088
rect 519910 83952 519966 84008
rect 521566 86672 521622 86728
rect 520094 83544 520150 83600
rect 520002 82592 520058 82648
rect 519726 81232 519782 81288
rect 115938 79872 115994 79928
rect 519082 79872 519138 79928
rect 520186 82048 520242 82104
rect 520094 78512 520150 78568
rect 116214 77968 116270 78024
rect 521106 80688 521162 80744
rect 520554 79192 520610 79248
rect 520186 77152 520242 77208
rect 521014 77696 521070 77752
rect 520554 74568 520610 74624
rect 116674 74024 116730 74080
rect 116582 72120 116638 72176
rect 113362 64504 113418 64560
rect 110326 59336 110382 59392
rect 109406 3576 109462 3632
rect 109498 3440 109554 3496
rect 109406 3168 109462 3224
rect 33046 2624 33102 2680
rect 76194 2624 76250 2680
rect 88890 2624 88946 2680
rect 98274 2624 98330 2680
rect 100298 2624 100354 2680
rect 102138 2624 102194 2680
rect 102322 2624 102378 2680
rect 26054 2080 26110 2136
rect 22926 1944 22982 2000
rect 19338 1808 19394 1864
rect 15934 1672 15990 1728
rect 12622 1536 12678 1592
rect 55954 1400 56010 1456
rect 94410 2352 94466 2408
rect 98274 2216 98330 2272
rect 102138 2352 102194 2408
rect 109498 2216 109554 2272
rect 110326 53896 110382 53952
rect 110326 51040 110382 51096
rect 110326 48320 110382 48376
rect 110326 47096 110382 47152
rect 110326 42880 110382 42936
rect 110142 3984 110198 4040
rect 110142 2896 110198 2952
rect 111062 2796 111064 2816
rect 111064 2796 111116 2816
rect 111116 2796 111118 2816
rect 111062 2760 111118 2796
rect 98274 1264 98330 1320
rect 102322 1264 102378 1320
rect 116306 70216 116362 70272
rect 116122 68312 116178 68368
rect 116582 66408 116638 66464
rect 521198 76200 521254 76256
rect 521106 75928 521162 75984
rect 521106 74704 521162 74760
rect 521014 73752 521070 73808
rect 521014 73208 521070 73264
rect 520002 71712 520058 71768
rect 519266 70216 519322 70272
rect 521198 71848 521254 71904
rect 521106 70488 521162 70544
rect 521014 69128 521070 69184
rect 520186 68720 520242 68776
rect 520002 67768 520058 67824
rect 519910 67360 519966 67416
rect 519266 66408 519322 66464
rect 519818 65864 519874 65920
rect 116214 64504 116270 64560
rect 519082 64368 519138 64424
rect 116122 62600 116178 62656
rect 520186 65048 520242 65104
rect 519910 63688 519966 63744
rect 520094 62872 520150 62928
rect 519818 62328 519874 62384
rect 519082 60968 519138 61024
rect 519082 59880 519138 59936
rect 116582 58656 116638 58712
rect 114190 53080 114246 53136
rect 116122 45192 116178 45248
rect 114098 41792 114154 41848
rect 115202 39480 115258 39536
rect 114006 30368 114062 30424
rect 113914 18944 113970 19000
rect 113822 7656 113878 7712
rect 115938 35672 115994 35728
rect 115938 33768 115994 33824
rect 115294 31728 115350 31784
rect 116122 29824 116178 29880
rect 115386 27920 115442 27976
rect 116122 26016 116178 26072
rect 115938 24112 115994 24168
rect 116122 22208 116178 22264
rect 116490 14456 116546 14512
rect 116214 12552 116270 12608
rect 115938 6840 115994 6896
rect 116122 10648 116178 10704
rect 116122 4936 116178 4992
rect 116122 3032 116178 3088
rect 116030 1672 116086 1728
rect 116214 1808 116270 1864
rect 116490 1944 116546 2000
rect 520186 61376 520242 61432
rect 520094 59608 520150 59664
rect 520002 58384 520058 58440
rect 519082 56888 519138 56944
rect 519450 56888 519506 56944
rect 116674 56752 116730 56808
rect 520186 58248 520242 58304
rect 520002 55528 520058 55584
rect 519818 55392 519874 55448
rect 519450 54168 519506 54224
rect 116766 52944 116822 53000
rect 520002 54032 520058 54088
rect 519818 52808 519874 52864
rect 520094 52536 520150 52592
rect 520002 51448 520058 51504
rect 520186 51040 520242 51096
rect 520094 50088 520150 50144
rect 521106 49544 521162 49600
rect 520186 48728 520242 48784
rect 520922 48048 520978 48104
rect 521106 47368 521162 47424
rect 520922 46688 520978 46744
rect 521566 46552 521622 46608
rect 521566 45600 521622 45656
rect 521106 45056 521162 45112
rect 521106 43968 521162 44024
rect 520922 43560 520978 43616
rect 520922 42608 520978 42664
rect 521106 42064 521162 42120
rect 116950 41384 117006 41440
rect 116858 20304 116914 20360
rect 521106 41248 521162 41304
rect 521106 40704 521162 40760
rect 521106 39888 521162 39944
rect 521106 39208 521162 39264
rect 521106 37848 521162 37904
rect 117134 37576 117190 37632
rect 117042 18400 117098 18456
rect 117042 8744 117098 8800
rect 116858 3712 116914 3768
rect 116766 3576 116822 3632
rect 520922 30232 520978 30288
rect 520922 29008 520978 29064
rect 521106 28736 521162 28792
rect 521106 27648 521162 27704
rect 521106 27376 521162 27432
rect 521106 26288 521162 26344
rect 520922 25880 520978 25936
rect 520922 24928 520978 24984
rect 519082 24384 519138 24440
rect 519082 23568 519138 23624
rect 521106 22888 521162 22944
rect 521106 22208 521162 22264
rect 117226 16360 117282 16416
rect 117134 3440 117190 3496
rect 521106 10648 521162 10704
rect 521106 9560 521162 9616
rect 520922 9288 520978 9344
rect 520922 8064 520978 8120
rect 520278 7928 520334 7984
rect 520278 6568 520334 6624
rect 521106 6432 521162 6488
rect 521014 5208 521070 5264
rect 521106 5072 521162 5128
rect 521198 3848 521254 3904
rect 521014 3576 521070 3632
rect 521106 2624 521162 2680
rect 117226 2080 117282 2136
rect 117042 1536 117098 1592
rect 163778 1536 163834 1592
rect 229282 1672 229338 1728
rect 293590 1672 293646 1728
rect 243634 1536 243690 1592
rect 294786 1420 294842 1456
rect 294786 1400 294788 1420
rect 294788 1400 294840 1420
rect 294840 1400 294842 1420
rect 360290 1400 360346 1456
rect 393594 1400 393650 1456
rect 521198 2080 521254 2136
rect 521106 720 521162 776
<< metal3 >>
rect 520917 159218 520983 159221
rect 523200 159218 524400 159248
rect 520917 159216 524400 159218
rect 520917 159160 520922 159216
rect 520978 159160 524400 159216
rect 520917 159158 524400 159160
rect 520917 159155 520983 159158
rect 523200 159128 524400 159158
rect 519537 157722 519603 157725
rect 523200 157722 524400 157752
rect 519537 157720 524400 157722
rect 519537 157664 519542 157720
rect 519598 157664 524400 157720
rect 519537 157662 524400 157664
rect 519537 157659 519603 157662
rect 523200 157632 524400 157662
rect 104433 157042 104499 157045
rect 198825 157042 198891 157045
rect 104433 157040 198891 157042
rect 104433 156984 104438 157040
rect 104494 156984 198830 157040
rect 198886 156984 198891 157040
rect 104433 156982 198891 156984
rect 104433 156979 104499 156982
rect 198825 156979 198891 156982
rect 101949 156906 102015 156909
rect 196801 156906 196867 156909
rect 101949 156904 196867 156906
rect 101949 156848 101954 156904
rect 102010 156848 196806 156904
rect 196862 156848 196867 156904
rect 101949 156846 196867 156848
rect 101949 156843 102015 156846
rect 196801 156843 196867 156846
rect 91829 156770 91895 156773
rect 189165 156770 189231 156773
rect 91829 156768 189231 156770
rect 91829 156712 91834 156768
rect 91890 156712 189170 156768
rect 189226 156712 189231 156768
rect 91829 156710 189231 156712
rect 91829 156707 91895 156710
rect 189165 156707 189231 156710
rect 33961 156634 34027 156637
rect 145189 156634 145255 156637
rect 33961 156632 145255 156634
rect 33961 156576 33966 156632
rect 34022 156576 145194 156632
rect 145250 156576 145255 156632
rect 33961 156574 145255 156576
rect 33961 156571 34027 156574
rect 145189 156571 145255 156574
rect 519629 156226 519695 156229
rect 523200 156226 524400 156256
rect 519629 156224 524400 156226
rect 519629 156168 519634 156224
rect 519690 156168 524400 156224
rect 519629 156166 524400 156168
rect 519629 156163 519695 156166
rect 523200 156136 524400 156166
rect 8293 156090 8359 156093
rect 124949 156090 125015 156093
rect 8293 156088 125015 156090
rect 8293 156032 8298 156088
rect 8354 156032 124954 156088
rect 125010 156032 125015 156088
rect 8293 156030 125015 156032
rect 8293 156027 8359 156030
rect 124949 156027 125015 156030
rect 28901 155954 28967 155957
rect 131113 155954 131179 155957
rect 28901 155952 131179 155954
rect 28901 155896 28906 155952
rect 28962 155896 131118 155952
rect 131174 155896 131179 155952
rect 28901 155894 131179 155896
rect 28901 155891 28967 155894
rect 131113 155891 131179 155894
rect 29729 155818 29795 155821
rect 138013 155818 138079 155821
rect 29729 155816 138079 155818
rect 29729 155760 29734 155816
rect 29790 155760 138018 155816
rect 138074 155760 138079 155816
rect 29729 155758 138079 155760
rect 29729 155755 29795 155758
rect 138013 155755 138079 155758
rect 173433 155818 173499 155821
rect 175825 155818 175891 155821
rect 173433 155816 175891 155818
rect 173433 155760 173438 155816
rect 173494 155760 175830 155816
rect 175886 155760 175891 155816
rect 173433 155758 175891 155760
rect 173433 155755 173499 155758
rect 175825 155755 175891 155758
rect 23013 155682 23079 155685
rect 134517 155682 134583 155685
rect 23013 155680 134583 155682
rect 23013 155624 23018 155680
rect 23074 155624 134522 155680
rect 134578 155624 134583 155680
rect 23013 155622 134583 155624
rect 23013 155619 23079 155622
rect 134517 155619 134583 155622
rect 207749 155682 207815 155685
rect 273345 155682 273411 155685
rect 207749 155680 273411 155682
rect 207749 155624 207754 155680
rect 207810 155624 273350 155680
rect 273406 155624 273411 155680
rect 207749 155622 273411 155624
rect 207749 155619 207815 155622
rect 273345 155619 273411 155622
rect 274909 155682 274975 155685
rect 329189 155682 329255 155685
rect 274909 155680 329255 155682
rect 274909 155624 274914 155680
rect 274970 155624 329194 155680
rect 329250 155624 329255 155680
rect 274909 155622 329255 155624
rect 274909 155619 274975 155622
rect 329189 155619 329255 155622
rect 16297 155546 16363 155549
rect 131021 155546 131087 155549
rect 16297 155544 131087 155546
rect 16297 155488 16302 155544
rect 16358 155488 131026 155544
rect 131082 155488 131087 155544
rect 16297 155486 131087 155488
rect 16297 155483 16363 155486
rect 131021 155483 131087 155486
rect 147305 155546 147371 155549
rect 222561 155546 222627 155549
rect 147305 155544 222627 155546
rect 147305 155488 147310 155544
rect 147366 155488 222566 155544
rect 222622 155488 222627 155544
rect 147305 155486 222627 155488
rect 147305 155483 147371 155486
rect 222561 155483 222627 155486
rect 222745 155546 222811 155549
rect 223573 155546 223639 155549
rect 222745 155544 223639 155546
rect 222745 155488 222750 155544
rect 222806 155488 223578 155544
rect 223634 155488 223639 155544
rect 222745 155486 223639 155488
rect 222745 155483 222811 155486
rect 223573 155483 223639 155486
rect 240409 155546 240475 155549
rect 242985 155546 243051 155549
rect 240409 155544 243051 155546
rect 240409 155488 240414 155544
rect 240470 155488 242990 155544
rect 243046 155488 243051 155544
rect 240409 155486 243051 155488
rect 240409 155483 240475 155486
rect 242985 155483 243051 155486
rect 254761 155546 254827 155549
rect 310605 155546 310671 155549
rect 254761 155544 310671 155546
rect 254761 155488 254766 155544
rect 254822 155488 310610 155544
rect 310666 155488 310671 155544
rect 254761 155486 310671 155488
rect 254761 155483 254827 155486
rect 310605 155483 310671 155486
rect 311893 155546 311959 155549
rect 316769 155546 316835 155549
rect 311893 155544 316835 155546
rect 311893 155488 311898 155544
rect 311954 155488 316774 155544
rect 316830 155488 316835 155544
rect 311893 155486 316835 155488
rect 311893 155483 311959 155486
rect 316769 155483 316835 155486
rect 107745 155410 107811 155413
rect 109033 155410 109099 155413
rect 107745 155408 109099 155410
rect 107745 155352 107750 155408
rect 107806 155352 109038 155408
rect 109094 155352 109099 155408
rect 107745 155350 109099 155352
rect 107745 155347 107811 155350
rect 109033 155347 109099 155350
rect 120441 155410 120507 155413
rect 208669 155410 208735 155413
rect 120441 155408 208735 155410
rect 120441 155352 120446 155408
rect 120502 155352 208674 155408
rect 208730 155352 208735 155408
rect 120441 155350 208735 155352
rect 120441 155347 120507 155350
rect 208669 155347 208735 155350
rect 214465 155410 214531 155413
rect 279509 155410 279575 155413
rect 214465 155408 279575 155410
rect 214465 155352 214470 155408
rect 214526 155352 279514 155408
rect 279570 155352 279575 155408
rect 214465 155350 279575 155352
rect 214465 155347 214531 155350
rect 279509 155347 279575 155350
rect 299565 155410 299631 155413
rect 309133 155410 309199 155413
rect 299565 155408 309199 155410
rect 299565 155352 299570 155408
rect 299626 155352 309138 155408
rect 309194 155352 309199 155408
rect 299565 155350 309199 155352
rect 299565 155347 299631 155350
rect 309133 155347 309199 155350
rect 311709 155410 311775 155413
rect 312077 155410 312143 155413
rect 311709 155408 312143 155410
rect 311709 155352 311714 155408
rect 311770 155352 312082 155408
rect 312138 155352 312143 155408
rect 311709 155350 312143 155352
rect 311709 155347 311775 155350
rect 312077 155347 312143 155350
rect 9581 155274 9647 155277
rect 126237 155274 126303 155277
rect 9581 155272 126303 155274
rect 9581 155216 9586 155272
rect 9642 155216 126242 155272
rect 126298 155216 126303 155272
rect 9581 155214 126303 155216
rect 9581 155211 9647 155214
rect 126237 155211 126303 155214
rect 132953 155274 133019 155277
rect 137369 155274 137435 155277
rect 132953 155272 137435 155274
rect 132953 155216 132958 155272
rect 133014 155216 137374 155272
rect 137430 155216 137435 155272
rect 132953 155214 137435 155216
rect 132953 155211 133019 155214
rect 137369 155211 137435 155214
rect 140589 155274 140655 155277
rect 223573 155274 223639 155277
rect 140589 155272 223639 155274
rect 140589 155216 140594 155272
rect 140650 155216 223578 155272
rect 223634 155216 223639 155272
rect 140589 155214 223639 155216
rect 140589 155211 140655 155214
rect 223573 155211 223639 155214
rect 227897 155274 227963 155277
rect 293217 155274 293283 155277
rect 227897 155272 293283 155274
rect 227897 155216 227902 155272
rect 227958 155216 293222 155272
rect 293278 155216 293283 155272
rect 227897 155214 293283 155216
rect 227897 155211 227963 155214
rect 293217 155211 293283 155214
rect 295149 155274 295215 155277
rect 342161 155274 342227 155277
rect 295149 155272 342227 155274
rect 295149 155216 295154 155272
rect 295210 155216 342166 155272
rect 342222 155216 342227 155272
rect 295149 155214 342227 155216
rect 295149 155211 295215 155214
rect 342161 155211 342227 155214
rect 349889 155274 349955 155277
rect 354581 155274 354647 155277
rect 349889 155272 354647 155274
rect 349889 155216 349894 155272
rect 349950 155216 354586 155272
rect 354642 155216 354647 155272
rect 349889 155214 354647 155216
rect 349889 155211 349955 155214
rect 354581 155211 354647 155214
rect 2865 155138 2931 155141
rect 121085 155138 121151 155141
rect 2865 155136 121151 155138
rect 2865 155080 2870 155136
rect 2926 155080 121090 155136
rect 121146 155080 121151 155136
rect 2865 155078 121151 155080
rect 2865 155075 2931 155078
rect 121085 155075 121151 155078
rect 222561 155138 222627 155141
rect 227805 155138 227871 155141
rect 222561 155136 227871 155138
rect 222561 155080 222566 155136
rect 222622 155080 227810 155136
rect 227866 155080 227871 155136
rect 222561 155078 227871 155080
rect 222561 155075 222627 155078
rect 227805 155075 227871 155078
rect 260557 155138 260623 155141
rect 263685 155138 263751 155141
rect 260557 155136 263751 155138
rect 260557 155080 260562 155136
rect 260618 155080 263690 155136
rect 263746 155080 263751 155136
rect 260557 155078 263751 155080
rect 260557 155075 260623 155078
rect 263685 155075 263751 155078
rect 348785 155138 348851 155141
rect 354213 155138 354279 155141
rect 348785 155136 354279 155138
rect 348785 155080 348790 155136
rect 348846 155080 354218 155136
rect 354274 155080 354279 155136
rect 348785 155078 354279 155080
rect 348785 155075 348851 155078
rect 354213 155075 354279 155078
rect 211889 155002 211955 155005
rect 212533 155002 212599 155005
rect 211889 155000 212599 155002
rect 211889 154944 211894 155000
rect 211950 154944 212538 155000
rect 212594 154944 212599 155000
rect 211889 154942 212599 154944
rect 211889 154939 211955 154942
rect 212533 154939 212599 154942
rect 232037 155002 232103 155005
rect 233233 155002 233299 155005
rect 232037 155000 233299 155002
rect 232037 154944 232042 155000
rect 232098 154944 233238 155000
rect 233294 154944 233299 155000
rect 232037 154942 233299 154944
rect 232037 154939 232103 154942
rect 233233 154939 233299 154942
rect 279877 155002 279943 155005
rect 282913 155002 282979 155005
rect 279877 155000 282979 155002
rect 279877 154944 279882 155000
rect 279938 154944 282918 155000
rect 282974 154944 282979 155000
rect 279877 154942 282979 154944
rect 279877 154939 279943 154942
rect 282913 154939 282979 154942
rect 292389 155002 292455 155005
rect 293953 155002 294019 155005
rect 292389 155000 294019 155002
rect 292389 154944 292394 155000
rect 292450 154944 293958 155000
rect 294014 154944 294019 155000
rect 292389 154942 294019 154944
rect 292389 154939 292455 154942
rect 293953 154939 294019 154942
rect 311433 155002 311499 155005
rect 311801 155002 311867 155005
rect 311433 155000 311867 155002
rect 311433 154944 311438 155000
rect 311494 154944 311806 155000
rect 311862 154944 311867 155000
rect 311433 154942 311867 154944
rect 311433 154939 311499 154942
rect 311801 154939 311867 154942
rect 321829 155002 321895 155005
rect 322197 155002 322263 155005
rect 321829 155000 322263 155002
rect 321829 154944 321834 155000
rect 321890 154944 322202 155000
rect 322258 154944 322263 155000
rect 321829 154942 322263 154944
rect 321829 154939 321895 154942
rect 322197 154939 322263 154942
rect 340505 155002 340571 155005
rect 341241 155002 341307 155005
rect 340505 155000 341307 155002
rect 340505 154944 340510 155000
rect 340566 154944 341246 155000
rect 341302 154944 341307 155000
rect 340505 154942 341307 154944
rect 340505 154939 340571 154942
rect 341241 154939 341307 154942
rect 113173 154866 113239 154869
rect 115933 154866 115999 154869
rect 113173 154864 115999 154866
rect 113173 154808 113178 154864
rect 113234 154808 115938 154864
rect 115994 154808 115999 154864
rect 113173 154806 115999 154808
rect 113173 154803 113239 154806
rect 115933 154803 115999 154806
rect 136909 154866 136975 154869
rect 137553 154866 137619 154869
rect 136909 154864 137619 154866
rect 136909 154808 136914 154864
rect 136970 154808 137558 154864
rect 137614 154808 137619 154864
rect 136909 154806 137619 154808
rect 136909 154803 136975 154806
rect 137553 154803 137619 154806
rect 238569 154866 238635 154869
rect 239029 154866 239095 154869
rect 238569 154864 239095 154866
rect 238569 154808 238574 154864
rect 238630 154808 239034 154864
rect 239090 154808 239095 154864
rect 238569 154806 239095 154808
rect 238569 154803 238635 154806
rect 239029 154803 239095 154806
rect 299657 154866 299723 154869
rect 303521 154866 303587 154869
rect 299657 154864 303587 154866
rect 299657 154808 299662 154864
rect 299718 154808 303526 154864
rect 303582 154808 303587 154864
rect 299657 154806 303587 154808
rect 299657 154803 299723 154806
rect 303521 154803 303587 154806
rect 340229 154866 340295 154869
rect 340873 154866 340939 154869
rect 340229 154864 340939 154866
rect 340229 154808 340234 154864
rect 340290 154808 340878 154864
rect 340934 154808 340939 154864
rect 340229 154806 340939 154808
rect 340229 154803 340295 154806
rect 340873 154803 340939 154806
rect 112897 154730 112963 154733
rect 113449 154730 113515 154733
rect 112897 154728 113515 154730
rect 112897 154672 112902 154728
rect 112958 154672 113454 154728
rect 113510 154672 113515 154728
rect 112897 154670 113515 154672
rect 112897 154667 112963 154670
rect 113449 154667 113515 154670
rect 113633 154730 113699 154733
rect 116853 154730 116919 154733
rect 113633 154728 116919 154730
rect 113633 154672 113638 154728
rect 113694 154672 116858 154728
rect 116914 154672 116919 154728
rect 113633 154670 116919 154672
rect 113633 154667 113699 154670
rect 116853 154667 116919 154670
rect 190821 154730 190887 154733
rect 192017 154730 192083 154733
rect 190821 154728 192083 154730
rect 190821 154672 190826 154728
rect 190882 154672 192022 154728
rect 192078 154672 192083 154728
rect 190821 154670 192083 154672
rect 190821 154667 190887 154670
rect 192017 154667 192083 154670
rect 340321 154730 340387 154733
rect 342805 154730 342871 154733
rect 340321 154728 342871 154730
rect 340321 154672 340326 154728
rect 340382 154672 342810 154728
rect 342866 154672 342871 154728
rect 340321 154670 342871 154672
rect 340321 154667 340387 154670
rect 342805 154667 342871 154670
rect 519721 154730 519787 154733
rect 523200 154730 524400 154760
rect 519721 154728 524400 154730
rect 519721 154672 519726 154728
rect 519782 154672 524400 154728
rect 519721 154670 524400 154672
rect 519721 154667 519787 154670
rect 523200 154640 524400 154670
rect 326061 154594 326127 154597
rect 327625 154594 327691 154597
rect 326061 154592 327691 154594
rect 326061 154536 326066 154592
rect 326122 154536 327630 154592
rect 327686 154536 327691 154592
rect 326061 154534 327691 154536
rect 326061 154531 326127 154534
rect 327625 154531 327691 154534
rect 108665 154458 108731 154461
rect 202045 154458 202111 154461
rect 108665 154456 202111 154458
rect 108665 154400 108670 154456
rect 108726 154400 202050 154456
rect 202106 154400 202111 154456
rect 108665 154398 202111 154400
rect 108665 154395 108731 154398
rect 202045 154395 202111 154398
rect 262397 154458 262463 154461
rect 319529 154458 319595 154461
rect 262397 154456 319595 154458
rect 262397 154400 262402 154456
rect 262458 154400 319534 154456
rect 319590 154400 319595 154456
rect 262397 154398 319595 154400
rect 262397 154395 262463 154398
rect 319529 154395 319595 154398
rect 98637 154322 98703 154325
rect 193213 154322 193279 154325
rect 218053 154322 218119 154325
rect 98637 154320 186330 154322
rect 98637 154264 98642 154320
rect 98698 154264 186330 154320
rect 98637 154262 186330 154264
rect 98637 154259 98703 154262
rect 61653 154186 61719 154189
rect 166073 154186 166139 154189
rect 61653 154184 166139 154186
rect 61653 154128 61658 154184
rect 61714 154128 166078 154184
rect 166134 154128 166139 154184
rect 61653 154126 166139 154128
rect 186270 154186 186330 154262
rect 193213 154320 218119 154322
rect 193213 154264 193218 154320
rect 193274 154264 218058 154320
rect 218114 154264 218119 154320
rect 193213 154262 218119 154264
rect 193213 154259 193279 154262
rect 218053 154259 218119 154262
rect 220721 154322 220787 154325
rect 233509 154322 233575 154325
rect 220721 154320 233575 154322
rect 220721 154264 220726 154320
rect 220782 154264 233514 154320
rect 233570 154264 233575 154320
rect 220721 154262 233575 154264
rect 220721 154259 220787 154262
rect 233509 154259 233575 154262
rect 265709 154322 265775 154325
rect 322105 154322 322171 154325
rect 265709 154320 322171 154322
rect 265709 154264 265714 154320
rect 265770 154264 322110 154320
rect 322166 154264 322171 154320
rect 265709 154262 322171 154264
rect 265709 154259 265775 154262
rect 322105 154259 322171 154262
rect 331213 154322 331279 154325
rect 336181 154322 336247 154325
rect 331213 154320 336247 154322
rect 331213 154264 331218 154320
rect 331274 154264 336186 154320
rect 336242 154264 336247 154320
rect 331213 154262 336247 154264
rect 331213 154259 331279 154262
rect 336181 154259 336247 154262
rect 342713 154322 342779 154325
rect 345749 154322 345815 154325
rect 342713 154320 345815 154322
rect 342713 154264 342718 154320
rect 342774 154264 345754 154320
rect 345810 154264 345815 154320
rect 342713 154262 345815 154264
rect 342713 154259 342779 154262
rect 345749 154259 345815 154262
rect 194317 154186 194383 154189
rect 186270 154184 194383 154186
rect 186270 154128 194322 154184
rect 194378 154128 194383 154184
rect 186270 154126 194383 154128
rect 61653 154123 61719 154126
rect 166073 154123 166139 154126
rect 194317 154123 194383 154126
rect 206093 154186 206159 154189
rect 276473 154186 276539 154189
rect 206093 154184 276539 154186
rect 206093 154128 206098 154184
rect 206154 154128 276478 154184
rect 276534 154128 276539 154184
rect 206093 154126 276539 154128
rect 206093 154123 206159 154126
rect 276473 154123 276539 154126
rect 292297 154186 292363 154189
rect 292665 154186 292731 154189
rect 292297 154184 292731 154186
rect 292297 154128 292302 154184
rect 292358 154128 292670 154184
rect 292726 154128 292731 154184
rect 292297 154126 292731 154128
rect 292297 154123 292363 154126
rect 292665 154123 292731 154126
rect 292849 154186 292915 154189
rect 299657 154186 299723 154189
rect 292849 154184 299723 154186
rect 292849 154128 292854 154184
rect 292910 154128 299662 154184
rect 299718 154128 299723 154184
rect 292849 154126 299723 154128
rect 292849 154123 292915 154126
rect 299657 154123 299723 154126
rect 44817 154050 44883 154053
rect 153193 154050 153259 154053
rect 44817 154048 153259 154050
rect 44817 153992 44822 154048
rect 44878 153992 153198 154048
rect 153254 153992 153259 154048
rect 44817 153990 153259 153992
rect 44817 153987 44883 153990
rect 153193 153987 153259 153990
rect 205265 154050 205331 154053
rect 275737 154050 275803 154053
rect 205265 154048 275803 154050
rect 205265 153992 205270 154048
rect 205326 153992 275742 154048
rect 275798 153992 275803 154048
rect 205265 153990 275803 153992
rect 205265 153987 205331 153990
rect 275737 153987 275803 153990
rect 278681 154050 278747 154053
rect 312261 154050 312327 154053
rect 278681 154048 312327 154050
rect 278681 153992 278686 154048
rect 278742 153992 312266 154048
rect 312322 153992 312327 154048
rect 278681 153990 312327 153992
rect 278681 153987 278747 153990
rect 312261 153987 312327 153990
rect 20529 153914 20595 153917
rect 134609 153914 134675 153917
rect 20529 153912 134675 153914
rect 20529 153856 20534 153912
rect 20590 153856 134614 153912
rect 134670 153856 134675 153912
rect 20529 153854 134675 153856
rect 20529 153851 20595 153854
rect 134609 153851 134675 153854
rect 164233 153914 164299 153917
rect 200113 153914 200179 153917
rect 164233 153912 200179 153914
rect 164233 153856 164238 153912
rect 164294 153856 200118 153912
rect 200174 153856 200179 153912
rect 164233 153854 200179 153856
rect 164233 153851 164299 153854
rect 200113 153851 200179 153854
rect 201861 153914 201927 153917
rect 273253 153914 273319 153917
rect 201861 153912 273319 153914
rect 201861 153856 201866 153912
rect 201922 153856 273258 153912
rect 273314 153856 273319 153912
rect 201861 153854 273319 153856
rect 201861 153851 201927 153854
rect 273253 153851 273319 153854
rect 275829 153914 275895 153917
rect 329833 153914 329899 153917
rect 275829 153912 329899 153914
rect 275829 153856 275834 153912
rect 275890 153856 329838 153912
rect 329894 153856 329899 153912
rect 275829 153854 329899 153856
rect 275829 153851 275895 153854
rect 329833 153851 329899 153854
rect 2037 153778 2103 153781
rect 120441 153778 120507 153781
rect 2037 153776 120507 153778
rect 2037 153720 2042 153776
rect 2098 153720 120446 153776
rect 120502 153720 120507 153776
rect 2037 153718 120507 153720
rect 2037 153715 2103 153718
rect 120441 153715 120507 153718
rect 138933 153778 138999 153781
rect 225137 153778 225203 153781
rect 138933 153776 225203 153778
rect 138933 153720 138938 153776
rect 138994 153720 225142 153776
rect 225198 153720 225203 153776
rect 138933 153718 225203 153720
rect 138933 153715 138999 153718
rect 225137 153715 225203 153718
rect 229645 153778 229711 153781
rect 294505 153778 294571 153781
rect 229645 153776 294571 153778
rect 229645 153720 229650 153776
rect 229706 153720 294510 153776
rect 294566 153720 294571 153776
rect 229645 153718 294571 153720
rect 229645 153715 229711 153718
rect 294505 153715 294571 153718
rect 320173 153778 320239 153781
rect 338113 153778 338179 153781
rect 320173 153776 338179 153778
rect 320173 153720 320178 153776
rect 320234 153720 338118 153776
rect 338174 153720 338179 153776
rect 320173 153718 338179 153720
rect 320173 153715 320239 153718
rect 338113 153715 338179 153718
rect 118785 153642 118851 153645
rect 209773 153642 209839 153645
rect 118785 153640 209839 153642
rect 118785 153584 118790 153640
rect 118846 153584 209778 153640
rect 209834 153584 209839 153640
rect 118785 153582 209839 153584
rect 118785 153579 118851 153582
rect 209773 153579 209839 153582
rect 312353 153642 312419 153645
rect 312905 153642 312971 153645
rect 312353 153640 312971 153642
rect 312353 153584 312358 153640
rect 312414 153584 312910 153640
rect 312966 153584 312971 153640
rect 312353 153582 312971 153584
rect 312353 153579 312419 153582
rect 312905 153579 312971 153582
rect 325233 153506 325299 153509
rect 327533 153506 327599 153509
rect 325233 153504 327599 153506
rect 325233 153448 325238 153504
rect 325294 153448 327538 153504
rect 327594 153448 327599 153504
rect 325233 153446 327599 153448
rect 325233 153443 325299 153446
rect 327533 153443 327599 153446
rect 311709 153370 311775 153373
rect 311893 153370 311959 153373
rect 311709 153368 311959 153370
rect 311709 153312 311714 153368
rect 311770 153312 311898 153368
rect 311954 153312 311959 153368
rect 311709 153310 311959 153312
rect 311709 153307 311775 153310
rect 311893 153307 311959 153310
rect 337009 153370 337075 153373
rect 339401 153370 339467 153373
rect 337009 153368 339467 153370
rect 337009 153312 337014 153368
rect 337070 153312 339406 153368
rect 339462 153312 339467 153368
rect 337009 153310 339467 153312
rect 337009 153307 337075 153310
rect 339401 153307 339467 153310
rect 342897 153370 342963 153373
rect 345381 153370 345447 153373
rect 342897 153368 345447 153370
rect 342897 153312 342902 153368
rect 342958 153312 345386 153368
rect 345442 153312 345447 153368
rect 342897 153310 345447 153312
rect 342897 153307 342963 153310
rect 345381 153307 345447 153310
rect 286869 153234 286935 153237
rect 291469 153234 291535 153237
rect 286869 153232 291535 153234
rect 286869 153176 286874 153232
rect 286930 153176 291474 153232
rect 291530 153176 291535 153232
rect 286869 153174 291535 153176
rect 286869 153171 286935 153174
rect 291469 153171 291535 153174
rect 316217 153234 316283 153237
rect 317137 153234 317203 153237
rect 316217 153232 317203 153234
rect 316217 153176 316222 153232
rect 316278 153176 317142 153232
rect 317198 153176 317203 153232
rect 316217 153174 317203 153176
rect 316217 153171 316283 153174
rect 317137 153171 317203 153174
rect 328637 153234 328703 153237
rect 332777 153234 332843 153237
rect 328637 153232 332843 153234
rect 328637 153176 328642 153232
rect 328698 153176 332782 153232
rect 332838 153176 332843 153232
rect 328637 153174 332843 153176
rect 328637 153171 328703 153174
rect 332777 153171 332843 153174
rect 519813 153234 519879 153237
rect 523200 153234 524400 153264
rect 519813 153232 524400 153234
rect 519813 153176 519818 153232
rect 519874 153176 524400 153232
rect 519813 153174 524400 153176
rect 519813 153171 519879 153174
rect 523200 153144 524400 153174
rect 91093 153098 91159 153101
rect 130745 153098 130811 153101
rect 91093 153096 130811 153098
rect 91093 153040 91098 153096
rect 91154 153040 130750 153096
rect 130806 153040 130811 153096
rect 91093 153038 130811 153040
rect 91093 153035 91159 153038
rect 130745 153035 130811 153038
rect 131113 153098 131179 153101
rect 141049 153098 141115 153101
rect 131113 153096 141115 153098
rect 131113 153040 131118 153096
rect 131174 153040 141054 153096
rect 141110 153040 141115 153096
rect 131113 153038 141115 153040
rect 131113 153035 131179 153038
rect 141049 153035 141115 153038
rect 270217 153098 270283 153101
rect 272701 153098 272767 153101
rect 270217 153096 272767 153098
rect 270217 153040 270222 153096
rect 270278 153040 272706 153096
rect 272762 153040 272767 153096
rect 270217 153038 272767 153040
rect 270217 153035 270283 153038
rect 272701 153035 272767 153038
rect 320265 153098 320331 153101
rect 323393 153098 323459 153101
rect 320265 153096 323459 153098
rect 320265 153040 320270 153096
rect 320326 153040 323398 153096
rect 323454 153040 323459 153096
rect 320265 153038 323459 153040
rect 320265 153035 320331 153038
rect 323393 153035 323459 153038
rect 109125 152962 109191 152965
rect 162853 152962 162919 152965
rect 109125 152960 162919 152962
rect 109125 152904 109130 152960
rect 109186 152904 162858 152960
rect 162914 152904 162919 152960
rect 109125 152902 162919 152904
rect 109125 152899 109191 152902
rect 162853 152899 162919 152902
rect 93577 152826 93643 152829
rect 190453 152826 190519 152829
rect 93577 152824 190519 152826
rect 93577 152768 93582 152824
rect 93638 152768 190458 152824
rect 190514 152768 190519 152824
rect 93577 152766 190519 152768
rect 93577 152763 93643 152766
rect 190453 152763 190519 152766
rect 200205 152826 200271 152829
rect 269481 152826 269547 152829
rect 200205 152824 269547 152826
rect 200205 152768 200210 152824
rect 200266 152768 269486 152824
rect 269542 152768 269547 152824
rect 200205 152766 269547 152768
rect 200205 152763 200271 152766
rect 269481 152763 269547 152766
rect 278313 152826 278379 152829
rect 331765 152826 331831 152829
rect 278313 152824 331831 152826
rect 278313 152768 278318 152824
rect 278374 152768 331770 152824
rect 331826 152768 331831 152824
rect 278313 152766 331831 152768
rect 278313 152763 278379 152766
rect 331765 152763 331831 152766
rect 19609 152690 19675 152693
rect 133965 152690 134031 152693
rect 19609 152688 134031 152690
rect 19609 152632 19614 152688
rect 19670 152632 133970 152688
rect 134026 152632 134031 152688
rect 19609 152630 134031 152632
rect 19609 152627 19675 152630
rect 133965 152627 134031 152630
rect 134517 152690 134583 152693
rect 136541 152690 136607 152693
rect 134517 152688 136607 152690
rect 134517 152632 134522 152688
rect 134578 152632 136546 152688
rect 136602 152632 136607 152688
rect 134517 152630 136607 152632
rect 134517 152627 134583 152630
rect 136541 152627 136607 152630
rect 191833 152690 191899 152693
rect 264973 152690 265039 152693
rect 191833 152688 265039 152690
rect 191833 152632 191838 152688
rect 191894 152632 264978 152688
rect 265034 152632 265039 152688
rect 191833 152630 265039 152632
rect 191833 152627 191899 152630
rect 264973 152627 265039 152630
rect 266445 152690 266511 152693
rect 321461 152690 321527 152693
rect 266445 152688 321527 152690
rect 266445 152632 266450 152688
rect 266506 152632 321466 152688
rect 321522 152632 321527 152688
rect 266445 152630 321527 152632
rect 266445 152627 266511 152630
rect 321461 152627 321527 152630
rect 18781 152554 18847 152557
rect 133229 152554 133295 152557
rect 218697 152554 218763 152557
rect 18781 152552 132510 152554
rect 18781 152496 18786 152552
rect 18842 152496 132510 152552
rect 18781 152494 132510 152496
rect 18781 152491 18847 152494
rect 6177 152418 6243 152421
rect 123661 152418 123727 152421
rect 6177 152416 123727 152418
rect 6177 152360 6182 152416
rect 6238 152360 123666 152416
rect 123722 152360 123727 152416
rect 6177 152358 123727 152360
rect 132450 152418 132510 152494
rect 133229 152552 218763 152554
rect 133229 152496 133234 152552
rect 133290 152496 218702 152552
rect 218758 152496 218763 152552
rect 133229 152494 218763 152496
rect 133229 152491 133295 152494
rect 218697 152491 218763 152494
rect 220813 152554 220879 152557
rect 287421 152554 287487 152557
rect 220813 152552 287487 152554
rect 220813 152496 220818 152552
rect 220874 152496 287426 152552
rect 287482 152496 287487 152552
rect 220813 152494 287487 152496
rect 220813 152491 220879 152494
rect 287421 152491 287487 152494
rect 133321 152418 133387 152421
rect 215477 152418 215543 152421
rect 132450 152416 133387 152418
rect 132450 152360 133326 152416
rect 133382 152360 133387 152416
rect 132450 152358 133387 152360
rect 6177 152355 6243 152358
rect 123661 152355 123727 152358
rect 133321 152355 133387 152358
rect 142110 152416 215543 152418
rect 142110 152360 215482 152416
rect 215538 152360 215543 152416
rect 142110 152358 215543 152360
rect 109033 152282 109099 152285
rect 125593 152282 125659 152285
rect 109033 152280 125659 152282
rect 109033 152224 109038 152280
rect 109094 152224 125598 152280
rect 125654 152224 125659 152280
rect 109033 152222 125659 152224
rect 109033 152219 109099 152222
rect 125593 152219 125659 152222
rect 126329 152282 126395 152285
rect 142110 152282 142170 152358
rect 215477 152355 215543 152358
rect 217869 152418 217935 152421
rect 285489 152418 285555 152421
rect 217869 152416 285555 152418
rect 217869 152360 217874 152416
rect 217930 152360 285494 152416
rect 285550 152360 285555 152416
rect 217869 152358 285555 152360
rect 217869 152355 217935 152358
rect 285489 152355 285555 152358
rect 287053 152418 287119 152421
rect 336825 152418 336891 152421
rect 287053 152416 336891 152418
rect 287053 152360 287058 152416
rect 287114 152360 336830 152416
rect 336886 152360 336891 152416
rect 287053 152358 336891 152360
rect 287053 152355 287119 152358
rect 336825 152355 336891 152358
rect 432873 152418 432939 152421
rect 449893 152418 449959 152421
rect 432873 152416 449959 152418
rect 432873 152360 432878 152416
rect 432934 152360 449898 152416
rect 449954 152360 449959 152416
rect 432873 152358 449959 152360
rect 432873 152355 432939 152358
rect 449893 152355 449959 152358
rect 126329 152280 142170 152282
rect 126329 152224 126334 152280
rect 126390 152224 142170 152280
rect 126329 152222 142170 152224
rect 126329 152219 126395 152222
rect 36997 152146 37063 152149
rect 109861 152146 109927 152149
rect 36997 152144 109927 152146
rect 36997 152088 37002 152144
rect 37058 152088 109866 152144
rect 109922 152088 109927 152144
rect 36997 152086 109927 152088
rect 36997 152083 37063 152086
rect 109861 152083 109927 152086
rect 16389 152010 16455 152013
rect 116209 152010 116275 152013
rect 16389 152008 116275 152010
rect 16389 151952 16394 152008
rect 16450 151952 116214 152008
rect 116270 151952 116275 152008
rect 16389 151950 116275 151952
rect 16389 151947 16455 151950
rect 116209 151947 116275 151950
rect 2681 151874 2747 151877
rect 109677 151874 109743 151877
rect 2681 151872 109743 151874
rect 2681 151816 2686 151872
rect 2742 151816 109682 151872
rect 109738 151816 109743 151872
rect 2681 151814 109743 151816
rect 2681 151811 2747 151814
rect 109677 151811 109743 151814
rect 273345 151874 273411 151877
rect 277761 151874 277827 151877
rect 273345 151872 277827 151874
rect 273345 151816 273350 151872
rect 273406 151816 277766 151872
rect 277822 151816 277827 151872
rect 273345 151814 277827 151816
rect 273345 151811 273411 151814
rect 277761 151811 277827 151814
rect 521009 151738 521075 151741
rect 523200 151738 524400 151768
rect 521009 151736 524400 151738
rect 521009 151680 521014 151736
rect 521070 151680 524400 151736
rect 521009 151678 524400 151680
rect 521009 151675 521075 151678
rect 523200 151648 524400 151678
rect 33593 151602 33659 151605
rect 112437 151602 112503 151605
rect 33593 151600 112503 151602
rect 33593 151544 33598 151600
rect 33654 151544 112442 151600
rect 112498 151544 112503 151600
rect 33593 151542 112503 151544
rect 33593 151539 33659 151542
rect 112437 151539 112503 151542
rect 9489 151466 9555 151469
rect 110873 151466 110939 151469
rect 9489 151464 110939 151466
rect 9489 151408 9494 151464
rect 9550 151408 110878 151464
rect 110934 151408 110939 151464
rect 9489 151406 110939 151408
rect 9489 151403 9555 151406
rect 110873 151403 110939 151406
rect 116577 151466 116643 151469
rect 184657 151466 184723 151469
rect 116577 151464 184723 151466
rect 116577 151408 116582 151464
rect 116638 151408 184662 151464
rect 184718 151408 184723 151464
rect 116577 151406 184723 151408
rect 116577 151403 116643 151406
rect 184657 151403 184723 151406
rect 111701 151330 111767 151333
rect 203977 151330 204043 151333
rect 111701 151328 204043 151330
rect 111701 151272 111706 151328
rect 111762 151272 203982 151328
rect 204038 151272 204043 151328
rect 111701 151270 204043 151272
rect 111701 151267 111767 151270
rect 203977 151267 204043 151270
rect 30189 151194 30255 151197
rect 111701 151194 111767 151197
rect 30189 151192 111767 151194
rect 30189 151136 30194 151192
rect 30250 151136 111706 151192
rect 111762 151136 111767 151192
rect 30189 151134 111767 151136
rect 30189 151131 30255 151134
rect 111701 151131 111767 151134
rect 115841 151194 115907 151197
rect 207197 151194 207263 151197
rect 115841 151192 207263 151194
rect 115841 151136 115846 151192
rect 115902 151136 207202 151192
rect 207258 151136 207263 151192
rect 115841 151134 207263 151136
rect 115841 151131 115907 151134
rect 207197 151131 207263 151134
rect 67541 151058 67607 151061
rect 170581 151058 170647 151061
rect 67541 151056 170647 151058
rect 67541 151000 67546 151056
rect 67602 151000 170586 151056
rect 170642 151000 170647 151056
rect 67541 150998 170647 151000
rect 67541 150995 67607 150998
rect 170581 150995 170647 150998
rect 23289 150922 23355 150925
rect 110965 150922 111031 150925
rect 23289 150920 111031 150922
rect 23289 150864 23294 150920
rect 23350 150864 110970 150920
rect 111026 150864 111031 150920
rect 23289 150862 111031 150864
rect 23289 150859 23355 150862
rect 110965 150859 111031 150862
rect 19793 150786 19859 150789
rect 109769 150786 109835 150789
rect 19793 150784 109835 150786
rect 19793 150728 19798 150784
rect 19854 150728 109774 150784
rect 109830 150728 109835 150784
rect 19793 150726 109835 150728
rect 19793 150723 19859 150726
rect 109769 150723 109835 150726
rect 12985 150650 13051 150653
rect 111333 150650 111399 150653
rect 12985 150648 111399 150650
rect 12985 150592 12990 150648
rect 13046 150592 111338 150648
rect 111394 150592 111399 150648
rect 12985 150590 111399 150592
rect 12985 150587 13051 150590
rect 111333 150587 111399 150590
rect 109217 150514 109283 150517
rect 111149 150514 111215 150517
rect 109217 150512 111215 150514
rect 109217 150456 109222 150512
rect 109278 150456 111154 150512
rect 111210 150456 111215 150512
rect 109217 150454 111215 150456
rect 109217 150451 109283 150454
rect 111149 150451 111215 150454
rect 519905 150242 519971 150245
rect 523200 150242 524400 150272
rect 519905 150240 524400 150242
rect 519905 150184 519910 150240
rect 519966 150184 524400 150240
rect 519905 150182 524400 150184
rect 519905 150179 519971 150182
rect 523200 150152 524400 150182
rect 80605 149698 80671 149701
rect 116393 149698 116459 149701
rect 80605 149696 116459 149698
rect 80605 149640 80610 149696
rect 80666 149640 116398 149696
rect 116454 149640 116459 149696
rect 80605 149638 116459 149640
rect 80605 149635 80671 149638
rect 116393 149635 116459 149638
rect 64689 149562 64755 149565
rect 112897 149562 112963 149565
rect 64689 149560 112963 149562
rect 64689 149504 64694 149560
rect 64750 149504 112902 149560
rect 112958 149504 112963 149560
rect 64689 149502 112963 149504
rect 64689 149499 64755 149502
rect 112897 149499 112963 149502
rect 26969 149426 27035 149429
rect 57881 149426 57947 149429
rect 61469 149426 61535 149429
rect 112713 149426 112779 149429
rect 26969 149424 35910 149426
rect 26969 149368 26974 149424
rect 27030 149368 35910 149424
rect 26969 149366 35910 149368
rect 26969 149363 27035 149366
rect 35850 149154 35910 149366
rect 57881 149424 61394 149426
rect 57881 149368 57886 149424
rect 57942 149368 61394 149424
rect 57881 149366 61394 149368
rect 57881 149363 57947 149366
rect 61334 149290 61394 149366
rect 61469 149424 112779 149426
rect 61469 149368 61474 149424
rect 61530 149368 112718 149424
rect 112774 149368 112779 149424
rect 61469 149366 112779 149368
rect 61469 149363 61535 149366
rect 112713 149363 112779 149366
rect 112529 149290 112595 149293
rect 520917 149290 520983 149293
rect 61334 149288 112595 149290
rect 61334 149232 112534 149288
rect 112590 149232 112595 149288
rect 61334 149230 112595 149232
rect 518788 149288 520983 149290
rect 518788 149232 520922 149288
rect 520978 149232 520983 149288
rect 518788 149230 520983 149232
rect 112529 149227 112595 149230
rect 520917 149227 520983 149230
rect 116577 149154 116643 149157
rect 35850 149152 116643 149154
rect 35850 149096 116582 149152
rect 116638 149096 116643 149152
rect 35850 149094 116643 149096
rect 116577 149091 116643 149094
rect 116117 149018 116183 149021
rect 116117 149016 119140 149018
rect 116117 148960 116122 149016
rect 116178 148960 119140 149016
rect 116117 148958 119140 148960
rect 116117 148955 116183 148958
rect 521101 148746 521167 148749
rect 523200 148746 524400 148776
rect 521101 148744 524400 148746
rect 521101 148688 521106 148744
rect 521162 148688 524400 148744
rect 521101 148686 524400 148688
rect 521101 148683 521167 148686
rect 523200 148656 524400 148686
rect 519537 147930 519603 147933
rect 518788 147928 519603 147930
rect 518788 147872 519542 147928
rect 519598 147872 519603 147928
rect 518788 147870 519603 147872
rect 519537 147867 519603 147870
rect 521193 147386 521259 147389
rect 523200 147386 524400 147416
rect 521193 147384 524400 147386
rect 521193 147328 521198 147384
rect 521254 147328 524400 147384
rect 521193 147326 524400 147328
rect 521193 147323 521259 147326
rect 523200 147296 524400 147326
rect 116485 147114 116551 147117
rect 116485 147112 119140 147114
rect 116485 147056 116490 147112
rect 116546 147056 119140 147112
rect 116485 147054 119140 147056
rect 116485 147051 116551 147054
rect 519629 146570 519695 146573
rect 518788 146568 519695 146570
rect 518788 146512 519634 146568
rect 519690 146512 519695 146568
rect 518788 146510 519695 146512
rect 519629 146507 519695 146510
rect 520917 145890 520983 145893
rect 523200 145890 524400 145920
rect 520917 145888 524400 145890
rect 520917 145832 520922 145888
rect 520978 145832 524400 145888
rect 520917 145830 524400 145832
rect 520917 145827 520983 145830
rect 523200 145800 524400 145830
rect 116025 145210 116091 145213
rect 519721 145210 519787 145213
rect 116025 145208 119140 145210
rect 116025 145152 116030 145208
rect 116086 145152 119140 145208
rect 116025 145150 119140 145152
rect 518788 145208 519787 145210
rect 518788 145152 519726 145208
rect 519782 145152 519787 145208
rect 518788 145150 519787 145152
rect 116025 145147 116091 145150
rect 519721 145147 519787 145150
rect 520273 144394 520339 144397
rect 523200 144394 524400 144424
rect 520273 144392 524400 144394
rect 520273 144336 520278 144392
rect 520334 144336 524400 144392
rect 520273 144334 524400 144336
rect 520273 144331 520339 144334
rect 523200 144304 524400 144334
rect 113817 144258 113883 144261
rect 110860 144256 113883 144258
rect 110860 144200 113822 144256
rect 113878 144200 113883 144256
rect 110860 144198 113883 144200
rect 113817 144195 113883 144198
rect 519813 143850 519879 143853
rect 518788 143848 519879 143850
rect 518788 143792 519818 143848
rect 519874 143792 519879 143848
rect 518788 143790 519879 143792
rect 519813 143787 519879 143790
rect 116117 143306 116183 143309
rect 116117 143304 119140 143306
rect 116117 143248 116122 143304
rect 116178 143248 119140 143304
rect 116117 143246 119140 143248
rect 116117 143243 116183 143246
rect 520733 142898 520799 142901
rect 523200 142898 524400 142928
rect 520733 142896 524400 142898
rect 520733 142840 520738 142896
rect 520794 142840 524400 142896
rect 520733 142838 524400 142840
rect 520733 142835 520799 142838
rect 523200 142808 524400 142838
rect 521009 142490 521075 142493
rect 518788 142488 521075 142490
rect 518788 142432 521014 142488
rect 521070 142432 521075 142488
rect 518788 142430 521075 142432
rect 521009 142427 521075 142430
rect 521009 141402 521075 141405
rect 523200 141402 524400 141432
rect 521009 141400 524400 141402
rect 110321 140858 110387 140861
rect 119110 140858 119170 141372
rect 521009 141344 521014 141400
rect 521070 141344 524400 141400
rect 521009 141342 524400 141344
rect 521009 141339 521075 141342
rect 523200 141312 524400 141342
rect 519905 141130 519971 141133
rect 518788 141128 519971 141130
rect 518788 141072 519910 141128
rect 519966 141072 519971 141128
rect 518788 141070 519971 141072
rect 519905 141067 519971 141070
rect 110321 140856 119170 140858
rect 110321 140800 110326 140856
rect 110382 140800 119170 140856
rect 110321 140798 119170 140800
rect 110321 140795 110387 140798
rect 521285 139906 521351 139909
rect 523200 139906 524400 139936
rect 521285 139904 524400 139906
rect 521285 139848 521290 139904
rect 521346 139848 524400 139904
rect 521285 139846 524400 139848
rect 521285 139843 521351 139846
rect 523200 139816 524400 139846
rect 521101 139770 521167 139773
rect 518788 139768 521167 139770
rect 518788 139712 521106 139768
rect 521162 139712 521167 139768
rect 518788 139710 521167 139712
rect 521101 139707 521167 139710
rect 116117 139498 116183 139501
rect 116117 139496 119140 139498
rect 116117 139440 116122 139496
rect 116178 139440 119140 139496
rect 116117 139438 119140 139440
rect 116117 139435 116183 139438
rect 521193 138410 521259 138413
rect 518788 138408 521259 138410
rect 518788 138352 521198 138408
rect 521254 138352 521259 138408
rect 518788 138350 521259 138352
rect 521193 138347 521259 138350
rect 521377 138410 521443 138413
rect 523200 138410 524400 138440
rect 521377 138408 524400 138410
rect 521377 138352 521382 138408
rect 521438 138352 524400 138408
rect 521377 138350 524400 138352
rect 521377 138347 521443 138350
rect 523200 138320 524400 138350
rect 116117 137594 116183 137597
rect 116117 137592 119140 137594
rect 116117 137536 116122 137592
rect 116178 137536 119140 137592
rect 116117 137534 119140 137536
rect 116117 137531 116183 137534
rect 520917 137050 520983 137053
rect 518788 137048 520983 137050
rect 518788 136992 520922 137048
rect 520978 136992 520983 137048
rect 518788 136990 520983 136992
rect 520917 136987 520983 136990
rect 521193 136914 521259 136917
rect 523200 136914 524400 136944
rect 521193 136912 524400 136914
rect 521193 136856 521198 136912
rect 521254 136856 524400 136912
rect 521193 136854 524400 136856
rect 521193 136851 521259 136854
rect 523200 136824 524400 136854
rect 520273 135690 520339 135693
rect 518788 135688 520339 135690
rect 518788 135632 520278 135688
rect 520334 135632 520339 135688
rect 518788 135630 520339 135632
rect 520273 135627 520339 135630
rect 117221 135554 117287 135557
rect 117221 135552 119140 135554
rect 117221 135496 117226 135552
rect 117282 135496 119140 135552
rect 117221 135494 119140 135496
rect 117221 135491 117287 135494
rect 521101 135418 521167 135421
rect 523200 135418 524400 135448
rect 521101 135416 524400 135418
rect 521101 135360 521106 135416
rect 521162 135360 524400 135416
rect 521101 135358 524400 135360
rect 521101 135355 521167 135358
rect 523200 135328 524400 135358
rect 520733 134330 520799 134333
rect 518788 134328 520799 134330
rect 518788 134272 520738 134328
rect 520794 134272 520799 134328
rect 518788 134270 520799 134272
rect 520733 134267 520799 134270
rect 520273 134058 520339 134061
rect 523200 134058 524400 134088
rect 520273 134056 524400 134058
rect 520273 134000 520278 134056
rect 520334 134000 524400 134056
rect 520273 133998 524400 134000
rect 520273 133995 520339 133998
rect 523200 133968 524400 133998
rect 117129 133650 117195 133653
rect 117129 133648 119140 133650
rect 117129 133592 117134 133648
rect 117190 133592 119140 133648
rect 117129 133590 119140 133592
rect 117129 133587 117195 133590
rect 521009 132970 521075 132973
rect 518788 132968 521075 132970
rect 518788 132912 521014 132968
rect 521070 132912 521075 132968
rect 518788 132910 521075 132912
rect 521009 132907 521075 132910
rect 113909 132834 113975 132837
rect 110860 132832 113975 132834
rect 110860 132776 113914 132832
rect 113970 132776 113975 132832
rect 110860 132774 113975 132776
rect 113909 132771 113975 132774
rect 521009 132562 521075 132565
rect 523200 132562 524400 132592
rect 521009 132560 524400 132562
rect 521009 132504 521014 132560
rect 521070 132504 524400 132560
rect 521009 132502 524400 132504
rect 521009 132499 521075 132502
rect 523200 132472 524400 132502
rect 115933 131746 115999 131749
rect 115933 131744 119140 131746
rect 115933 131688 115938 131744
rect 115994 131688 119140 131744
rect 115933 131686 119140 131688
rect 115933 131683 115999 131686
rect 521285 131610 521351 131613
rect 518788 131608 521351 131610
rect 518788 131552 521290 131608
rect 521346 131552 521351 131608
rect 518788 131550 521351 131552
rect 521285 131547 521351 131550
rect 520181 131066 520247 131069
rect 523200 131066 524400 131096
rect 520181 131064 524400 131066
rect 520181 131008 520186 131064
rect 520242 131008 524400 131064
rect 520181 131006 524400 131008
rect 520181 131003 520247 131006
rect 523200 130976 524400 131006
rect 521377 130250 521443 130253
rect 518788 130248 521443 130250
rect 518788 130192 521382 130248
rect 521438 130192 521443 130248
rect 518788 130190 521443 130192
rect 521377 130187 521443 130190
rect 115933 129842 115999 129845
rect 115933 129840 119140 129842
rect 115933 129784 115938 129840
rect 115994 129784 119140 129840
rect 115933 129782 119140 129784
rect 115933 129779 115999 129782
rect 519905 129570 519971 129573
rect 523200 129570 524400 129600
rect 519905 129568 524400 129570
rect 519905 129512 519910 129568
rect 519966 129512 524400 129568
rect 519905 129510 524400 129512
rect 519905 129507 519971 129510
rect 523200 129480 524400 129510
rect 521193 128890 521259 128893
rect 518788 128888 521259 128890
rect 518788 128832 521198 128888
rect 521254 128832 521259 128888
rect 518788 128830 521259 128832
rect 521193 128827 521259 128830
rect 519537 128074 519603 128077
rect 523200 128074 524400 128104
rect 519537 128072 524400 128074
rect 519537 128016 519542 128072
rect 519598 128016 524400 128072
rect 519537 128014 524400 128016
rect 519537 128011 519603 128014
rect 523200 127984 524400 128014
rect 115197 127938 115263 127941
rect 115197 127936 119140 127938
rect 115197 127880 115202 127936
rect 115258 127880 119140 127936
rect 115197 127878 119140 127880
rect 115197 127875 115263 127878
rect 521101 127530 521167 127533
rect 518788 127528 521167 127530
rect 518788 127472 521106 127528
rect 521162 127472 521167 127528
rect 518788 127470 521167 127472
rect 521101 127467 521167 127470
rect 519721 126578 519787 126581
rect 523200 126578 524400 126608
rect 519721 126576 524400 126578
rect 519721 126520 519726 126576
rect 519782 126520 524400 126576
rect 519721 126518 524400 126520
rect 519721 126515 519787 126518
rect 523200 126488 524400 126518
rect 520273 126170 520339 126173
rect 518788 126168 520339 126170
rect 518788 126112 520278 126168
rect 520334 126112 520339 126168
rect 518788 126110 520339 126112
rect 520273 126107 520339 126110
rect 116117 126034 116183 126037
rect 116117 126032 119140 126034
rect 116117 125976 116122 126032
rect 116178 125976 119140 126032
rect 116117 125974 119140 125976
rect 116117 125971 116183 125974
rect 519813 125082 519879 125085
rect 523200 125082 524400 125112
rect 519813 125080 524400 125082
rect 519813 125024 519818 125080
rect 519874 125024 524400 125080
rect 519813 125022 524400 125024
rect 519813 125019 519879 125022
rect 523200 124992 524400 125022
rect 521009 124810 521075 124813
rect 518788 124808 521075 124810
rect 518788 124752 521014 124808
rect 521070 124752 521075 124808
rect 518788 124750 521075 124752
rect 521009 124747 521075 124750
rect 116117 124130 116183 124133
rect 116117 124128 119140 124130
rect 116117 124072 116122 124128
rect 116178 124072 119140 124128
rect 116117 124070 119140 124072
rect 116117 124067 116183 124070
rect 519261 123586 519327 123589
rect 523200 123586 524400 123616
rect 519261 123584 524400 123586
rect 519261 123528 519266 123584
rect 519322 123528 524400 123584
rect 519261 123526 524400 123528
rect 519261 123523 519327 123526
rect 523200 123496 524400 123526
rect 520181 123450 520247 123453
rect 518788 123448 520247 123450
rect 518788 123392 520186 123448
rect 520242 123392 520247 123448
rect 518788 123390 520247 123392
rect 520181 123387 520247 123390
rect 116117 122226 116183 122229
rect 116117 122224 119140 122226
rect 116117 122168 116122 122224
rect 116178 122168 119140 122224
rect 116117 122166 119140 122168
rect 116117 122163 116183 122166
rect 519905 122090 519971 122093
rect 518788 122088 519971 122090
rect 518788 122032 519910 122088
rect 519966 122032 519971 122088
rect 518788 122030 519971 122032
rect 519905 122027 519971 122030
rect 520089 122090 520155 122093
rect 523200 122090 524400 122120
rect 520089 122088 524400 122090
rect 520089 122032 520094 122088
rect 520150 122032 524400 122088
rect 520089 122030 524400 122032
rect 520089 122027 520155 122030
rect 523200 122000 524400 122030
rect 114001 121410 114067 121413
rect 110860 121408 114067 121410
rect 110860 121352 114006 121408
rect 114062 121352 114067 121408
rect 110860 121350 114067 121352
rect 114001 121347 114067 121350
rect 519537 120730 519603 120733
rect 518788 120728 519603 120730
rect 518788 120672 519542 120728
rect 519598 120672 519603 120728
rect 518788 120670 519603 120672
rect 519537 120667 519603 120670
rect 520181 120730 520247 120733
rect 523200 120730 524400 120760
rect 520181 120728 524400 120730
rect 520181 120672 520186 120728
rect 520242 120672 524400 120728
rect 520181 120670 524400 120672
rect 520181 120667 520247 120670
rect 523200 120640 524400 120670
rect 116117 120186 116183 120189
rect 116117 120184 119140 120186
rect 116117 120128 116122 120184
rect 116178 120128 119140 120184
rect 116117 120126 119140 120128
rect 116117 120123 116183 120126
rect 519721 119370 519787 119373
rect 518788 119368 519787 119370
rect 518788 119312 519726 119368
rect 519782 119312 519787 119368
rect 518788 119310 519787 119312
rect 519721 119307 519787 119310
rect 519905 119234 519971 119237
rect 523200 119234 524400 119264
rect 519905 119232 524400 119234
rect 519905 119176 519910 119232
rect 519966 119176 524400 119232
rect 519905 119174 524400 119176
rect 519905 119171 519971 119174
rect 523200 119144 524400 119174
rect 117037 118282 117103 118285
rect 117037 118280 119140 118282
rect 117037 118224 117042 118280
rect 117098 118224 119140 118280
rect 117037 118222 119140 118224
rect 117037 118219 117103 118222
rect 519813 118010 519879 118013
rect 518788 118008 519879 118010
rect 518788 117952 519818 118008
rect 519874 117952 519879 118008
rect 518788 117950 519879 117952
rect 519813 117947 519879 117950
rect 519721 117738 519787 117741
rect 523200 117738 524400 117768
rect 519721 117736 524400 117738
rect 519721 117680 519726 117736
rect 519782 117680 524400 117736
rect 519721 117678 524400 117680
rect 519721 117675 519787 117678
rect 523200 117648 524400 117678
rect 519261 116650 519327 116653
rect 518788 116648 519327 116650
rect 518788 116592 519266 116648
rect 519322 116592 519327 116648
rect 518788 116590 519327 116592
rect 519261 116587 519327 116590
rect 116945 116378 117011 116381
rect 116945 116376 119140 116378
rect 116945 116320 116950 116376
rect 117006 116320 119140 116376
rect 116945 116318 119140 116320
rect 116945 116315 117011 116318
rect 519997 116242 520063 116245
rect 523200 116242 524400 116272
rect 519997 116240 524400 116242
rect 519997 116184 520002 116240
rect 520058 116184 524400 116240
rect 519997 116182 524400 116184
rect 519997 116179 520063 116182
rect 523200 116152 524400 116182
rect 520089 115290 520155 115293
rect 518788 115288 520155 115290
rect 518788 115232 520094 115288
rect 520150 115232 520155 115288
rect 518788 115230 520155 115232
rect 520089 115227 520155 115230
rect 519813 114746 519879 114749
rect 523200 114746 524400 114776
rect 519813 114744 524400 114746
rect 519813 114688 519818 114744
rect 519874 114688 524400 114744
rect 519813 114686 524400 114688
rect 519813 114683 519879 114686
rect 523200 114656 524400 114686
rect 110321 113250 110387 113253
rect 119110 113250 119170 114444
rect 520181 113930 520247 113933
rect 518788 113928 520247 113930
rect 518788 113872 520186 113928
rect 520242 113872 520247 113928
rect 518788 113870 520247 113872
rect 520181 113867 520247 113870
rect 110321 113248 119170 113250
rect 110321 113192 110326 113248
rect 110382 113192 119170 113248
rect 110321 113190 119170 113192
rect 519261 113250 519327 113253
rect 523200 113250 524400 113280
rect 519261 113248 524400 113250
rect 519261 113192 519266 113248
rect 519322 113192 524400 113248
rect 519261 113190 524400 113192
rect 110321 113187 110387 113190
rect 519261 113187 519327 113190
rect 523200 113160 524400 113190
rect 116853 112570 116919 112573
rect 519905 112570 519971 112573
rect 116853 112568 119140 112570
rect 116853 112512 116858 112568
rect 116914 112512 119140 112568
rect 116853 112510 119140 112512
rect 518788 112568 519971 112570
rect 518788 112512 519910 112568
rect 519966 112512 519971 112568
rect 518788 112510 519971 112512
rect 116853 112507 116919 112510
rect 519905 112507 519971 112510
rect 520089 111754 520155 111757
rect 523200 111754 524400 111784
rect 520089 111752 524400 111754
rect 520089 111696 520094 111752
rect 520150 111696 524400 111752
rect 520089 111694 524400 111696
rect 520089 111691 520155 111694
rect 523200 111664 524400 111694
rect 519721 111210 519787 111213
rect 518788 111208 519787 111210
rect 518788 111152 519726 111208
rect 519782 111152 519787 111208
rect 518788 111150 519787 111152
rect 519721 111147 519787 111150
rect 110321 110666 110387 110669
rect 110321 110664 119140 110666
rect 110321 110608 110326 110664
rect 110382 110608 119140 110664
rect 110321 110606 119140 110608
rect 110321 110603 110387 110606
rect 520181 110258 520247 110261
rect 523200 110258 524400 110288
rect 520181 110256 524400 110258
rect 520181 110200 520186 110256
rect 520242 110200 524400 110256
rect 520181 110198 524400 110200
rect 520181 110195 520247 110198
rect 523200 110168 524400 110198
rect 114093 110122 114159 110125
rect 110860 110120 114159 110122
rect 110860 110064 114098 110120
rect 114154 110064 114159 110120
rect 110860 110062 114159 110064
rect 114093 110059 114159 110062
rect 519997 109850 520063 109853
rect 518788 109848 520063 109850
rect 518788 109792 520002 109848
rect 520058 109792 520063 109848
rect 518788 109790 520063 109792
rect 519997 109787 520063 109790
rect 519629 108762 519695 108765
rect 523200 108762 524400 108792
rect 519629 108760 524400 108762
rect 110321 107674 110387 107677
rect 119110 107674 119170 108732
rect 519629 108704 519634 108760
rect 519690 108704 524400 108760
rect 519629 108702 524400 108704
rect 519629 108699 519695 108702
rect 523200 108672 524400 108702
rect 519813 108490 519879 108493
rect 518788 108488 519879 108490
rect 518788 108432 519818 108488
rect 519874 108432 519879 108488
rect 518788 108430 519879 108432
rect 519813 108427 519879 108430
rect 110321 107672 119170 107674
rect 110321 107616 110326 107672
rect 110382 107616 119170 107672
rect 110321 107614 119170 107616
rect 110321 107611 110387 107614
rect 519721 107402 519787 107405
rect 523200 107402 524400 107432
rect 519721 107400 524400 107402
rect 519721 107344 519726 107400
rect 519782 107344 524400 107400
rect 519721 107342 524400 107344
rect 519721 107339 519787 107342
rect 523200 107312 524400 107342
rect 519261 107130 519327 107133
rect 518788 107128 519327 107130
rect 518788 107072 519266 107128
rect 519322 107072 519327 107128
rect 518788 107070 519327 107072
rect 519261 107067 519327 107070
rect 116117 106858 116183 106861
rect 116117 106856 119140 106858
rect 116117 106800 116122 106856
rect 116178 106800 119140 106856
rect 116117 106798 119140 106800
rect 116117 106795 116183 106798
rect 519905 105906 519971 105909
rect 523200 105906 524400 105936
rect 519905 105904 524400 105906
rect 519905 105848 519910 105904
rect 519966 105848 524400 105904
rect 519905 105846 524400 105848
rect 519905 105843 519971 105846
rect 523200 105816 524400 105846
rect 520089 105770 520155 105773
rect 518788 105768 520155 105770
rect 518788 105712 520094 105768
rect 520150 105712 520155 105768
rect 518788 105710 520155 105712
rect 520089 105707 520155 105710
rect 116117 104818 116183 104821
rect 116117 104816 119140 104818
rect 116117 104760 116122 104816
rect 116178 104760 119140 104816
rect 116117 104758 119140 104760
rect 116117 104755 116183 104758
rect 520181 104546 520247 104549
rect 518758 104544 520247 104546
rect 518758 104488 520186 104544
rect 520242 104488 520247 104544
rect 518758 104486 520247 104488
rect 518758 104380 518818 104486
rect 520181 104483 520247 104486
rect 519077 104410 519143 104413
rect 523200 104410 524400 104440
rect 519077 104408 524400 104410
rect 519077 104352 519082 104408
rect 519138 104352 524400 104408
rect 519077 104350 524400 104352
rect 519077 104347 519143 104350
rect 523200 104320 524400 104350
rect 519629 103050 519695 103053
rect 518788 103048 519695 103050
rect 518788 102992 519634 103048
rect 519690 102992 519695 103048
rect 518788 102990 519695 102992
rect 519629 102987 519695 102990
rect 116761 102914 116827 102917
rect 520089 102914 520155 102917
rect 523200 102914 524400 102944
rect 116761 102912 119140 102914
rect 116761 102856 116766 102912
rect 116822 102856 119140 102912
rect 116761 102854 119140 102856
rect 520089 102912 524400 102914
rect 520089 102856 520094 102912
rect 520150 102856 524400 102912
rect 520089 102854 524400 102856
rect 116761 102851 116827 102854
rect 520089 102851 520155 102854
rect 523200 102824 524400 102854
rect 519721 101690 519787 101693
rect 518788 101688 519787 101690
rect 518788 101632 519726 101688
rect 519782 101632 519787 101688
rect 518788 101630 519787 101632
rect 519721 101627 519787 101630
rect 520181 101418 520247 101421
rect 523200 101418 524400 101448
rect 520181 101416 524400 101418
rect 520181 101360 520186 101416
rect 520242 101360 524400 101416
rect 520181 101358 524400 101360
rect 520181 101355 520247 101358
rect 523200 101328 524400 101358
rect 115933 101010 115999 101013
rect 115933 101008 119140 101010
rect 115933 100952 115938 101008
rect 115994 100952 119140 101008
rect 115933 100950 119140 100952
rect 115933 100947 115999 100950
rect 519905 100330 519971 100333
rect 518788 100328 519971 100330
rect 518788 100272 519910 100328
rect 519966 100272 519971 100328
rect 518788 100270 519971 100272
rect 519905 100267 519971 100270
rect 519445 99922 519511 99925
rect 523200 99922 524400 99952
rect 519445 99920 524400 99922
rect 519445 99864 519450 99920
rect 519506 99864 524400 99920
rect 519445 99862 524400 99864
rect 519445 99859 519511 99862
rect 523200 99832 524400 99862
rect 114185 98698 114251 98701
rect 110860 98696 114251 98698
rect 110860 98640 114190 98696
rect 114246 98640 114251 98696
rect 110860 98638 114251 98640
rect 114185 98635 114251 98638
rect 110321 98154 110387 98157
rect 119110 98154 119170 99076
rect 519077 98970 519143 98973
rect 518788 98968 519143 98970
rect 518788 98912 519082 98968
rect 519138 98912 519143 98968
rect 518788 98910 519143 98912
rect 519077 98907 519143 98910
rect 519813 98426 519879 98429
rect 523200 98426 524400 98456
rect 519813 98424 524400 98426
rect 519813 98368 519818 98424
rect 519874 98368 524400 98424
rect 519813 98366 524400 98368
rect 519813 98363 519879 98366
rect 523200 98336 524400 98366
rect 110321 98152 119170 98154
rect 110321 98096 110326 98152
rect 110382 98096 119170 98152
rect 110321 98094 119170 98096
rect 110321 98091 110387 98094
rect 520089 97610 520155 97613
rect 518788 97608 520155 97610
rect 518788 97552 520094 97608
rect 520150 97552 520155 97608
rect 518788 97550 520155 97552
rect 520089 97547 520155 97550
rect 116209 97202 116275 97205
rect 116209 97200 119140 97202
rect 116209 97144 116214 97200
rect 116270 97144 119140 97200
rect 116209 97142 119140 97144
rect 116209 97139 116275 97142
rect 519537 96930 519603 96933
rect 523200 96930 524400 96960
rect 519537 96928 524400 96930
rect 519537 96872 519542 96928
rect 519598 96872 524400 96928
rect 519537 96870 524400 96872
rect 519537 96867 519603 96870
rect 523200 96840 524400 96870
rect 520181 96250 520247 96253
rect 518788 96248 520247 96250
rect 518788 96192 520186 96248
rect 520242 96192 520247 96248
rect 518788 96190 520247 96192
rect 520181 96187 520247 96190
rect 519721 95434 519787 95437
rect 523200 95434 524400 95464
rect 519721 95432 524400 95434
rect 519721 95376 519726 95432
rect 519782 95376 524400 95432
rect 519721 95374 524400 95376
rect 519721 95371 519787 95374
rect 523200 95344 524400 95374
rect 116117 95298 116183 95301
rect 116117 95296 119140 95298
rect 116117 95240 116122 95296
rect 116178 95240 119140 95296
rect 116117 95238 119140 95240
rect 116117 95235 116183 95238
rect 519445 94890 519511 94893
rect 518788 94888 519511 94890
rect 518788 94832 519450 94888
rect 519506 94832 519511 94888
rect 518788 94830 519511 94832
rect 519445 94827 519511 94830
rect 519077 94074 519143 94077
rect 523200 94074 524400 94104
rect 519077 94072 524400 94074
rect 519077 94016 519082 94072
rect 519138 94016 524400 94072
rect 519077 94014 524400 94016
rect 519077 94011 519143 94014
rect 523200 93984 524400 94014
rect 519813 93530 519879 93533
rect 518788 93528 519879 93530
rect 518788 93472 519818 93528
rect 519874 93472 519879 93528
rect 518788 93470 519879 93472
rect 519813 93467 519879 93470
rect 116117 93394 116183 93397
rect 116117 93392 119140 93394
rect 116117 93336 116122 93392
rect 116178 93336 119140 93392
rect 116117 93334 119140 93336
rect 116117 93331 116183 93334
rect 519261 92578 519327 92581
rect 523200 92578 524400 92608
rect 519261 92576 524400 92578
rect 519261 92520 519266 92576
rect 519322 92520 524400 92576
rect 519261 92518 524400 92520
rect 519261 92515 519327 92518
rect 523200 92488 524400 92518
rect 519537 92170 519603 92173
rect 518788 92168 519603 92170
rect 518788 92112 519542 92168
rect 519598 92112 519603 92168
rect 518788 92110 519603 92112
rect 519537 92107 519603 92110
rect 116577 91354 116643 91357
rect 116577 91352 119140 91354
rect 116577 91296 116582 91352
rect 116638 91296 119140 91352
rect 116577 91294 119140 91296
rect 116577 91291 116643 91294
rect 519445 91082 519511 91085
rect 523200 91082 524400 91112
rect 519445 91080 524400 91082
rect 519445 91024 519450 91080
rect 519506 91024 524400 91080
rect 519445 91022 524400 91024
rect 519445 91019 519511 91022
rect 523200 90992 524400 91022
rect 519721 90810 519787 90813
rect 518788 90808 519787 90810
rect 518788 90752 519726 90808
rect 519782 90752 519787 90808
rect 518788 90750 519787 90752
rect 519721 90747 519787 90750
rect 519905 89586 519971 89589
rect 523200 89586 524400 89616
rect 519905 89584 524400 89586
rect 519905 89528 519910 89584
rect 519966 89528 524400 89584
rect 519905 89526 524400 89528
rect 519905 89523 519971 89526
rect 523200 89496 524400 89526
rect 519077 89450 519143 89453
rect 518788 89448 519143 89450
rect 110321 88362 110387 88365
rect 119110 88362 119170 89420
rect 518788 89392 519082 89448
rect 519138 89392 519143 89448
rect 518788 89390 519143 89392
rect 519077 89387 519143 89390
rect 110321 88360 119170 88362
rect 110321 88304 110326 88360
rect 110382 88304 119170 88360
rect 110321 88302 119170 88304
rect 110321 88299 110387 88302
rect 519261 88090 519327 88093
rect 518788 88088 519327 88090
rect 518788 88032 519266 88088
rect 519322 88032 519327 88088
rect 518788 88030 519327 88032
rect 519261 88027 519327 88030
rect 519997 88090 520063 88093
rect 523200 88090 524400 88120
rect 519997 88088 524400 88090
rect 519997 88032 520002 88088
rect 520058 88032 524400 88088
rect 519997 88030 524400 88032
rect 519997 88027 520063 88030
rect 523200 88000 524400 88030
rect 115933 87546 115999 87549
rect 115933 87544 119140 87546
rect 115933 87488 115938 87544
rect 115994 87488 119140 87544
rect 115933 87486 119140 87488
rect 115933 87483 115999 87486
rect 114277 87274 114343 87277
rect 110860 87272 114343 87274
rect 110860 87216 114282 87272
rect 114338 87216 114343 87272
rect 110860 87214 114343 87216
rect 114277 87211 114343 87214
rect 521561 86730 521627 86733
rect 518788 86728 521627 86730
rect 518788 86672 521566 86728
rect 521622 86672 521627 86728
rect 518788 86670 521627 86672
rect 521561 86667 521627 86670
rect 519721 86594 519787 86597
rect 523200 86594 524400 86624
rect 519721 86592 524400 86594
rect 519721 86536 519726 86592
rect 519782 86536 524400 86592
rect 519721 86534 524400 86536
rect 519721 86531 519787 86534
rect 523200 86504 524400 86534
rect 116393 85642 116459 85645
rect 116393 85640 119140 85642
rect 116393 85584 116398 85640
rect 116454 85584 119140 85640
rect 116393 85582 119140 85584
rect 116393 85579 116459 85582
rect 519445 85370 519511 85373
rect 518788 85368 519511 85370
rect 518788 85312 519450 85368
rect 519506 85312 519511 85368
rect 518788 85310 519511 85312
rect 519445 85307 519511 85310
rect 519077 85098 519143 85101
rect 523200 85098 524400 85128
rect 519077 85096 524400 85098
rect 519077 85040 519082 85096
rect 519138 85040 524400 85096
rect 519077 85038 524400 85040
rect 519077 85035 519143 85038
rect 523200 85008 524400 85038
rect 519905 84010 519971 84013
rect 518788 84008 519971 84010
rect 518788 83952 519910 84008
rect 519966 83952 519971 84008
rect 518788 83950 519971 83952
rect 519905 83947 519971 83950
rect 116577 83738 116643 83741
rect 116577 83736 119140 83738
rect 116577 83680 116582 83736
rect 116638 83680 119140 83736
rect 116577 83678 119140 83680
rect 116577 83675 116643 83678
rect 520089 83602 520155 83605
rect 523200 83602 524400 83632
rect 520089 83600 524400 83602
rect 520089 83544 520094 83600
rect 520150 83544 524400 83600
rect 520089 83542 524400 83544
rect 520089 83539 520155 83542
rect 523200 83512 524400 83542
rect 519997 82650 520063 82653
rect 518788 82648 520063 82650
rect 518788 82592 520002 82648
rect 520058 82592 520063 82648
rect 518788 82590 520063 82592
rect 519997 82587 520063 82590
rect 520181 82106 520247 82109
rect 523200 82106 524400 82136
rect 520181 82104 524400 82106
rect 520181 82048 520186 82104
rect 520242 82048 524400 82104
rect 520181 82046 524400 82048
rect 520181 82043 520247 82046
rect 523200 82016 524400 82046
rect 116301 81834 116367 81837
rect 116301 81832 119140 81834
rect 116301 81776 116306 81832
rect 116362 81776 119140 81832
rect 116301 81774 119140 81776
rect 116301 81771 116367 81774
rect 519721 81290 519787 81293
rect 518788 81288 519787 81290
rect 518788 81232 519726 81288
rect 519782 81232 519787 81288
rect 518788 81230 519787 81232
rect 519721 81227 519787 81230
rect 521101 80746 521167 80749
rect 523200 80746 524400 80776
rect 521101 80744 524400 80746
rect 521101 80688 521106 80744
rect 521162 80688 524400 80744
rect 521101 80686 524400 80688
rect 521101 80683 521167 80686
rect 523200 80656 524400 80686
rect 115933 79930 115999 79933
rect 519077 79930 519143 79933
rect 115933 79928 119140 79930
rect 115933 79872 115938 79928
rect 115994 79872 119140 79928
rect 115933 79870 119140 79872
rect 518788 79928 519143 79930
rect 518788 79872 519082 79928
rect 519138 79872 519143 79928
rect 518788 79870 519143 79872
rect 115933 79867 115999 79870
rect 519077 79867 519143 79870
rect 520549 79250 520615 79253
rect 523200 79250 524400 79280
rect 520549 79248 524400 79250
rect 520549 79192 520554 79248
rect 520610 79192 524400 79248
rect 520549 79190 524400 79192
rect 520549 79187 520615 79190
rect 523200 79160 524400 79190
rect 520089 78570 520155 78573
rect 518788 78568 520155 78570
rect 518788 78512 520094 78568
rect 520150 78512 520155 78568
rect 518788 78510 520155 78512
rect 520089 78507 520155 78510
rect 116209 78026 116275 78029
rect 116209 78024 119140 78026
rect 116209 77968 116214 78024
rect 116270 77968 119140 78024
rect 116209 77966 119140 77968
rect 116209 77963 116275 77966
rect 521009 77754 521075 77757
rect 523200 77754 524400 77784
rect 521009 77752 524400 77754
rect 521009 77696 521014 77752
rect 521070 77696 524400 77752
rect 521009 77694 524400 77696
rect 521009 77691 521075 77694
rect 523200 77664 524400 77694
rect 520181 77210 520247 77213
rect 518788 77208 520247 77210
rect 518788 77152 520186 77208
rect 520242 77152 520247 77208
rect 518788 77150 520247 77152
rect 520181 77147 520247 77150
rect 521193 76258 521259 76261
rect 523200 76258 524400 76288
rect 521193 76256 524400 76258
rect 521193 76200 521198 76256
rect 521254 76200 524400 76256
rect 521193 76198 524400 76200
rect 521193 76195 521259 76198
rect 523200 76168 524400 76198
rect 521101 75986 521167 75989
rect 110860 75926 119140 75986
rect 518788 75984 521167 75986
rect 518788 75928 521106 75984
rect 521162 75928 521167 75984
rect 518788 75926 521167 75928
rect 521101 75923 521167 75926
rect 521101 74762 521167 74765
rect 523200 74762 524400 74792
rect 521101 74760 524400 74762
rect 521101 74704 521106 74760
rect 521162 74704 524400 74760
rect 521101 74702 524400 74704
rect 521101 74699 521167 74702
rect 523200 74672 524400 74702
rect 520549 74626 520615 74629
rect 518788 74624 520615 74626
rect 518788 74568 520554 74624
rect 520610 74568 520615 74624
rect 518788 74566 520615 74568
rect 520549 74563 520615 74566
rect 116669 74082 116735 74085
rect 116669 74080 119140 74082
rect 116669 74024 116674 74080
rect 116730 74024 119140 74080
rect 116669 74022 119140 74024
rect 116669 74019 116735 74022
rect 521009 73810 521075 73813
rect 518758 73808 521075 73810
rect 518758 73752 521014 73808
rect 521070 73752 521075 73808
rect 518758 73750 521075 73752
rect 518758 73236 518818 73750
rect 521009 73747 521075 73750
rect 521009 73266 521075 73269
rect 523200 73266 524400 73296
rect 521009 73264 524400 73266
rect 521009 73208 521014 73264
rect 521070 73208 524400 73264
rect 521009 73206 524400 73208
rect 521009 73203 521075 73206
rect 523200 73176 524400 73206
rect 116577 72178 116643 72181
rect 116577 72176 119140 72178
rect 116577 72120 116582 72176
rect 116638 72120 119140 72176
rect 116577 72118 119140 72120
rect 116577 72115 116643 72118
rect 521193 71906 521259 71909
rect 518788 71904 521259 71906
rect 518788 71848 521198 71904
rect 521254 71848 521259 71904
rect 518788 71846 521259 71848
rect 521193 71843 521259 71846
rect 519997 71770 520063 71773
rect 523200 71770 524400 71800
rect 519997 71768 524400 71770
rect 519997 71712 520002 71768
rect 520058 71712 524400 71768
rect 519997 71710 524400 71712
rect 519997 71707 520063 71710
rect 523200 71680 524400 71710
rect 521101 70546 521167 70549
rect 518788 70544 521167 70546
rect 518788 70488 521106 70544
rect 521162 70488 521167 70544
rect 518788 70486 521167 70488
rect 521101 70483 521167 70486
rect 116301 70274 116367 70277
rect 519261 70274 519327 70277
rect 523200 70274 524400 70304
rect 116301 70272 119140 70274
rect 116301 70216 116306 70272
rect 116362 70216 119140 70272
rect 116301 70214 119140 70216
rect 519261 70272 524400 70274
rect 519261 70216 519266 70272
rect 519322 70216 524400 70272
rect 519261 70214 524400 70216
rect 116301 70211 116367 70214
rect 519261 70211 519327 70214
rect 523200 70184 524400 70214
rect 521009 69186 521075 69189
rect 518788 69184 521075 69186
rect 518788 69128 521014 69184
rect 521070 69128 521075 69184
rect 518788 69126 521075 69128
rect 521009 69123 521075 69126
rect 520181 68778 520247 68781
rect 523200 68778 524400 68808
rect 520181 68776 524400 68778
rect 520181 68720 520186 68776
rect 520242 68720 524400 68776
rect 520181 68718 524400 68720
rect 520181 68715 520247 68718
rect 523200 68688 524400 68718
rect 116117 68370 116183 68373
rect 116117 68368 119140 68370
rect 116117 68312 116122 68368
rect 116178 68312 119140 68368
rect 116117 68310 119140 68312
rect 116117 68307 116183 68310
rect 519997 67826 520063 67829
rect 518788 67824 520063 67826
rect 518788 67768 520002 67824
rect 520058 67768 520063 67824
rect 518788 67766 520063 67768
rect 519997 67763 520063 67766
rect 519905 67418 519971 67421
rect 523200 67418 524400 67448
rect 519905 67416 524400 67418
rect 519905 67360 519910 67416
rect 519966 67360 524400 67416
rect 519905 67358 524400 67360
rect 519905 67355 519971 67358
rect 523200 67328 524400 67358
rect 116577 66466 116643 66469
rect 519261 66466 519327 66469
rect 116577 66464 119140 66466
rect 116577 66408 116582 66464
rect 116638 66408 119140 66464
rect 116577 66406 119140 66408
rect 518788 66464 519327 66466
rect 518788 66408 519266 66464
rect 519322 66408 519327 66464
rect 518788 66406 519327 66408
rect 116577 66403 116643 66406
rect 519261 66403 519327 66406
rect 519813 65922 519879 65925
rect 523200 65922 524400 65952
rect 519813 65920 524400 65922
rect 519813 65864 519818 65920
rect 519874 65864 524400 65920
rect 519813 65862 524400 65864
rect 519813 65859 519879 65862
rect 523200 65832 524400 65862
rect 520181 65106 520247 65109
rect 518788 65104 520247 65106
rect 518788 65048 520186 65104
rect 520242 65048 520247 65104
rect 518788 65046 520247 65048
rect 520181 65043 520247 65046
rect 113357 64562 113423 64565
rect 110860 64560 113423 64562
rect 110860 64504 113362 64560
rect 113418 64504 113423 64560
rect 110860 64502 113423 64504
rect 113357 64499 113423 64502
rect 116209 64562 116275 64565
rect 116209 64560 119140 64562
rect 116209 64504 116214 64560
rect 116270 64504 119140 64560
rect 116209 64502 119140 64504
rect 116209 64499 116275 64502
rect 519077 64426 519143 64429
rect 523200 64426 524400 64456
rect 519077 64424 524400 64426
rect 519077 64368 519082 64424
rect 519138 64368 524400 64424
rect 519077 64366 524400 64368
rect 519077 64363 519143 64366
rect 523200 64336 524400 64366
rect 519905 63746 519971 63749
rect 518788 63744 519971 63746
rect 518788 63688 519910 63744
rect 519966 63688 519971 63744
rect 518788 63686 519971 63688
rect 519905 63683 519971 63686
rect 520089 62930 520155 62933
rect 523200 62930 524400 62960
rect 520089 62928 524400 62930
rect 520089 62872 520094 62928
rect 520150 62872 524400 62928
rect 520089 62870 524400 62872
rect 520089 62867 520155 62870
rect 523200 62840 524400 62870
rect 116117 62658 116183 62661
rect 116117 62656 119140 62658
rect 116117 62600 116122 62656
rect 116178 62600 119140 62656
rect 116117 62598 119140 62600
rect 116117 62595 116183 62598
rect 519813 62386 519879 62389
rect 518788 62384 519879 62386
rect 518788 62328 519818 62384
rect 519874 62328 519879 62384
rect 518788 62326 519879 62328
rect 519813 62323 519879 62326
rect 520181 61434 520247 61437
rect 523200 61434 524400 61464
rect 520181 61432 524400 61434
rect 520181 61376 520186 61432
rect 520242 61376 524400 61432
rect 520181 61374 524400 61376
rect 520181 61371 520247 61374
rect 523200 61344 524400 61374
rect 519077 61026 519143 61029
rect 518788 61024 519143 61026
rect 518788 60968 519082 61024
rect 519138 60968 519143 61024
rect 518788 60966 519143 60968
rect 519077 60963 519143 60966
rect 110321 59394 110387 59397
rect 119110 59394 119170 60588
rect 519077 59938 519143 59941
rect 523200 59938 524400 59968
rect 519077 59936 524400 59938
rect 519077 59880 519082 59936
rect 519138 59880 524400 59936
rect 519077 59878 524400 59880
rect 519077 59875 519143 59878
rect 523200 59848 524400 59878
rect 520089 59666 520155 59669
rect 518788 59664 520155 59666
rect 518788 59608 520094 59664
rect 520150 59608 520155 59664
rect 518788 59606 520155 59608
rect 520089 59603 520155 59606
rect 110321 59392 119170 59394
rect 110321 59336 110326 59392
rect 110382 59336 119170 59392
rect 110321 59334 119170 59336
rect 110321 59331 110387 59334
rect 116577 58714 116643 58717
rect 116577 58712 119140 58714
rect 116577 58656 116582 58712
rect 116638 58656 119140 58712
rect 116577 58654 119140 58656
rect 116577 58651 116643 58654
rect 519997 58442 520063 58445
rect 523200 58442 524400 58472
rect 519997 58440 524400 58442
rect 519997 58384 520002 58440
rect 520058 58384 524400 58440
rect 519997 58382 524400 58384
rect 519997 58379 520063 58382
rect 523200 58352 524400 58382
rect 520181 58306 520247 58309
rect 518788 58304 520247 58306
rect 518788 58248 520186 58304
rect 520242 58248 520247 58304
rect 518788 58246 520247 58248
rect 520181 58243 520247 58246
rect 519077 56946 519143 56949
rect 518788 56944 519143 56946
rect 518788 56888 519082 56944
rect 519138 56888 519143 56944
rect 518788 56886 519143 56888
rect 519077 56883 519143 56886
rect 519445 56946 519511 56949
rect 523200 56946 524400 56976
rect 519445 56944 524400 56946
rect 519445 56888 519450 56944
rect 519506 56888 524400 56944
rect 519445 56886 524400 56888
rect 519445 56883 519511 56886
rect 523200 56856 524400 56886
rect 116669 56810 116735 56813
rect 116669 56808 119140 56810
rect 116669 56752 116674 56808
rect 116730 56752 119140 56808
rect 116669 56750 119140 56752
rect 116669 56747 116735 56750
rect 519997 55586 520063 55589
rect 518788 55584 520063 55586
rect 518788 55528 520002 55584
rect 520058 55528 520063 55584
rect 518788 55526 520063 55528
rect 519997 55523 520063 55526
rect 519813 55450 519879 55453
rect 523200 55450 524400 55480
rect 519813 55448 524400 55450
rect 519813 55392 519818 55448
rect 519874 55392 524400 55448
rect 519813 55390 524400 55392
rect 519813 55387 519879 55390
rect 523200 55360 524400 55390
rect 110321 53954 110387 53957
rect 119110 53954 119170 54876
rect 519445 54226 519511 54229
rect 518788 54224 519511 54226
rect 518788 54168 519450 54224
rect 519506 54168 519511 54224
rect 518788 54166 519511 54168
rect 519445 54163 519511 54166
rect 519997 54090 520063 54093
rect 523200 54090 524400 54120
rect 519997 54088 524400 54090
rect 519997 54032 520002 54088
rect 520058 54032 524400 54088
rect 519997 54030 524400 54032
rect 519997 54027 520063 54030
rect 523200 54000 524400 54030
rect 110321 53952 119170 53954
rect 110321 53896 110326 53952
rect 110382 53896 119170 53952
rect 110321 53894 119170 53896
rect 110321 53891 110387 53894
rect 114185 53138 114251 53141
rect 110860 53136 114251 53138
rect 110860 53080 114190 53136
rect 114246 53080 114251 53136
rect 110860 53078 114251 53080
rect 114185 53075 114251 53078
rect 116761 53002 116827 53005
rect 116761 53000 119140 53002
rect 116761 52944 116766 53000
rect 116822 52944 119140 53000
rect 116761 52942 119140 52944
rect 116761 52939 116827 52942
rect 519813 52866 519879 52869
rect 518788 52864 519879 52866
rect 518788 52808 519818 52864
rect 519874 52808 519879 52864
rect 518788 52806 519879 52808
rect 519813 52803 519879 52806
rect 520089 52594 520155 52597
rect 523200 52594 524400 52624
rect 520089 52592 524400 52594
rect 520089 52536 520094 52592
rect 520150 52536 524400 52592
rect 520089 52534 524400 52536
rect 520089 52531 520155 52534
rect 523200 52504 524400 52534
rect 519997 51506 520063 51509
rect 518788 51504 520063 51506
rect 518788 51448 520002 51504
rect 520058 51448 520063 51504
rect 518788 51446 520063 51448
rect 519997 51443 520063 51446
rect 110321 51098 110387 51101
rect 520181 51098 520247 51101
rect 523200 51098 524400 51128
rect 110321 51096 119140 51098
rect 110321 51040 110326 51096
rect 110382 51040 119140 51096
rect 110321 51038 119140 51040
rect 520181 51096 524400 51098
rect 520181 51040 520186 51096
rect 520242 51040 524400 51096
rect 520181 51038 524400 51040
rect 110321 51035 110387 51038
rect 520181 51035 520247 51038
rect 523200 51008 524400 51038
rect 520089 50146 520155 50149
rect 518788 50144 520155 50146
rect 518788 50088 520094 50144
rect 520150 50088 520155 50144
rect 518788 50086 520155 50088
rect 520089 50083 520155 50086
rect 521101 49602 521167 49605
rect 523200 49602 524400 49632
rect 521101 49600 524400 49602
rect 521101 49544 521106 49600
rect 521162 49544 524400 49600
rect 521101 49542 524400 49544
rect 521101 49539 521167 49542
rect 523200 49512 524400 49542
rect 110321 48378 110387 48381
rect 119110 48378 119170 49164
rect 520181 48786 520247 48789
rect 518788 48784 520247 48786
rect 518788 48728 520186 48784
rect 520242 48728 520247 48784
rect 518788 48726 520247 48728
rect 520181 48723 520247 48726
rect 110321 48376 119170 48378
rect 110321 48320 110326 48376
rect 110382 48320 119170 48376
rect 110321 48318 119170 48320
rect 110321 48315 110387 48318
rect 520917 48106 520983 48109
rect 523200 48106 524400 48136
rect 520917 48104 524400 48106
rect 520917 48048 520922 48104
rect 520978 48048 524400 48104
rect 520917 48046 524400 48048
rect 520917 48043 520983 48046
rect 523200 48016 524400 48046
rect 521101 47426 521167 47429
rect 518788 47424 521167 47426
rect 518788 47368 521106 47424
rect 521162 47368 521167 47424
rect 518788 47366 521167 47368
rect 521101 47363 521167 47366
rect 110321 47154 110387 47157
rect 110321 47152 119140 47154
rect 110321 47096 110326 47152
rect 110382 47096 119140 47152
rect 110321 47094 119140 47096
rect 110321 47091 110387 47094
rect 520917 46746 520983 46749
rect 518758 46744 520983 46746
rect 518758 46688 520922 46744
rect 520978 46688 520983 46744
rect 518758 46686 520983 46688
rect 518758 46036 518818 46686
rect 520917 46683 520983 46686
rect 521561 46610 521627 46613
rect 523200 46610 524400 46640
rect 521561 46608 524400 46610
rect 521561 46552 521566 46608
rect 521622 46552 524400 46608
rect 521561 46550 524400 46552
rect 521561 46547 521627 46550
rect 523200 46520 524400 46550
rect 521561 45658 521627 45661
rect 521561 45656 521670 45658
rect 521561 45600 521566 45656
rect 521622 45600 521670 45656
rect 521561 45595 521670 45600
rect 521610 45386 521670 45595
rect 518758 45326 521670 45386
rect 116117 45250 116183 45253
rect 116117 45248 119140 45250
rect 116117 45192 116122 45248
rect 116178 45192 119140 45248
rect 116117 45190 119140 45192
rect 116117 45187 116183 45190
rect 518758 44676 518818 45326
rect 521101 45114 521167 45117
rect 523200 45114 524400 45144
rect 521101 45112 524400 45114
rect 521101 45056 521106 45112
rect 521162 45056 524400 45112
rect 521101 45054 524400 45056
rect 521101 45051 521167 45054
rect 523200 45024 524400 45054
rect 521101 44026 521167 44029
rect 518758 44024 521167 44026
rect 518758 43968 521106 44024
rect 521162 43968 521167 44024
rect 518758 43966 521167 43968
rect 518758 43316 518818 43966
rect 521101 43963 521167 43966
rect 520917 43618 520983 43621
rect 523200 43618 524400 43648
rect 520917 43616 524400 43618
rect 520917 43560 520922 43616
rect 520978 43560 524400 43616
rect 520917 43558 524400 43560
rect 520917 43555 520983 43558
rect 523200 43528 524400 43558
rect 110321 42938 110387 42941
rect 119110 42938 119170 43316
rect 110321 42936 119170 42938
rect 110321 42880 110326 42936
rect 110382 42880 119170 42936
rect 110321 42878 119170 42880
rect 110321 42875 110387 42878
rect 520917 42666 520983 42669
rect 518758 42664 520983 42666
rect 518758 42608 520922 42664
rect 520978 42608 520983 42664
rect 518758 42606 520983 42608
rect 518758 41956 518818 42606
rect 520917 42603 520983 42606
rect 521101 42122 521167 42125
rect 523200 42122 524400 42152
rect 521101 42120 524400 42122
rect 521101 42064 521106 42120
rect 521162 42064 524400 42120
rect 521101 42062 524400 42064
rect 521101 42059 521167 42062
rect 523200 42032 524400 42062
rect 114093 41850 114159 41853
rect 110860 41848 114159 41850
rect 110860 41792 114098 41848
rect 114154 41792 114159 41848
rect 110860 41790 114159 41792
rect 114093 41787 114159 41790
rect 116945 41442 117011 41445
rect 116945 41440 119140 41442
rect 116945 41384 116950 41440
rect 117006 41384 119140 41440
rect 116945 41382 119140 41384
rect 116945 41379 117011 41382
rect 521101 41306 521167 41309
rect 518758 41304 521167 41306
rect 518758 41248 521106 41304
rect 521162 41248 521167 41304
rect 518758 41246 521167 41248
rect 518758 40596 518818 41246
rect 521101 41243 521167 41246
rect 521101 40762 521167 40765
rect 523200 40762 524400 40792
rect 521101 40760 524400 40762
rect 521101 40704 521106 40760
rect 521162 40704 524400 40760
rect 521101 40702 524400 40704
rect 521101 40699 521167 40702
rect 523200 40672 524400 40702
rect 521101 39946 521167 39949
rect 518758 39944 521167 39946
rect 518758 39888 521106 39944
rect 521162 39888 521167 39944
rect 518758 39886 521167 39888
rect 115197 39538 115263 39541
rect 115197 39536 119140 39538
rect 115197 39480 115202 39536
rect 115258 39480 119140 39536
rect 115197 39478 119140 39480
rect 115197 39475 115263 39478
rect 518758 39236 518818 39886
rect 521101 39883 521167 39886
rect 521101 39266 521167 39269
rect 523200 39266 524400 39296
rect 521101 39264 524400 39266
rect 521101 39208 521106 39264
rect 521162 39208 524400 39264
rect 521101 39206 524400 39208
rect 521101 39203 521167 39206
rect 523200 39176 524400 39206
rect 521101 37906 521167 37909
rect 518788 37904 521167 37906
rect 518788 37848 521106 37904
rect 521162 37848 521167 37904
rect 518788 37846 521167 37848
rect 521101 37843 521167 37846
rect 523200 37770 524400 37800
rect 521150 37710 524400 37770
rect 117129 37634 117195 37637
rect 117129 37632 119140 37634
rect 117129 37576 117134 37632
rect 117190 37576 119140 37632
rect 117129 37574 119140 37576
rect 117129 37571 117195 37574
rect 521150 37226 521210 37710
rect 523200 37680 524400 37710
rect 518758 37166 521210 37226
rect 518758 36516 518818 37166
rect 523200 36274 524400 36304
rect 521610 36214 524400 36274
rect 521610 35866 521670 36214
rect 523200 36184 524400 36214
rect 518758 35806 521670 35866
rect 115933 35730 115999 35733
rect 115933 35728 119140 35730
rect 115933 35672 115938 35728
rect 115994 35672 119140 35728
rect 115933 35670 119140 35672
rect 115933 35667 115999 35670
rect 518758 35156 518818 35806
rect 523200 34778 524400 34808
rect 518850 34718 524400 34778
rect 518850 34506 518910 34718
rect 523200 34688 524400 34718
rect 518758 34446 518910 34506
rect 115933 33826 115999 33829
rect 115933 33824 119140 33826
rect 115933 33768 115938 33824
rect 115994 33768 119140 33824
rect 518758 33796 518818 34446
rect 115933 33766 119140 33768
rect 115933 33763 115999 33766
rect 523200 33282 524400 33312
rect 518850 33222 524400 33282
rect 518850 33146 518910 33222
rect 523200 33192 524400 33222
rect 518758 33086 518910 33146
rect 518758 32436 518818 33086
rect 115289 31786 115355 31789
rect 523200 31786 524400 31816
rect 115289 31784 119140 31786
rect 115289 31728 115294 31784
rect 115350 31728 119140 31784
rect 115289 31726 119140 31728
rect 518850 31726 524400 31786
rect 115289 31723 115355 31726
rect 518850 31650 518910 31726
rect 523200 31696 524400 31726
rect 518758 31590 518910 31650
rect 518758 31076 518818 31590
rect 114001 30426 114067 30429
rect 110860 30424 114067 30426
rect 110860 30368 114006 30424
rect 114062 30368 114067 30424
rect 110860 30366 114067 30368
rect 114001 30363 114067 30366
rect 520917 30290 520983 30293
rect 523200 30290 524400 30320
rect 520917 30288 524400 30290
rect 520917 30232 520922 30288
rect 520978 30232 524400 30288
rect 520917 30230 524400 30232
rect 520917 30227 520983 30230
rect 523200 30200 524400 30230
rect 116117 29882 116183 29885
rect 116117 29880 119140 29882
rect 116117 29824 116122 29880
rect 116178 29824 119140 29880
rect 116117 29822 119140 29824
rect 116117 29819 116183 29822
rect 518758 29066 518818 29716
rect 520917 29066 520983 29069
rect 518758 29064 520983 29066
rect 518758 29008 520922 29064
rect 520978 29008 520983 29064
rect 518758 29006 520983 29008
rect 520917 29003 520983 29006
rect 521101 28794 521167 28797
rect 523200 28794 524400 28824
rect 521101 28792 524400 28794
rect 521101 28736 521106 28792
rect 521162 28736 524400 28792
rect 521101 28734 524400 28736
rect 521101 28731 521167 28734
rect 523200 28704 524400 28734
rect 115381 27978 115447 27981
rect 115381 27976 119140 27978
rect 115381 27920 115386 27976
rect 115442 27920 119140 27976
rect 115381 27918 119140 27920
rect 115381 27915 115447 27918
rect 518758 27706 518818 28356
rect 521101 27706 521167 27709
rect 518758 27704 521167 27706
rect 518758 27648 521106 27704
rect 521162 27648 521167 27704
rect 518758 27646 521167 27648
rect 521101 27643 521167 27646
rect 521101 27434 521167 27437
rect 523200 27434 524400 27464
rect 521101 27432 524400 27434
rect 521101 27376 521106 27432
rect 521162 27376 524400 27432
rect 521101 27374 524400 27376
rect 521101 27371 521167 27374
rect 523200 27344 524400 27374
rect 518758 26346 518818 26996
rect 521101 26346 521167 26349
rect 518758 26344 521167 26346
rect 518758 26288 521106 26344
rect 521162 26288 521167 26344
rect 518758 26286 521167 26288
rect 521101 26283 521167 26286
rect 116117 26074 116183 26077
rect 116117 26072 119140 26074
rect 116117 26016 116122 26072
rect 116178 26016 119140 26072
rect 116117 26014 119140 26016
rect 116117 26011 116183 26014
rect 520917 25938 520983 25941
rect 523200 25938 524400 25968
rect 520917 25936 524400 25938
rect 520917 25880 520922 25936
rect 520978 25880 524400 25936
rect 520917 25878 524400 25880
rect 520917 25875 520983 25878
rect 523200 25848 524400 25878
rect 518758 24986 518818 25636
rect 520917 24986 520983 24989
rect 518758 24984 520983 24986
rect 518758 24928 520922 24984
rect 520978 24928 520983 24984
rect 518758 24926 520983 24928
rect 520917 24923 520983 24926
rect 519077 24442 519143 24445
rect 523200 24442 524400 24472
rect 519077 24440 524400 24442
rect 519077 24384 519082 24440
rect 519138 24384 524400 24440
rect 519077 24382 524400 24384
rect 519077 24379 519143 24382
rect 523200 24352 524400 24382
rect 115933 24170 115999 24173
rect 115933 24168 119140 24170
rect 115933 24112 115938 24168
rect 115994 24112 119140 24168
rect 115933 24110 119140 24112
rect 115933 24107 115999 24110
rect 518758 23626 518818 24276
rect 519077 23626 519143 23629
rect 518758 23624 519143 23626
rect 518758 23568 519082 23624
rect 519138 23568 519143 23624
rect 518758 23566 519143 23568
rect 519077 23563 519143 23566
rect 521101 22946 521167 22949
rect 523200 22946 524400 22976
rect 521101 22944 524400 22946
rect 116117 22266 116183 22269
rect 518758 22266 518818 22916
rect 521101 22888 521106 22944
rect 521162 22888 524400 22944
rect 521101 22886 524400 22888
rect 521101 22883 521167 22886
rect 523200 22856 524400 22886
rect 521101 22266 521167 22269
rect 116117 22264 119140 22266
rect 116117 22208 116122 22264
rect 116178 22208 119140 22264
rect 116117 22206 119140 22208
rect 518758 22264 521167 22266
rect 518758 22208 521106 22264
rect 521162 22208 521167 22264
rect 518758 22206 521167 22208
rect 116117 22203 116183 22206
rect 521101 22203 521167 22206
rect 518758 20906 518818 21556
rect 523200 21450 524400 21480
rect 521150 21390 524400 21450
rect 521150 20906 521210 21390
rect 523200 21360 524400 21390
rect 518758 20846 521210 20906
rect 116853 20362 116919 20365
rect 116853 20360 119140 20362
rect 116853 20304 116858 20360
rect 116914 20304 119140 20360
rect 116853 20302 119140 20304
rect 116853 20299 116919 20302
rect 518758 19546 518818 20196
rect 523200 19954 524400 19984
rect 521150 19894 524400 19954
rect 521150 19546 521210 19894
rect 523200 19864 524400 19894
rect 518758 19486 521210 19546
rect 113909 19002 113975 19005
rect 110860 19000 113975 19002
rect 110860 18944 113914 19000
rect 113970 18944 113975 19000
rect 110860 18942 113975 18944
rect 113909 18939 113975 18942
rect 117037 18458 117103 18461
rect 117037 18456 119140 18458
rect 117037 18400 117042 18456
rect 117098 18400 119140 18456
rect 117037 18398 119140 18400
rect 117037 18395 117103 18398
rect 518758 18186 518818 18836
rect 523200 18458 524400 18488
rect 521150 18398 524400 18458
rect 521150 18186 521210 18398
rect 523200 18368 524400 18398
rect 518758 18126 521210 18186
rect 518758 16826 518818 17476
rect 523200 16962 524400 16992
rect 521150 16902 524400 16962
rect 521150 16826 521210 16902
rect 523200 16872 524400 16902
rect 518758 16766 521210 16826
rect 117221 16418 117287 16421
rect 117221 16416 119140 16418
rect 117221 16360 117226 16416
rect 117282 16360 119140 16416
rect 117221 16358 119140 16360
rect 117221 16355 117287 16358
rect 518758 15466 518818 16116
rect 523200 15466 524400 15496
rect 518758 15406 524400 15466
rect 523200 15376 524400 15406
rect 116485 14514 116551 14517
rect 116485 14512 119140 14514
rect 116485 14456 116490 14512
rect 116546 14456 119140 14512
rect 116485 14454 119140 14456
rect 116485 14451 116551 14454
rect 518758 14106 518818 14756
rect 523200 14106 524400 14136
rect 518758 14046 524400 14106
rect 523200 14016 524400 14046
rect 518758 12746 518818 13396
rect 518758 12686 518910 12746
rect 116209 12610 116275 12613
rect 518850 12610 518910 12686
rect 523200 12610 524400 12640
rect 116209 12608 119140 12610
rect 116209 12552 116214 12608
rect 116270 12552 119140 12608
rect 116209 12550 119140 12552
rect 518850 12550 524400 12610
rect 116209 12547 116275 12550
rect 523200 12520 524400 12550
rect 518758 11386 518818 12036
rect 518758 11326 518910 11386
rect 518850 11114 518910 11326
rect 523200 11114 524400 11144
rect 518850 11054 524400 11114
rect 523200 11024 524400 11054
rect 116117 10706 116183 10709
rect 521101 10706 521167 10709
rect 116117 10704 119140 10706
rect 116117 10648 116122 10704
rect 116178 10648 119140 10704
rect 116117 10646 119140 10648
rect 518788 10704 521167 10706
rect 518788 10648 521106 10704
rect 521162 10648 521167 10704
rect 518788 10646 521167 10648
rect 116117 10643 116183 10646
rect 521101 10643 521167 10646
rect 521101 9618 521167 9621
rect 523200 9618 524400 9648
rect 521101 9616 524400 9618
rect 521101 9560 521106 9616
rect 521162 9560 524400 9616
rect 521101 9558 524400 9560
rect 521101 9555 521167 9558
rect 523200 9528 524400 9558
rect 520917 9346 520983 9349
rect 518788 9344 520983 9346
rect 518788 9288 520922 9344
rect 520978 9288 520983 9344
rect 518788 9286 520983 9288
rect 520917 9283 520983 9286
rect 117037 8802 117103 8805
rect 117037 8800 119140 8802
rect 117037 8744 117042 8800
rect 117098 8744 119140 8800
rect 117037 8742 119140 8744
rect 117037 8739 117103 8742
rect 520917 8122 520983 8125
rect 523200 8122 524400 8152
rect 520917 8120 524400 8122
rect 520917 8064 520922 8120
rect 520978 8064 524400 8120
rect 520917 8062 524400 8064
rect 520917 8059 520983 8062
rect 523200 8032 524400 8062
rect 520273 7986 520339 7989
rect 518788 7984 520339 7986
rect 518788 7928 520278 7984
rect 520334 7928 520339 7984
rect 518788 7926 520339 7928
rect 520273 7923 520339 7926
rect 113817 7714 113883 7717
rect 110860 7712 113883 7714
rect 110860 7656 113822 7712
rect 113878 7656 113883 7712
rect 110860 7654 113883 7656
rect 113817 7651 113883 7654
rect 115933 6898 115999 6901
rect 115933 6896 119140 6898
rect 115933 6840 115938 6896
rect 115994 6840 119140 6896
rect 115933 6838 119140 6840
rect 115933 6835 115999 6838
rect 520273 6626 520339 6629
rect 523200 6626 524400 6656
rect 518788 6566 520106 6626
rect 520046 6490 520106 6566
rect 520273 6624 524400 6626
rect 520273 6568 520278 6624
rect 520334 6568 524400 6624
rect 520273 6566 524400 6568
rect 520273 6563 520339 6566
rect 523200 6536 524400 6566
rect 521101 6490 521167 6493
rect 520046 6488 521167 6490
rect 520046 6432 521106 6488
rect 521162 6432 521167 6488
rect 520046 6430 521167 6432
rect 521101 6427 521167 6430
rect 521009 5266 521075 5269
rect 518788 5264 521075 5266
rect 518788 5208 521014 5264
rect 521070 5208 521075 5264
rect 518788 5206 521075 5208
rect 521009 5203 521075 5206
rect 521101 5130 521167 5133
rect 523200 5130 524400 5160
rect 521101 5128 524400 5130
rect 521101 5072 521106 5128
rect 521162 5072 524400 5128
rect 521101 5070 524400 5072
rect 521101 5067 521167 5070
rect 523200 5040 524400 5070
rect 116117 4994 116183 4997
rect 116117 4992 119140 4994
rect 116117 4936 116122 4992
rect 116178 4936 119140 4992
rect 116117 4934 119140 4936
rect 116117 4931 116183 4934
rect 110137 4042 110203 4045
rect 93810 4040 110203 4042
rect 93810 3984 110142 4040
rect 110198 3984 110203 4040
rect 93810 3982 110203 3984
rect 84150 3302 89730 3362
rect 84150 2954 84210 3302
rect 89670 3226 89730 3302
rect 93810 3226 93870 3982
rect 110137 3979 110203 3982
rect 521193 3906 521259 3909
rect 518788 3904 521259 3906
rect 518788 3848 521198 3904
rect 521254 3848 521259 3904
rect 518788 3846 521259 3848
rect 521193 3843 521259 3846
rect 116853 3770 116919 3773
rect 100710 3768 116919 3770
rect 100710 3712 116858 3768
rect 116914 3712 116919 3768
rect 100710 3710 116919 3712
rect 100710 3362 100770 3710
rect 116853 3707 116919 3710
rect 109401 3634 109467 3637
rect 116761 3634 116827 3637
rect 109401 3632 116827 3634
rect 109401 3576 109406 3632
rect 109462 3576 116766 3632
rect 116822 3576 116827 3632
rect 109401 3574 116827 3576
rect 109401 3571 109467 3574
rect 116761 3571 116827 3574
rect 521009 3634 521075 3637
rect 523200 3634 524400 3664
rect 521009 3632 524400 3634
rect 521009 3576 521014 3632
rect 521070 3576 524400 3632
rect 521009 3574 524400 3576
rect 521009 3571 521075 3574
rect 523200 3544 524400 3574
rect 109493 3498 109559 3501
rect 117129 3498 117195 3501
rect 109493 3496 117195 3498
rect 109493 3440 109498 3496
rect 109554 3440 117134 3496
rect 117190 3440 117195 3496
rect 109493 3438 117195 3440
rect 109493 3435 109559 3438
rect 117129 3435 117195 3438
rect 89670 3166 93870 3226
rect 100296 3302 100770 3362
rect 89670 3030 98332 3090
rect 89670 2954 89730 3030
rect 76238 2894 84210 2954
rect 88934 2894 89730 2954
rect 33182 2758 76114 2818
rect 33041 2682 33107 2685
rect 33182 2682 33242 2758
rect 33041 2680 33242 2682
rect 33041 2624 33046 2680
rect 33102 2624 33242 2680
rect 33041 2622 33242 2624
rect 33041 2619 33107 2622
rect 76054 2546 76114 2758
rect 76238 2685 76298 2894
rect 76189 2680 76298 2685
rect 76189 2624 76194 2680
rect 76250 2624 76298 2680
rect 76189 2622 76298 2624
rect 76422 2758 88810 2818
rect 76189 2619 76255 2622
rect 76422 2546 76482 2758
rect 76054 2486 76482 2546
rect 88750 2546 88810 2758
rect 88934 2685 88994 2894
rect 88885 2680 88994 2685
rect 88885 2624 88890 2680
rect 88946 2624 88994 2680
rect 88885 2622 88994 2624
rect 89118 2758 93870 2818
rect 88885 2619 88951 2622
rect 89118 2546 89178 2758
rect 88750 2486 89178 2546
rect 93810 2546 93870 2758
rect 98272 2685 98332 3030
rect 100296 2685 100356 3302
rect 109401 3226 109467 3229
rect 108990 3224 109467 3226
rect 108990 3168 109406 3224
rect 109462 3168 109467 3224
rect 108990 3166 109467 3168
rect 108990 3090 109050 3166
rect 109401 3163 109467 3166
rect 102182 3030 109050 3090
rect 116117 3090 116183 3093
rect 116117 3088 119140 3090
rect 116117 3032 116122 3088
rect 116178 3032 119140 3088
rect 116117 3030 119140 3032
rect 102182 2685 102242 3030
rect 116117 3027 116183 3030
rect 110137 2954 110203 2957
rect 102366 2952 110203 2954
rect 102366 2896 110142 2952
rect 110198 2896 110203 2952
rect 102366 2894 110203 2896
rect 102366 2685 102426 2894
rect 110137 2891 110203 2894
rect 111057 2818 111123 2821
rect 98269 2680 98335 2685
rect 98269 2624 98274 2680
rect 98330 2624 98335 2680
rect 98269 2619 98335 2624
rect 100293 2680 100359 2685
rect 100293 2624 100298 2680
rect 100354 2624 100359 2680
rect 100293 2619 100359 2624
rect 102133 2680 102242 2685
rect 102133 2624 102138 2680
rect 102194 2624 102242 2680
rect 102133 2622 102242 2624
rect 102317 2680 102426 2685
rect 102317 2624 102322 2680
rect 102378 2624 102426 2680
rect 102317 2622 102426 2624
rect 103470 2816 111123 2818
rect 103470 2760 111062 2816
rect 111118 2760 111123 2816
rect 103470 2758 111123 2760
rect 102133 2619 102199 2622
rect 102317 2619 102383 2622
rect 103470 2546 103530 2758
rect 111057 2755 111123 2758
rect 521101 2682 521167 2685
rect 518788 2680 521167 2682
rect 518788 2624 521106 2680
rect 521162 2624 521167 2680
rect 518788 2622 521167 2624
rect 521101 2619 521167 2622
rect 93810 2486 103530 2546
rect 94405 2410 94471 2413
rect 102133 2410 102199 2413
rect 94405 2408 102199 2410
rect 94405 2352 94410 2408
rect 94466 2352 102138 2408
rect 102194 2352 102199 2408
rect 94405 2350 102199 2352
rect 94405 2347 94471 2350
rect 102133 2347 102199 2350
rect 98269 2274 98335 2277
rect 109493 2274 109559 2277
rect 98269 2272 109559 2274
rect 98269 2216 98274 2272
rect 98330 2216 109498 2272
rect 109554 2216 109559 2272
rect 98269 2214 109559 2216
rect 98269 2211 98335 2214
rect 109493 2211 109559 2214
rect 26049 2138 26115 2141
rect 117221 2138 117287 2141
rect 26049 2136 117287 2138
rect 26049 2080 26054 2136
rect 26110 2080 117226 2136
rect 117282 2080 117287 2136
rect 26049 2078 117287 2080
rect 26049 2075 26115 2078
rect 117221 2075 117287 2078
rect 521193 2138 521259 2141
rect 523200 2138 524400 2168
rect 521193 2136 524400 2138
rect 521193 2080 521198 2136
rect 521254 2080 524400 2136
rect 521193 2078 524400 2080
rect 521193 2075 521259 2078
rect 523200 2048 524400 2078
rect 22921 2002 22987 2005
rect 116485 2002 116551 2005
rect 22921 2000 116551 2002
rect 22921 1944 22926 2000
rect 22982 1944 116490 2000
rect 116546 1944 116551 2000
rect 22921 1942 116551 1944
rect 22921 1939 22987 1942
rect 116485 1939 116551 1942
rect 19333 1866 19399 1869
rect 116209 1866 116275 1869
rect 19333 1864 116275 1866
rect 19333 1808 19338 1864
rect 19394 1808 116214 1864
rect 116270 1808 116275 1864
rect 19333 1806 116275 1808
rect 19333 1803 19399 1806
rect 116209 1803 116275 1806
rect 15929 1730 15995 1733
rect 116025 1730 116091 1733
rect 15929 1728 116091 1730
rect 15929 1672 15934 1728
rect 15990 1672 116030 1728
rect 116086 1672 116091 1728
rect 15929 1670 116091 1672
rect 15929 1667 15995 1670
rect 116025 1667 116091 1670
rect 229277 1730 229343 1733
rect 293585 1730 293651 1733
rect 229277 1728 293651 1730
rect 229277 1672 229282 1728
rect 229338 1672 293590 1728
rect 293646 1672 293651 1728
rect 229277 1670 293651 1672
rect 229277 1667 229343 1670
rect 293585 1667 293651 1670
rect 12617 1594 12683 1597
rect 117037 1594 117103 1597
rect 12617 1592 117103 1594
rect 12617 1536 12622 1592
rect 12678 1536 117042 1592
rect 117098 1536 117103 1592
rect 12617 1534 117103 1536
rect 12617 1531 12683 1534
rect 117037 1531 117103 1534
rect 163773 1594 163839 1597
rect 243629 1594 243695 1597
rect 163773 1592 243695 1594
rect 163773 1536 163778 1592
rect 163834 1536 243634 1592
rect 243690 1536 243695 1592
rect 163773 1534 243695 1536
rect 163773 1531 163839 1534
rect 243629 1531 243695 1534
rect 55949 1458 56015 1461
rect 294781 1458 294847 1461
rect 55949 1456 294847 1458
rect 55949 1400 55954 1456
rect 56010 1400 294786 1456
rect 294842 1400 294847 1456
rect 55949 1398 294847 1400
rect 55949 1395 56015 1398
rect 294781 1395 294847 1398
rect 360285 1458 360351 1461
rect 393589 1458 393655 1461
rect 360285 1456 393655 1458
rect 360285 1400 360290 1456
rect 360346 1400 393594 1456
rect 393650 1400 393655 1456
rect 360285 1398 393655 1400
rect 360285 1395 360351 1398
rect 393589 1395 393655 1398
rect 98269 1322 98335 1325
rect 102317 1322 102383 1325
rect 98269 1320 102383 1322
rect 98269 1264 98274 1320
rect 98330 1264 102322 1320
rect 102378 1264 102383 1320
rect 98269 1262 102383 1264
rect 98269 1259 98335 1262
rect 102317 1259 102383 1262
rect 521101 778 521167 781
rect 523200 778 524400 808
rect 521101 776 524400 778
rect 521101 720 521106 776
rect 521162 720 524400 776
rect 521101 718 524400 720
rect 521101 715 521167 718
rect 523200 688 524400 718
<< metal4 >>
rect 1664 144454 1984 144496
rect 1664 144218 1706 144454
rect 1942 144218 1984 144454
rect 1664 144134 1984 144218
rect 1664 143898 1706 144134
rect 1942 143898 1984 144134
rect 1664 143856 1984 143898
rect 109956 144454 110276 144496
rect 109956 144218 109998 144454
rect 110234 144218 110276 144454
rect 109956 144134 110276 144218
rect 109956 143898 109998 144134
rect 110234 143898 110276 144134
rect 109956 143856 110276 143898
rect 119664 144454 119984 144496
rect 119664 144218 119706 144454
rect 119942 144218 119984 144454
rect 119664 144134 119984 144218
rect 119664 143898 119706 144134
rect 119942 143898 119984 144134
rect 119664 143856 119984 143898
rect 517940 144454 518260 144496
rect 517940 144218 517982 144454
rect 518218 144218 518260 144454
rect 517940 144134 518260 144218
rect 517940 143898 517982 144134
rect 518218 143898 518260 144134
rect 517940 143856 518260 143898
rect 1096 131454 1332 131496
rect 1096 131134 1332 131218
rect 1096 130856 1332 130898
rect 110616 131454 110936 131496
rect 110616 131218 110658 131454
rect 110894 131218 110936 131454
rect 110616 131134 110936 131218
rect 110616 130898 110658 131134
rect 110894 130898 110936 131134
rect 110616 130856 110936 130898
rect 119004 131454 119324 131496
rect 119004 131218 119046 131454
rect 119282 131218 119324 131454
rect 119004 131134 119324 131218
rect 119004 130898 119046 131134
rect 119282 130898 119324 131134
rect 119004 130856 119324 130898
rect 518600 131454 518920 131496
rect 518600 131218 518642 131454
rect 518878 131218 518920 131454
rect 518600 131134 518920 131218
rect 518600 130898 518642 131134
rect 518878 130898 518920 131134
rect 518600 130856 518920 130898
rect 1664 118454 1984 118496
rect 1664 118218 1706 118454
rect 1942 118218 1984 118454
rect 1664 118134 1984 118218
rect 1664 117898 1706 118134
rect 1942 117898 1984 118134
rect 1664 117856 1984 117898
rect 109956 118454 110276 118496
rect 109956 118218 109998 118454
rect 110234 118218 110276 118454
rect 109956 118134 110276 118218
rect 109956 117898 109998 118134
rect 110234 117898 110276 118134
rect 109956 117856 110276 117898
rect 119664 118454 119984 118496
rect 119664 118218 119706 118454
rect 119942 118218 119984 118454
rect 119664 118134 119984 118218
rect 119664 117898 119706 118134
rect 119942 117898 119984 118134
rect 119664 117856 119984 117898
rect 517940 118454 518260 118496
rect 517940 118218 517982 118454
rect 518218 118218 518260 118454
rect 517940 118134 518260 118218
rect 517940 117898 517982 118134
rect 518218 117898 518260 118134
rect 517940 117856 518260 117898
rect 1096 105454 1332 105496
rect 1096 105134 1332 105218
rect 1096 104856 1332 104898
rect 110616 105454 110936 105496
rect 110616 105218 110658 105454
rect 110894 105218 110936 105454
rect 110616 105134 110936 105218
rect 110616 104898 110658 105134
rect 110894 104898 110936 105134
rect 110616 104856 110936 104898
rect 119004 105454 119324 105496
rect 119004 105218 119046 105454
rect 119282 105218 119324 105454
rect 119004 105134 119324 105218
rect 119004 104898 119046 105134
rect 119282 104898 119324 105134
rect 119004 104856 119324 104898
rect 518600 105454 518920 105496
rect 518600 105218 518642 105454
rect 518878 105218 518920 105454
rect 518600 105134 518920 105218
rect 518600 104898 518642 105134
rect 518878 104898 518920 105134
rect 518600 104856 518920 104898
rect 1664 92454 1984 92496
rect 1664 92218 1706 92454
rect 1942 92218 1984 92454
rect 1664 92134 1984 92218
rect 1664 91898 1706 92134
rect 1942 91898 1984 92134
rect 1664 91856 1984 91898
rect 109956 92454 110276 92496
rect 109956 92218 109998 92454
rect 110234 92218 110276 92454
rect 109956 92134 110276 92218
rect 109956 91898 109998 92134
rect 110234 91898 110276 92134
rect 109956 91856 110276 91898
rect 119664 92454 119984 92496
rect 119664 92218 119706 92454
rect 119942 92218 119984 92454
rect 119664 92134 119984 92218
rect 119664 91898 119706 92134
rect 119942 91898 119984 92134
rect 119664 91856 119984 91898
rect 517940 92454 518260 92496
rect 517940 92218 517982 92454
rect 518218 92218 518260 92454
rect 517940 92134 518260 92218
rect 517940 91898 517982 92134
rect 518218 91898 518260 92134
rect 517940 91856 518260 91898
rect 1096 79454 1332 79496
rect 1096 79134 1332 79218
rect 1096 78856 1332 78898
rect 110616 79454 110936 79496
rect 110616 79218 110658 79454
rect 110894 79218 110936 79454
rect 110616 79134 110936 79218
rect 110616 78898 110658 79134
rect 110894 78898 110936 79134
rect 110616 78856 110936 78898
rect 119004 79454 119324 79496
rect 119004 79218 119046 79454
rect 119282 79218 119324 79454
rect 119004 79134 119324 79218
rect 119004 78898 119046 79134
rect 119282 78898 119324 79134
rect 119004 78856 119324 78898
rect 518600 79454 518920 79496
rect 518600 79218 518642 79454
rect 518878 79218 518920 79454
rect 518600 79134 518920 79218
rect 518600 78898 518642 79134
rect 518878 78898 518920 79134
rect 518600 78856 518920 78898
rect 1664 66454 1984 66496
rect 1664 66218 1706 66454
rect 1942 66218 1984 66454
rect 1664 66134 1984 66218
rect 1664 65898 1706 66134
rect 1942 65898 1984 66134
rect 1664 65856 1984 65898
rect 109956 66454 110276 66496
rect 109956 66218 109998 66454
rect 110234 66218 110276 66454
rect 109956 66134 110276 66218
rect 109956 65898 109998 66134
rect 110234 65898 110276 66134
rect 109956 65856 110276 65898
rect 119664 66454 119984 66496
rect 119664 66218 119706 66454
rect 119942 66218 119984 66454
rect 119664 66134 119984 66218
rect 119664 65898 119706 66134
rect 119942 65898 119984 66134
rect 119664 65856 119984 65898
rect 517940 66454 518260 66496
rect 517940 66218 517982 66454
rect 518218 66218 518260 66454
rect 517940 66134 518260 66218
rect 517940 65898 517982 66134
rect 518218 65898 518260 66134
rect 517940 65856 518260 65898
rect 1096 53454 1332 53496
rect 1096 53134 1332 53218
rect 1096 52856 1332 52898
rect 110616 53454 110936 53496
rect 110616 53218 110658 53454
rect 110894 53218 110936 53454
rect 110616 53134 110936 53218
rect 110616 52898 110658 53134
rect 110894 52898 110936 53134
rect 110616 52856 110936 52898
rect 119004 53454 119324 53496
rect 119004 53218 119046 53454
rect 119282 53218 119324 53454
rect 119004 53134 119324 53218
rect 119004 52898 119046 53134
rect 119282 52898 119324 53134
rect 119004 52856 119324 52898
rect 518600 53454 518920 53496
rect 518600 53218 518642 53454
rect 518878 53218 518920 53454
rect 518600 53134 518920 53218
rect 518600 52898 518642 53134
rect 518878 52898 518920 53134
rect 518600 52856 518920 52898
rect 1664 40454 1984 40496
rect 1664 40218 1706 40454
rect 1942 40218 1984 40454
rect 1664 40134 1984 40218
rect 1664 39898 1706 40134
rect 1942 39898 1984 40134
rect 1664 39856 1984 39898
rect 109956 40454 110276 40496
rect 109956 40218 109998 40454
rect 110234 40218 110276 40454
rect 109956 40134 110276 40218
rect 109956 39898 109998 40134
rect 110234 39898 110276 40134
rect 109956 39856 110276 39898
rect 119664 40454 119984 40496
rect 119664 40218 119706 40454
rect 119942 40218 119984 40454
rect 119664 40134 119984 40218
rect 119664 39898 119706 40134
rect 119942 39898 119984 40134
rect 119664 39856 119984 39898
rect 517940 40454 518260 40496
rect 517940 40218 517982 40454
rect 518218 40218 518260 40454
rect 517940 40134 518260 40218
rect 517940 39898 517982 40134
rect 518218 39898 518260 40134
rect 517940 39856 518260 39898
rect 1096 27454 1332 27496
rect 1096 27134 1332 27218
rect 1096 26856 1332 26898
rect 110616 27454 110936 27496
rect 110616 27218 110658 27454
rect 110894 27218 110936 27454
rect 110616 27134 110936 27218
rect 110616 26898 110658 27134
rect 110894 26898 110936 27134
rect 110616 26856 110936 26898
rect 119004 27454 119324 27496
rect 119004 27218 119046 27454
rect 119282 27218 119324 27454
rect 119004 27134 119324 27218
rect 119004 26898 119046 27134
rect 119282 26898 119324 27134
rect 119004 26856 119324 26898
rect 518600 27454 518920 27496
rect 518600 27218 518642 27454
rect 518878 27218 518920 27454
rect 518600 27134 518920 27218
rect 518600 26898 518642 27134
rect 518878 26898 518920 27134
rect 518600 26856 518920 26898
rect 1664 14454 1984 14496
rect 1664 14218 1706 14454
rect 1942 14218 1984 14454
rect 1664 14134 1984 14218
rect 1664 13898 1706 14134
rect 1942 13898 1984 14134
rect 1664 13856 1984 13898
rect 109956 14454 110276 14496
rect 109956 14218 109998 14454
rect 110234 14218 110276 14454
rect 109956 14134 110276 14218
rect 109956 13898 109998 14134
rect 110234 13898 110276 14134
rect 109956 13856 110276 13898
rect 119664 14454 119984 14496
rect 119664 14218 119706 14454
rect 119942 14218 119984 14454
rect 119664 14134 119984 14218
rect 119664 13898 119706 14134
rect 119942 13898 119984 14134
rect 119664 13856 119984 13898
rect 517940 14454 518260 14496
rect 517940 14218 517982 14454
rect 518218 14218 518260 14454
rect 517940 14134 518260 14218
rect 517940 13898 517982 14134
rect 518218 13898 518260 14134
rect 517940 13856 518260 13898
<< via4 >>
rect 1706 144218 1942 144454
rect 1706 143898 1942 144134
rect 109998 144218 110234 144454
rect 109998 143898 110234 144134
rect 119706 144218 119942 144454
rect 119706 143898 119942 144134
rect 517982 144218 518218 144454
rect 517982 143898 518218 144134
rect 1096 131218 1332 131454
rect 1096 130898 1332 131134
rect 110658 131218 110894 131454
rect 110658 130898 110894 131134
rect 119046 131218 119282 131454
rect 119046 130898 119282 131134
rect 518642 131218 518878 131454
rect 518642 130898 518878 131134
rect 1706 118218 1942 118454
rect 1706 117898 1942 118134
rect 109998 118218 110234 118454
rect 109998 117898 110234 118134
rect 119706 118218 119942 118454
rect 119706 117898 119942 118134
rect 517982 118218 518218 118454
rect 517982 117898 518218 118134
rect 1096 105218 1332 105454
rect 1096 104898 1332 105134
rect 110658 105218 110894 105454
rect 110658 104898 110894 105134
rect 119046 105218 119282 105454
rect 119046 104898 119282 105134
rect 518642 105218 518878 105454
rect 518642 104898 518878 105134
rect 1706 92218 1942 92454
rect 1706 91898 1942 92134
rect 109998 92218 110234 92454
rect 109998 91898 110234 92134
rect 119706 92218 119942 92454
rect 119706 91898 119942 92134
rect 517982 92218 518218 92454
rect 517982 91898 518218 92134
rect 1096 79218 1332 79454
rect 1096 78898 1332 79134
rect 110658 79218 110894 79454
rect 110658 78898 110894 79134
rect 119046 79218 119282 79454
rect 119046 78898 119282 79134
rect 518642 79218 518878 79454
rect 518642 78898 518878 79134
rect 1706 66218 1942 66454
rect 1706 65898 1942 66134
rect 109998 66218 110234 66454
rect 109998 65898 110234 66134
rect 119706 66218 119942 66454
rect 119706 65898 119942 66134
rect 517982 66218 518218 66454
rect 517982 65898 518218 66134
rect 1096 53218 1332 53454
rect 1096 52898 1332 53134
rect 110658 53218 110894 53454
rect 110658 52898 110894 53134
rect 119046 53218 119282 53454
rect 119046 52898 119282 53134
rect 518642 53218 518878 53454
rect 518642 52898 518878 53134
rect 1706 40218 1942 40454
rect 1706 39898 1942 40134
rect 109998 40218 110234 40454
rect 109998 39898 110234 40134
rect 119706 40218 119942 40454
rect 119706 39898 119942 40134
rect 517982 40218 518218 40454
rect 517982 39898 518218 40134
rect 1096 27218 1332 27454
rect 1096 26898 1332 27134
rect 110658 27218 110894 27454
rect 110658 26898 110894 27134
rect 119046 27218 119282 27454
rect 119046 26898 119282 27134
rect 518642 27218 518878 27454
rect 518642 26898 518878 27134
rect 1706 14218 1942 14454
rect 1706 13898 1942 14134
rect 109998 14218 110234 14454
rect 109998 13898 110234 14134
rect 119706 14218 119942 14454
rect 119706 13898 119942 14134
rect 517982 14218 518218 14454
rect 517982 13898 518218 14134
<< metal5 >>
rect 1104 144454 2200 144496
rect 1104 144218 1706 144454
rect 1942 144218 2200 144454
rect 1104 144134 2200 144218
rect 1104 143898 1706 144134
rect 1942 143898 2200 144134
rect 1104 143856 2200 143898
rect 109800 144454 120200 144496
rect 109800 144218 109998 144454
rect 110234 144218 119706 144454
rect 119942 144218 120200 144454
rect 109800 144134 120200 144218
rect 109800 143898 109998 144134
rect 110234 143898 119706 144134
rect 119942 143898 120200 144134
rect 109800 143856 120200 143898
rect 517800 144454 522836 144496
rect 517800 144218 517982 144454
rect 518218 144218 522836 144454
rect 517800 144134 522836 144218
rect 517800 143898 517982 144134
rect 518218 143898 522836 144134
rect 517800 143856 522836 143898
rect 1072 131454 2200 131496
rect 1072 131218 1096 131454
rect 1332 131218 2200 131454
rect 1072 131134 2200 131218
rect 1072 130898 1096 131134
rect 1332 130898 2200 131134
rect 1072 130856 2200 130898
rect 109800 131454 120200 131496
rect 109800 131218 110658 131454
rect 110894 131218 119046 131454
rect 119282 131218 120200 131454
rect 109800 131134 120200 131218
rect 109800 130898 110658 131134
rect 110894 130898 119046 131134
rect 119282 130898 120200 131134
rect 109800 130856 120200 130898
rect 517800 131454 522836 131496
rect 517800 131218 518642 131454
rect 518878 131218 522836 131454
rect 517800 131134 522836 131218
rect 517800 130898 518642 131134
rect 518878 130898 522836 131134
rect 517800 130856 522836 130898
rect 1104 118454 2200 118496
rect 1104 118218 1706 118454
rect 1942 118218 2200 118454
rect 1104 118134 2200 118218
rect 1104 117898 1706 118134
rect 1942 117898 2200 118134
rect 1104 117856 2200 117898
rect 109800 118454 120200 118496
rect 109800 118218 109998 118454
rect 110234 118218 119706 118454
rect 119942 118218 120200 118454
rect 109800 118134 120200 118218
rect 109800 117898 109998 118134
rect 110234 117898 119706 118134
rect 119942 117898 120200 118134
rect 109800 117856 120200 117898
rect 517800 118454 522836 118496
rect 517800 118218 517982 118454
rect 518218 118218 522836 118454
rect 517800 118134 522836 118218
rect 517800 117898 517982 118134
rect 518218 117898 522836 118134
rect 517800 117856 522836 117898
rect 1072 105454 2200 105496
rect 1072 105218 1096 105454
rect 1332 105218 2200 105454
rect 1072 105134 2200 105218
rect 1072 104898 1096 105134
rect 1332 104898 2200 105134
rect 1072 104856 2200 104898
rect 109800 105454 120200 105496
rect 109800 105218 110658 105454
rect 110894 105218 119046 105454
rect 119282 105218 120200 105454
rect 109800 105134 120200 105218
rect 109800 104898 110658 105134
rect 110894 104898 119046 105134
rect 119282 104898 120200 105134
rect 109800 104856 120200 104898
rect 517800 105454 522836 105496
rect 517800 105218 518642 105454
rect 518878 105218 522836 105454
rect 517800 105134 522836 105218
rect 517800 104898 518642 105134
rect 518878 104898 522836 105134
rect 517800 104856 522836 104898
rect 1104 92454 2200 92496
rect 1104 92218 1706 92454
rect 1942 92218 2200 92454
rect 1104 92134 2200 92218
rect 1104 91898 1706 92134
rect 1942 91898 2200 92134
rect 1104 91856 2200 91898
rect 109800 92454 120200 92496
rect 109800 92218 109998 92454
rect 110234 92218 119706 92454
rect 119942 92218 120200 92454
rect 109800 92134 120200 92218
rect 109800 91898 109998 92134
rect 110234 91898 119706 92134
rect 119942 91898 120200 92134
rect 109800 91856 120200 91898
rect 517800 92454 522836 92496
rect 517800 92218 517982 92454
rect 518218 92218 522836 92454
rect 517800 92134 522836 92218
rect 517800 91898 517982 92134
rect 518218 91898 522836 92134
rect 517800 91856 522836 91898
rect 1072 79454 2200 79496
rect 1072 79218 1096 79454
rect 1332 79218 2200 79454
rect 1072 79134 2200 79218
rect 1072 78898 1096 79134
rect 1332 78898 2200 79134
rect 1072 78856 2200 78898
rect 109800 79454 120200 79496
rect 109800 79218 110658 79454
rect 110894 79218 119046 79454
rect 119282 79218 120200 79454
rect 109800 79134 120200 79218
rect 109800 78898 110658 79134
rect 110894 78898 119046 79134
rect 119282 78898 120200 79134
rect 109800 78856 120200 78898
rect 517800 79454 522836 79496
rect 517800 79218 518642 79454
rect 518878 79218 522836 79454
rect 517800 79134 522836 79218
rect 517800 78898 518642 79134
rect 518878 78898 522836 79134
rect 517800 78856 522836 78898
rect 1104 66454 2200 66496
rect 1104 66218 1706 66454
rect 1942 66218 2200 66454
rect 1104 66134 2200 66218
rect 1104 65898 1706 66134
rect 1942 65898 2200 66134
rect 1104 65856 2200 65898
rect 109800 66454 120200 66496
rect 109800 66218 109998 66454
rect 110234 66218 119706 66454
rect 119942 66218 120200 66454
rect 109800 66134 120200 66218
rect 109800 65898 109998 66134
rect 110234 65898 119706 66134
rect 119942 65898 120200 66134
rect 109800 65856 120200 65898
rect 517800 66454 522836 66496
rect 517800 66218 517982 66454
rect 518218 66218 522836 66454
rect 517800 66134 522836 66218
rect 517800 65898 517982 66134
rect 518218 65898 522836 66134
rect 517800 65856 522836 65898
rect 1072 53454 2200 53496
rect 1072 53218 1096 53454
rect 1332 53218 2200 53454
rect 1072 53134 2200 53218
rect 1072 52898 1096 53134
rect 1332 52898 2200 53134
rect 1072 52856 2200 52898
rect 109800 53454 120200 53496
rect 109800 53218 110658 53454
rect 110894 53218 119046 53454
rect 119282 53218 120200 53454
rect 109800 53134 120200 53218
rect 109800 52898 110658 53134
rect 110894 52898 119046 53134
rect 119282 52898 120200 53134
rect 109800 52856 120200 52898
rect 517800 53454 522836 53496
rect 517800 53218 518642 53454
rect 518878 53218 522836 53454
rect 517800 53134 522836 53218
rect 517800 52898 518642 53134
rect 518878 52898 522836 53134
rect 517800 52856 522836 52898
rect 1104 40454 2200 40496
rect 1104 40218 1706 40454
rect 1942 40218 2200 40454
rect 1104 40134 2200 40218
rect 1104 39898 1706 40134
rect 1942 39898 2200 40134
rect 1104 39856 2200 39898
rect 109800 40454 120200 40496
rect 109800 40218 109998 40454
rect 110234 40218 119706 40454
rect 119942 40218 120200 40454
rect 109800 40134 120200 40218
rect 109800 39898 109998 40134
rect 110234 39898 119706 40134
rect 119942 39898 120200 40134
rect 109800 39856 120200 39898
rect 517800 40454 522836 40496
rect 517800 40218 517982 40454
rect 518218 40218 522836 40454
rect 517800 40134 522836 40218
rect 517800 39898 517982 40134
rect 518218 39898 522836 40134
rect 517800 39856 522836 39898
rect 1072 27454 2200 27496
rect 1072 27218 1096 27454
rect 1332 27218 2200 27454
rect 1072 27134 2200 27218
rect 1072 26898 1096 27134
rect 1332 26898 2200 27134
rect 1072 26856 2200 26898
rect 109800 27454 120200 27496
rect 109800 27218 110658 27454
rect 110894 27218 119046 27454
rect 119282 27218 120200 27454
rect 109800 27134 120200 27218
rect 109800 26898 110658 27134
rect 110894 26898 119046 27134
rect 119282 26898 120200 27134
rect 109800 26856 120200 26898
rect 517800 27454 522836 27496
rect 517800 27218 518642 27454
rect 518878 27218 522836 27454
rect 517800 27134 522836 27218
rect 517800 26898 518642 27134
rect 518878 26898 522836 27134
rect 517800 26856 522836 26898
rect 1104 14454 2200 14496
rect 1104 14218 1706 14454
rect 1942 14218 2200 14454
rect 1104 14134 2200 14218
rect 1104 13898 1706 14134
rect 1942 13898 2200 14134
rect 1104 13856 2200 13898
rect 109800 14454 120200 14496
rect 109800 14218 109998 14454
rect 110234 14218 119706 14454
rect 119942 14218 120200 14454
rect 109800 14134 120200 14218
rect 109800 13898 109998 14134
rect 110234 13898 119706 14134
rect 119942 13898 120200 14134
rect 109800 13856 120200 13898
rect 517800 14454 522836 14496
rect 517800 14218 517982 14454
rect 518218 14218 522836 14454
rect 517800 14134 522836 14218
rect 517800 13898 517982 14134
rect 518218 13898 522836 14134
rect 517800 13856 522836 13898
use mgmt_core  core
timestamp 1638311292
transform 1 0 119000 0 1 2000
box 0 0 400000 148000
use DFFRAM  DFFRAM
timestamp 1638311292
transform 1 0 1000 0 1 2000
box 4 0 110000 148000
<< labels >>
rlabel metal5 s 1104 26856 2200 27496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 26856 120200 27496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 26856 522836 27496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 52856 2200 53496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 52856 120200 53496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 52856 522836 53496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 78856 2200 79496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 78856 120200 79496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 78856 522836 79496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 104856 2200 105496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 104856 120200 105496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 104856 522836 105496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 130856 2200 131496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 130856 120200 131496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 130856 522836 131496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 13856 2200 14496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 13856 120200 14496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 13856 522836 14496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 39856 2200 40496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 39856 120200 40496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 39856 522836 40496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 65856 2200 66496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 65856 120200 66496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 65856 522836 66496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 91856 2200 92496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 91856 120200 92496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 91856 522836 92496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 117856 2200 118496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 117856 120200 118496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 117856 522836 118496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 143856 2200 144496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 143856 120200 144496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 143856 522836 144496 6 VPWR
port 1 nsew power input
rlabel metal2 s 294786 -400 294842 800 6 core_clk
port 2 nsew signal input
rlabel metal2 s 98274 -400 98330 800 6 core_rstn
port 3 nsew signal input
rlabel metal3 s 523200 62840 524400 62960 6 debug_in
port 4 nsew signal input
rlabel metal3 s 523200 64336 524400 64456 6 debug_mode
port 5 nsew signal tristate
rlabel metal3 s 523200 65832 524400 65952 6 debug_oeb
port 6 nsew signal tristate
rlabel metal3 s 523200 67328 524400 67448 6 debug_out
port 7 nsew signal tristate
rlabel metal3 s 523200 141312 524400 141432 6 flash_clk
port 8 nsew signal tristate
rlabel metal3 s 523200 139816 524400 139936 6 flash_csb
port 9 nsew signal tristate
rlabel metal3 s 523200 142808 524400 142928 6 flash_io0_di
port 10 nsew signal input
rlabel metal3 s 523200 144304 524400 144424 6 flash_io0_do
port 11 nsew signal tristate
rlabel metal3 s 523200 145800 524400 145920 6 flash_io0_oeb
port 12 nsew signal tristate
rlabel metal3 s 523200 147296 524400 147416 6 flash_io1_di
port 13 nsew signal input
rlabel metal3 s 523200 148656 524400 148776 6 flash_io1_do
port 14 nsew signal tristate
rlabel metal3 s 523200 150152 524400 150272 6 flash_io1_oeb
port 15 nsew signal tristate
rlabel metal3 s 523200 151648 524400 151768 6 flash_io2_di
port 16 nsew signal input
rlabel metal3 s 523200 153144 524400 153264 6 flash_io2_do
port 17 nsew signal tristate
rlabel metal3 s 523200 154640 524400 154760 6 flash_io2_oeb
port 18 nsew signal tristate
rlabel metal3 s 523200 156136 524400 156256 6 flash_io3_di
port 19 nsew signal input
rlabel metal3 s 523200 157632 524400 157752 6 flash_io3_do
port 20 nsew signal tristate
rlabel metal3 s 523200 159128 524400 159248 6 flash_io3_oeb
port 21 nsew signal tristate
rlabel metal2 s 32770 -400 32826 800 6 gpio_in_pad
port 22 nsew signal input
rlabel metal2 s 163778 -400 163834 800 6 gpio_inenb_pad
port 23 nsew signal tristate
rlabel metal2 s 229282 -400 229338 800 6 gpio_mode0_pad
port 24 nsew signal tristate
rlabel metal2 s 360290 -400 360346 800 6 gpio_mode1_pad
port 25 nsew signal tristate
rlabel metal2 s 425794 -400 425850 800 6 gpio_out_pad
port 26 nsew signal tristate
rlabel metal2 s 491298 -400 491354 800 6 gpio_outenb_pad
port 27 nsew signal tristate
rlabel metal3 s 523200 89496 524400 89616 6 hk_ack_i
port 28 nsew signal input
rlabel metal2 s 523498 159200 523554 160400 6 hk_cyc_o
port 29 nsew signal tristate
rlabel metal3 s 523200 92488 524400 92608 6 hk_dat_i[0]
port 30 nsew signal input
rlabel metal3 s 523200 107312 524400 107432 6 hk_dat_i[10]
port 31 nsew signal input
rlabel metal3 s 523200 108672 524400 108792 6 hk_dat_i[11]
port 32 nsew signal input
rlabel metal3 s 523200 110168 524400 110288 6 hk_dat_i[12]
port 33 nsew signal input
rlabel metal3 s 523200 111664 524400 111784 6 hk_dat_i[13]
port 34 nsew signal input
rlabel metal3 s 523200 113160 524400 113280 6 hk_dat_i[14]
port 35 nsew signal input
rlabel metal3 s 523200 114656 524400 114776 6 hk_dat_i[15]
port 36 nsew signal input
rlabel metal3 s 523200 116152 524400 116272 6 hk_dat_i[16]
port 37 nsew signal input
rlabel metal3 s 523200 117648 524400 117768 6 hk_dat_i[17]
port 38 nsew signal input
rlabel metal3 s 523200 119144 524400 119264 6 hk_dat_i[18]
port 39 nsew signal input
rlabel metal3 s 523200 120640 524400 120760 6 hk_dat_i[19]
port 40 nsew signal input
rlabel metal3 s 523200 93984 524400 94104 6 hk_dat_i[1]
port 41 nsew signal input
rlabel metal3 s 523200 122000 524400 122120 6 hk_dat_i[20]
port 42 nsew signal input
rlabel metal3 s 523200 123496 524400 123616 6 hk_dat_i[21]
port 43 nsew signal input
rlabel metal3 s 523200 124992 524400 125112 6 hk_dat_i[22]
port 44 nsew signal input
rlabel metal3 s 523200 126488 524400 126608 6 hk_dat_i[23]
port 45 nsew signal input
rlabel metal3 s 523200 127984 524400 128104 6 hk_dat_i[24]
port 46 nsew signal input
rlabel metal3 s 523200 129480 524400 129600 6 hk_dat_i[25]
port 47 nsew signal input
rlabel metal3 s 523200 130976 524400 131096 6 hk_dat_i[26]
port 48 nsew signal input
rlabel metal3 s 523200 132472 524400 132592 6 hk_dat_i[27]
port 49 nsew signal input
rlabel metal3 s 523200 133968 524400 134088 6 hk_dat_i[28]
port 50 nsew signal input
rlabel metal3 s 523200 135328 524400 135448 6 hk_dat_i[29]
port 51 nsew signal input
rlabel metal3 s 523200 95344 524400 95464 6 hk_dat_i[2]
port 52 nsew signal input
rlabel metal3 s 523200 136824 524400 136944 6 hk_dat_i[30]
port 53 nsew signal input
rlabel metal3 s 523200 138320 524400 138440 6 hk_dat_i[31]
port 54 nsew signal input
rlabel metal3 s 523200 96840 524400 96960 6 hk_dat_i[3]
port 55 nsew signal input
rlabel metal3 s 523200 98336 524400 98456 6 hk_dat_i[4]
port 56 nsew signal input
rlabel metal3 s 523200 99832 524400 99952 6 hk_dat_i[5]
port 57 nsew signal input
rlabel metal3 s 523200 101328 524400 101448 6 hk_dat_i[6]
port 58 nsew signal input
rlabel metal3 s 523200 102824 524400 102944 6 hk_dat_i[7]
port 59 nsew signal input
rlabel metal3 s 523200 104320 524400 104440 6 hk_dat_i[8]
port 60 nsew signal input
rlabel metal3 s 523200 105816 524400 105936 6 hk_dat_i[9]
port 61 nsew signal input
rlabel metal3 s 523200 90992 524400 91112 6 hk_stb_o
port 62 nsew signal tristate
rlabel metal2 s 521014 159200 521070 160400 6 irq[0]
port 63 nsew signal input
rlabel metal2 s 521842 159200 521898 160400 6 irq[1]
port 64 nsew signal input
rlabel metal2 s 522670 159200 522726 160400 6 irq[2]
port 65 nsew signal input
rlabel metal3 s 523200 73176 524400 73296 6 irq[3]
port 66 nsew signal input
rlabel metal3 s 523200 71680 524400 71800 6 irq[4]
port 67 nsew signal input
rlabel metal3 s 523200 70184 524400 70304 6 irq[5]
port 68 nsew signal input
rlabel metal2 s 386 159200 442 160400 6 la_iena[0]
port 69 nsew signal tristate
rlabel metal2 s 336278 159200 336334 160400 6 la_iena[100]
port 70 nsew signal tristate
rlabel metal2 s 339590 159200 339646 160400 6 la_iena[101]
port 71 nsew signal tristate
rlabel metal2 s 342994 159200 343050 160400 6 la_iena[102]
port 72 nsew signal tristate
rlabel metal2 s 346306 159200 346362 160400 6 la_iena[103]
port 73 nsew signal tristate
rlabel metal2 s 349710 159200 349766 160400 6 la_iena[104]
port 74 nsew signal tristate
rlabel metal2 s 353022 159200 353078 160400 6 la_iena[105]
port 75 nsew signal tristate
rlabel metal2 s 356426 159200 356482 160400 6 la_iena[106]
port 76 nsew signal tristate
rlabel metal2 s 359738 159200 359794 160400 6 la_iena[107]
port 77 nsew signal tristate
rlabel metal2 s 363142 159200 363198 160400 6 la_iena[108]
port 78 nsew signal tristate
rlabel metal2 s 366454 159200 366510 160400 6 la_iena[109]
port 79 nsew signal tristate
rlabel metal2 s 33966 159200 34022 160400 6 la_iena[10]
port 80 nsew signal tristate
rlabel metal2 s 369858 159200 369914 160400 6 la_iena[110]
port 81 nsew signal tristate
rlabel metal2 s 373170 159200 373226 160400 6 la_iena[111]
port 82 nsew signal tristate
rlabel metal2 s 376574 159200 376630 160400 6 la_iena[112]
port 83 nsew signal tristate
rlabel metal2 s 379886 159200 379942 160400 6 la_iena[113]
port 84 nsew signal tristate
rlabel metal2 s 383290 159200 383346 160400 6 la_iena[114]
port 85 nsew signal tristate
rlabel metal2 s 386602 159200 386658 160400 6 la_iena[115]
port 86 nsew signal tristate
rlabel metal2 s 390006 159200 390062 160400 6 la_iena[116]
port 87 nsew signal tristate
rlabel metal2 s 393410 159200 393466 160400 6 la_iena[117]
port 88 nsew signal tristate
rlabel metal2 s 396722 159200 396778 160400 6 la_iena[118]
port 89 nsew signal tristate
rlabel metal2 s 400126 159200 400182 160400 6 la_iena[119]
port 90 nsew signal tristate
rlabel metal2 s 37278 159200 37334 160400 6 la_iena[11]
port 91 nsew signal tristate
rlabel metal2 s 403438 159200 403494 160400 6 la_iena[120]
port 92 nsew signal tristate
rlabel metal2 s 406842 159200 406898 160400 6 la_iena[121]
port 93 nsew signal tristate
rlabel metal2 s 410154 159200 410210 160400 6 la_iena[122]
port 94 nsew signal tristate
rlabel metal2 s 413558 159200 413614 160400 6 la_iena[123]
port 95 nsew signal tristate
rlabel metal2 s 416870 159200 416926 160400 6 la_iena[124]
port 96 nsew signal tristate
rlabel metal2 s 420274 159200 420330 160400 6 la_iena[125]
port 97 nsew signal tristate
rlabel metal2 s 423586 159200 423642 160400 6 la_iena[126]
port 98 nsew signal tristate
rlabel metal2 s 426990 159200 427046 160400 6 la_iena[127]
port 99 nsew signal tristate
rlabel metal2 s 40682 159200 40738 160400 6 la_iena[12]
port 100 nsew signal tristate
rlabel metal2 s 43994 159200 44050 160400 6 la_iena[13]
port 101 nsew signal tristate
rlabel metal2 s 47398 159200 47454 160400 6 la_iena[14]
port 102 nsew signal tristate
rlabel metal2 s 50710 159200 50766 160400 6 la_iena[15]
port 103 nsew signal tristate
rlabel metal2 s 54114 159200 54170 160400 6 la_iena[16]
port 104 nsew signal tristate
rlabel metal2 s 57426 159200 57482 160400 6 la_iena[17]
port 105 nsew signal tristate
rlabel metal2 s 60830 159200 60886 160400 6 la_iena[18]
port 106 nsew signal tristate
rlabel metal2 s 64142 159200 64198 160400 6 la_iena[19]
port 107 nsew signal tristate
rlabel metal2 s 3698 159200 3754 160400 6 la_iena[1]
port 108 nsew signal tristate
rlabel metal2 s 67546 159200 67602 160400 6 la_iena[20]
port 109 nsew signal tristate
rlabel metal2 s 70858 159200 70914 160400 6 la_iena[21]
port 110 nsew signal tristate
rlabel metal2 s 74262 159200 74318 160400 6 la_iena[22]
port 111 nsew signal tristate
rlabel metal2 s 77574 159200 77630 160400 6 la_iena[23]
port 112 nsew signal tristate
rlabel metal2 s 80978 159200 81034 160400 6 la_iena[24]
port 113 nsew signal tristate
rlabel metal2 s 84290 159200 84346 160400 6 la_iena[25]
port 114 nsew signal tristate
rlabel metal2 s 87694 159200 87750 160400 6 la_iena[26]
port 115 nsew signal tristate
rlabel metal2 s 91006 159200 91062 160400 6 la_iena[27]
port 116 nsew signal tristate
rlabel metal2 s 94410 159200 94466 160400 6 la_iena[28]
port 117 nsew signal tristate
rlabel metal2 s 97722 159200 97778 160400 6 la_iena[29]
port 118 nsew signal tristate
rlabel metal2 s 7102 159200 7158 160400 6 la_iena[2]
port 119 nsew signal tristate
rlabel metal2 s 101126 159200 101182 160400 6 la_iena[30]
port 120 nsew signal tristate
rlabel metal2 s 104438 159200 104494 160400 6 la_iena[31]
port 121 nsew signal tristate
rlabel metal2 s 107842 159200 107898 160400 6 la_iena[32]
port 122 nsew signal tristate
rlabel metal2 s 111154 159200 111210 160400 6 la_iena[33]
port 123 nsew signal tristate
rlabel metal2 s 114558 159200 114614 160400 6 la_iena[34]
port 124 nsew signal tristate
rlabel metal2 s 117870 159200 117926 160400 6 la_iena[35]
port 125 nsew signal tristate
rlabel metal2 s 121274 159200 121330 160400 6 la_iena[36]
port 126 nsew signal tristate
rlabel metal2 s 124586 159200 124642 160400 6 la_iena[37]
port 127 nsew signal tristate
rlabel metal2 s 127990 159200 128046 160400 6 la_iena[38]
port 128 nsew signal tristate
rlabel metal2 s 131394 159200 131450 160400 6 la_iena[39]
port 129 nsew signal tristate
rlabel metal2 s 10414 159200 10470 160400 6 la_iena[3]
port 130 nsew signal tristate
rlabel metal2 s 134706 159200 134762 160400 6 la_iena[40]
port 131 nsew signal tristate
rlabel metal2 s 138110 159200 138166 160400 6 la_iena[41]
port 132 nsew signal tristate
rlabel metal2 s 141422 159200 141478 160400 6 la_iena[42]
port 133 nsew signal tristate
rlabel metal2 s 144826 159200 144882 160400 6 la_iena[43]
port 134 nsew signal tristate
rlabel metal2 s 148138 159200 148194 160400 6 la_iena[44]
port 135 nsew signal tristate
rlabel metal2 s 151542 159200 151598 160400 6 la_iena[45]
port 136 nsew signal tristate
rlabel metal2 s 154854 159200 154910 160400 6 la_iena[46]
port 137 nsew signal tristate
rlabel metal2 s 158258 159200 158314 160400 6 la_iena[47]
port 138 nsew signal tristate
rlabel metal2 s 161570 159200 161626 160400 6 la_iena[48]
port 139 nsew signal tristate
rlabel metal2 s 164974 159200 165030 160400 6 la_iena[49]
port 140 nsew signal tristate
rlabel metal2 s 13818 159200 13874 160400 6 la_iena[4]
port 141 nsew signal tristate
rlabel metal2 s 168286 159200 168342 160400 6 la_iena[50]
port 142 nsew signal tristate
rlabel metal2 s 171690 159200 171746 160400 6 la_iena[51]
port 143 nsew signal tristate
rlabel metal2 s 175002 159200 175058 160400 6 la_iena[52]
port 144 nsew signal tristate
rlabel metal2 s 178406 159200 178462 160400 6 la_iena[53]
port 145 nsew signal tristate
rlabel metal2 s 181718 159200 181774 160400 6 la_iena[54]
port 146 nsew signal tristate
rlabel metal2 s 185122 159200 185178 160400 6 la_iena[55]
port 147 nsew signal tristate
rlabel metal2 s 188434 159200 188490 160400 6 la_iena[56]
port 148 nsew signal tristate
rlabel metal2 s 191838 159200 191894 160400 6 la_iena[57]
port 149 nsew signal tristate
rlabel metal2 s 195150 159200 195206 160400 6 la_iena[58]
port 150 nsew signal tristate
rlabel metal2 s 198554 159200 198610 160400 6 la_iena[59]
port 151 nsew signal tristate
rlabel metal2 s 17130 159200 17186 160400 6 la_iena[5]
port 152 nsew signal tristate
rlabel metal2 s 201866 159200 201922 160400 6 la_iena[60]
port 153 nsew signal tristate
rlabel metal2 s 205270 159200 205326 160400 6 la_iena[61]
port 154 nsew signal tristate
rlabel metal2 s 208582 159200 208638 160400 6 la_iena[62]
port 155 nsew signal tristate
rlabel metal2 s 211986 159200 212042 160400 6 la_iena[63]
port 156 nsew signal tristate
rlabel metal2 s 215298 159200 215354 160400 6 la_iena[64]
port 157 nsew signal tristate
rlabel metal2 s 218702 159200 218758 160400 6 la_iena[65]
port 158 nsew signal tristate
rlabel metal2 s 222014 159200 222070 160400 6 la_iena[66]
port 159 nsew signal tristate
rlabel metal2 s 225418 159200 225474 160400 6 la_iena[67]
port 160 nsew signal tristate
rlabel metal2 s 228730 159200 228786 160400 6 la_iena[68]
port 161 nsew signal tristate
rlabel metal2 s 232134 159200 232190 160400 6 la_iena[69]
port 162 nsew signal tristate
rlabel metal2 s 20534 159200 20590 160400 6 la_iena[6]
port 163 nsew signal tristate
rlabel metal2 s 235446 159200 235502 160400 6 la_iena[70]
port 164 nsew signal tristate
rlabel metal2 s 238850 159200 238906 160400 6 la_iena[71]
port 165 nsew signal tristate
rlabel metal2 s 242162 159200 242218 160400 6 la_iena[72]
port 166 nsew signal tristate
rlabel metal2 s 245566 159200 245622 160400 6 la_iena[73]
port 167 nsew signal tristate
rlabel metal2 s 248878 159200 248934 160400 6 la_iena[74]
port 168 nsew signal tristate
rlabel metal2 s 252282 159200 252338 160400 6 la_iena[75]
port 169 nsew signal tristate
rlabel metal2 s 255594 159200 255650 160400 6 la_iena[76]
port 170 nsew signal tristate
rlabel metal2 s 258998 159200 259054 160400 6 la_iena[77]
port 171 nsew signal tristate
rlabel metal2 s 262402 159200 262458 160400 6 la_iena[78]
port 172 nsew signal tristate
rlabel metal2 s 265714 159200 265770 160400 6 la_iena[79]
port 173 nsew signal tristate
rlabel metal2 s 23846 159200 23902 160400 6 la_iena[7]
port 174 nsew signal tristate
rlabel metal2 s 269118 159200 269174 160400 6 la_iena[80]
port 175 nsew signal tristate
rlabel metal2 s 272430 159200 272486 160400 6 la_iena[81]
port 176 nsew signal tristate
rlabel metal2 s 275834 159200 275890 160400 6 la_iena[82]
port 177 nsew signal tristate
rlabel metal2 s 279146 159200 279202 160400 6 la_iena[83]
port 178 nsew signal tristate
rlabel metal2 s 282550 159200 282606 160400 6 la_iena[84]
port 179 nsew signal tristate
rlabel metal2 s 285862 159200 285918 160400 6 la_iena[85]
port 180 nsew signal tristate
rlabel metal2 s 289266 159200 289322 160400 6 la_iena[86]
port 181 nsew signal tristate
rlabel metal2 s 292578 159200 292634 160400 6 la_iena[87]
port 182 nsew signal tristate
rlabel metal2 s 295982 159200 296038 160400 6 la_iena[88]
port 183 nsew signal tristate
rlabel metal2 s 299294 159200 299350 160400 6 la_iena[89]
port 184 nsew signal tristate
rlabel metal2 s 27250 159200 27306 160400 6 la_iena[8]
port 185 nsew signal tristate
rlabel metal2 s 302698 159200 302754 160400 6 la_iena[90]
port 186 nsew signal tristate
rlabel metal2 s 306010 159200 306066 160400 6 la_iena[91]
port 187 nsew signal tristate
rlabel metal2 s 309414 159200 309470 160400 6 la_iena[92]
port 188 nsew signal tristate
rlabel metal2 s 312726 159200 312782 160400 6 la_iena[93]
port 189 nsew signal tristate
rlabel metal2 s 316130 159200 316186 160400 6 la_iena[94]
port 190 nsew signal tristate
rlabel metal2 s 319442 159200 319498 160400 6 la_iena[95]
port 191 nsew signal tristate
rlabel metal2 s 322846 159200 322902 160400 6 la_iena[96]
port 192 nsew signal tristate
rlabel metal2 s 326158 159200 326214 160400 6 la_iena[97]
port 193 nsew signal tristate
rlabel metal2 s 329562 159200 329618 160400 6 la_iena[98]
port 194 nsew signal tristate
rlabel metal2 s 332874 159200 332930 160400 6 la_iena[99]
port 195 nsew signal tristate
rlabel metal2 s 30562 159200 30618 160400 6 la_iena[9]
port 196 nsew signal tristate
rlabel metal2 s 1214 159200 1270 160400 6 la_input[0]
port 197 nsew signal input
rlabel metal2 s 337106 159200 337162 160400 6 la_input[100]
port 198 nsew signal input
rlabel metal2 s 340418 159200 340474 160400 6 la_input[101]
port 199 nsew signal input
rlabel metal2 s 343822 159200 343878 160400 6 la_input[102]
port 200 nsew signal input
rlabel metal2 s 347134 159200 347190 160400 6 la_input[103]
port 201 nsew signal input
rlabel metal2 s 350538 159200 350594 160400 6 la_input[104]
port 202 nsew signal input
rlabel metal2 s 353850 159200 353906 160400 6 la_input[105]
port 203 nsew signal input
rlabel metal2 s 357254 159200 357310 160400 6 la_input[106]
port 204 nsew signal input
rlabel metal2 s 360658 159200 360714 160400 6 la_input[107]
port 205 nsew signal input
rlabel metal2 s 363970 159200 364026 160400 6 la_input[108]
port 206 nsew signal input
rlabel metal2 s 367374 159200 367430 160400 6 la_input[109]
port 207 nsew signal input
rlabel metal2 s 34794 159200 34850 160400 6 la_input[10]
port 208 nsew signal input
rlabel metal2 s 370686 159200 370742 160400 6 la_input[110]
port 209 nsew signal input
rlabel metal2 s 374090 159200 374146 160400 6 la_input[111]
port 210 nsew signal input
rlabel metal2 s 377402 159200 377458 160400 6 la_input[112]
port 211 nsew signal input
rlabel metal2 s 380806 159200 380862 160400 6 la_input[113]
port 212 nsew signal input
rlabel metal2 s 384118 159200 384174 160400 6 la_input[114]
port 213 nsew signal input
rlabel metal2 s 387522 159200 387578 160400 6 la_input[115]
port 214 nsew signal input
rlabel metal2 s 390834 159200 390890 160400 6 la_input[116]
port 215 nsew signal input
rlabel metal2 s 394238 159200 394294 160400 6 la_input[117]
port 216 nsew signal input
rlabel metal2 s 397550 159200 397606 160400 6 la_input[118]
port 217 nsew signal input
rlabel metal2 s 400954 159200 401010 160400 6 la_input[119]
port 218 nsew signal input
rlabel metal2 s 38106 159200 38162 160400 6 la_input[11]
port 219 nsew signal input
rlabel metal2 s 404266 159200 404322 160400 6 la_input[120]
port 220 nsew signal input
rlabel metal2 s 407670 159200 407726 160400 6 la_input[121]
port 221 nsew signal input
rlabel metal2 s 410982 159200 411038 160400 6 la_input[122]
port 222 nsew signal input
rlabel metal2 s 414386 159200 414442 160400 6 la_input[123]
port 223 nsew signal input
rlabel metal2 s 417698 159200 417754 160400 6 la_input[124]
port 224 nsew signal input
rlabel metal2 s 421102 159200 421158 160400 6 la_input[125]
port 225 nsew signal input
rlabel metal2 s 424414 159200 424470 160400 6 la_input[126]
port 226 nsew signal input
rlabel metal2 s 427818 159200 427874 160400 6 la_input[127]
port 227 nsew signal input
rlabel metal2 s 41510 159200 41566 160400 6 la_input[12]
port 228 nsew signal input
rlabel metal2 s 44822 159200 44878 160400 6 la_input[13]
port 229 nsew signal input
rlabel metal2 s 48226 159200 48282 160400 6 la_input[14]
port 230 nsew signal input
rlabel metal2 s 51538 159200 51594 160400 6 la_input[15]
port 231 nsew signal input
rlabel metal2 s 54942 159200 54998 160400 6 la_input[16]
port 232 nsew signal input
rlabel metal2 s 58254 159200 58310 160400 6 la_input[17]
port 233 nsew signal input
rlabel metal2 s 61658 159200 61714 160400 6 la_input[18]
port 234 nsew signal input
rlabel metal2 s 64970 159200 65026 160400 6 la_input[19]
port 235 nsew signal input
rlabel metal2 s 4526 159200 4582 160400 6 la_input[1]
port 236 nsew signal input
rlabel metal2 s 68374 159200 68430 160400 6 la_input[20]
port 237 nsew signal input
rlabel metal2 s 71686 159200 71742 160400 6 la_input[21]
port 238 nsew signal input
rlabel metal2 s 75090 159200 75146 160400 6 la_input[22]
port 239 nsew signal input
rlabel metal2 s 78402 159200 78458 160400 6 la_input[23]
port 240 nsew signal input
rlabel metal2 s 81806 159200 81862 160400 6 la_input[24]
port 241 nsew signal input
rlabel metal2 s 85118 159200 85174 160400 6 la_input[25]
port 242 nsew signal input
rlabel metal2 s 88522 159200 88578 160400 6 la_input[26]
port 243 nsew signal input
rlabel metal2 s 91834 159200 91890 160400 6 la_input[27]
port 244 nsew signal input
rlabel metal2 s 95238 159200 95294 160400 6 la_input[28]
port 245 nsew signal input
rlabel metal2 s 98642 159200 98698 160400 6 la_input[29]
port 246 nsew signal input
rlabel metal2 s 7930 159200 7986 160400 6 la_input[2]
port 247 nsew signal input
rlabel metal2 s 101954 159200 102010 160400 6 la_input[30]
port 248 nsew signal input
rlabel metal2 s 105358 159200 105414 160400 6 la_input[31]
port 249 nsew signal input
rlabel metal2 s 108670 159200 108726 160400 6 la_input[32]
port 250 nsew signal input
rlabel metal2 s 112074 159200 112130 160400 6 la_input[33]
port 251 nsew signal input
rlabel metal2 s 115386 159200 115442 160400 6 la_input[34]
port 252 nsew signal input
rlabel metal2 s 118790 159200 118846 160400 6 la_input[35]
port 253 nsew signal input
rlabel metal2 s 122102 159200 122158 160400 6 la_input[36]
port 254 nsew signal input
rlabel metal2 s 125506 159200 125562 160400 6 la_input[37]
port 255 nsew signal input
rlabel metal2 s 128818 159200 128874 160400 6 la_input[38]
port 256 nsew signal input
rlabel metal2 s 132222 159200 132278 160400 6 la_input[39]
port 257 nsew signal input
rlabel metal2 s 11242 159200 11298 160400 6 la_input[3]
port 258 nsew signal input
rlabel metal2 s 135534 159200 135590 160400 6 la_input[40]
port 259 nsew signal input
rlabel metal2 s 138938 159200 138994 160400 6 la_input[41]
port 260 nsew signal input
rlabel metal2 s 142250 159200 142306 160400 6 la_input[42]
port 261 nsew signal input
rlabel metal2 s 145654 159200 145710 160400 6 la_input[43]
port 262 nsew signal input
rlabel metal2 s 148966 159200 149022 160400 6 la_input[44]
port 263 nsew signal input
rlabel metal2 s 152370 159200 152426 160400 6 la_input[45]
port 264 nsew signal input
rlabel metal2 s 155682 159200 155738 160400 6 la_input[46]
port 265 nsew signal input
rlabel metal2 s 159086 159200 159142 160400 6 la_input[47]
port 266 nsew signal input
rlabel metal2 s 162398 159200 162454 160400 6 la_input[48]
port 267 nsew signal input
rlabel metal2 s 165802 159200 165858 160400 6 la_input[49]
port 268 nsew signal input
rlabel metal2 s 14646 159200 14702 160400 6 la_input[4]
port 269 nsew signal input
rlabel metal2 s 169114 159200 169170 160400 6 la_input[50]
port 270 nsew signal input
rlabel metal2 s 172518 159200 172574 160400 6 la_input[51]
port 271 nsew signal input
rlabel metal2 s 175830 159200 175886 160400 6 la_input[52]
port 272 nsew signal input
rlabel metal2 s 179234 159200 179290 160400 6 la_input[53]
port 273 nsew signal input
rlabel metal2 s 182546 159200 182602 160400 6 la_input[54]
port 274 nsew signal input
rlabel metal2 s 185950 159200 186006 160400 6 la_input[55]
port 275 nsew signal input
rlabel metal2 s 189262 159200 189318 160400 6 la_input[56]
port 276 nsew signal input
rlabel metal2 s 192666 159200 192722 160400 6 la_input[57]
port 277 nsew signal input
rlabel metal2 s 195978 159200 196034 160400 6 la_input[58]
port 278 nsew signal input
rlabel metal2 s 199382 159200 199438 160400 6 la_input[59]
port 279 nsew signal input
rlabel metal2 s 17958 159200 18014 160400 6 la_input[5]
port 280 nsew signal input
rlabel metal2 s 202694 159200 202750 160400 6 la_input[60]
port 281 nsew signal input
rlabel metal2 s 206098 159200 206154 160400 6 la_input[61]
port 282 nsew signal input
rlabel metal2 s 209410 159200 209466 160400 6 la_input[62]
port 283 nsew signal input
rlabel metal2 s 212814 159200 212870 160400 6 la_input[63]
port 284 nsew signal input
rlabel metal2 s 216126 159200 216182 160400 6 la_input[64]
port 285 nsew signal input
rlabel metal2 s 219530 159200 219586 160400 6 la_input[65]
port 286 nsew signal input
rlabel metal2 s 222842 159200 222898 160400 6 la_input[66]
port 287 nsew signal input
rlabel metal2 s 226246 159200 226302 160400 6 la_input[67]
port 288 nsew signal input
rlabel metal2 s 229650 159200 229706 160400 6 la_input[68]
port 289 nsew signal input
rlabel metal2 s 232962 159200 233018 160400 6 la_input[69]
port 290 nsew signal input
rlabel metal2 s 21362 159200 21418 160400 6 la_input[6]
port 291 nsew signal input
rlabel metal2 s 236366 159200 236422 160400 6 la_input[70]
port 292 nsew signal input
rlabel metal2 s 239678 159200 239734 160400 6 la_input[71]
port 293 nsew signal input
rlabel metal2 s 243082 159200 243138 160400 6 la_input[72]
port 294 nsew signal input
rlabel metal2 s 246394 159200 246450 160400 6 la_input[73]
port 295 nsew signal input
rlabel metal2 s 249798 159200 249854 160400 6 la_input[74]
port 296 nsew signal input
rlabel metal2 s 253110 159200 253166 160400 6 la_input[75]
port 297 nsew signal input
rlabel metal2 s 256514 159200 256570 160400 6 la_input[76]
port 298 nsew signal input
rlabel metal2 s 259826 159200 259882 160400 6 la_input[77]
port 299 nsew signal input
rlabel metal2 s 263230 159200 263286 160400 6 la_input[78]
port 300 nsew signal input
rlabel metal2 s 266542 159200 266598 160400 6 la_input[79]
port 301 nsew signal input
rlabel metal2 s 24674 159200 24730 160400 6 la_input[7]
port 302 nsew signal input
rlabel metal2 s 269946 159200 270002 160400 6 la_input[80]
port 303 nsew signal input
rlabel metal2 s 273258 159200 273314 160400 6 la_input[81]
port 304 nsew signal input
rlabel metal2 s 276662 159200 276718 160400 6 la_input[82]
port 305 nsew signal input
rlabel metal2 s 279974 159200 280030 160400 6 la_input[83]
port 306 nsew signal input
rlabel metal2 s 283378 159200 283434 160400 6 la_input[84]
port 307 nsew signal input
rlabel metal2 s 286690 159200 286746 160400 6 la_input[85]
port 308 nsew signal input
rlabel metal2 s 290094 159200 290150 160400 6 la_input[86]
port 309 nsew signal input
rlabel metal2 s 293406 159200 293462 160400 6 la_input[87]
port 310 nsew signal input
rlabel metal2 s 296810 159200 296866 160400 6 la_input[88]
port 311 nsew signal input
rlabel metal2 s 300122 159200 300178 160400 6 la_input[89]
port 312 nsew signal input
rlabel metal2 s 28078 159200 28134 160400 6 la_input[8]
port 313 nsew signal input
rlabel metal2 s 303526 159200 303582 160400 6 la_input[90]
port 314 nsew signal input
rlabel metal2 s 306838 159200 306894 160400 6 la_input[91]
port 315 nsew signal input
rlabel metal2 s 310242 159200 310298 160400 6 la_input[92]
port 316 nsew signal input
rlabel metal2 s 313554 159200 313610 160400 6 la_input[93]
port 317 nsew signal input
rlabel metal2 s 316958 159200 317014 160400 6 la_input[94]
port 318 nsew signal input
rlabel metal2 s 320270 159200 320326 160400 6 la_input[95]
port 319 nsew signal input
rlabel metal2 s 323674 159200 323730 160400 6 la_input[96]
port 320 nsew signal input
rlabel metal2 s 326986 159200 327042 160400 6 la_input[97]
port 321 nsew signal input
rlabel metal2 s 330390 159200 330446 160400 6 la_input[98]
port 322 nsew signal input
rlabel metal2 s 333702 159200 333758 160400 6 la_input[99]
port 323 nsew signal input
rlabel metal2 s 31390 159200 31446 160400 6 la_input[9]
port 324 nsew signal input
rlabel metal2 s 2042 159200 2098 160400 6 la_oenb[0]
port 325 nsew signal tristate
rlabel metal2 s 337934 159200 337990 160400 6 la_oenb[100]
port 326 nsew signal tristate
rlabel metal2 s 341338 159200 341394 160400 6 la_oenb[101]
port 327 nsew signal tristate
rlabel metal2 s 344650 159200 344706 160400 6 la_oenb[102]
port 328 nsew signal tristate
rlabel metal2 s 348054 159200 348110 160400 6 la_oenb[103]
port 329 nsew signal tristate
rlabel metal2 s 351366 159200 351422 160400 6 la_oenb[104]
port 330 nsew signal tristate
rlabel metal2 s 354770 159200 354826 160400 6 la_oenb[105]
port 331 nsew signal tristate
rlabel metal2 s 358082 159200 358138 160400 6 la_oenb[106]
port 332 nsew signal tristate
rlabel metal2 s 361486 159200 361542 160400 6 la_oenb[107]
port 333 nsew signal tristate
rlabel metal2 s 364798 159200 364854 160400 6 la_oenb[108]
port 334 nsew signal tristate
rlabel metal2 s 368202 159200 368258 160400 6 la_oenb[109]
port 335 nsew signal tristate
rlabel metal2 s 35622 159200 35678 160400 6 la_oenb[10]
port 336 nsew signal tristate
rlabel metal2 s 371514 159200 371570 160400 6 la_oenb[110]
port 337 nsew signal tristate
rlabel metal2 s 374918 159200 374974 160400 6 la_oenb[111]
port 338 nsew signal tristate
rlabel metal2 s 378230 159200 378286 160400 6 la_oenb[112]
port 339 nsew signal tristate
rlabel metal2 s 381634 159200 381690 160400 6 la_oenb[113]
port 340 nsew signal tristate
rlabel metal2 s 384946 159200 385002 160400 6 la_oenb[114]
port 341 nsew signal tristate
rlabel metal2 s 388350 159200 388406 160400 6 la_oenb[115]
port 342 nsew signal tristate
rlabel metal2 s 391662 159200 391718 160400 6 la_oenb[116]
port 343 nsew signal tristate
rlabel metal2 s 395066 159200 395122 160400 6 la_oenb[117]
port 344 nsew signal tristate
rlabel metal2 s 398378 159200 398434 160400 6 la_oenb[118]
port 345 nsew signal tristate
rlabel metal2 s 401782 159200 401838 160400 6 la_oenb[119]
port 346 nsew signal tristate
rlabel metal2 s 38934 159200 38990 160400 6 la_oenb[11]
port 347 nsew signal tristate
rlabel metal2 s 405094 159200 405150 160400 6 la_oenb[120]
port 348 nsew signal tristate
rlabel metal2 s 408498 159200 408554 160400 6 la_oenb[121]
port 349 nsew signal tristate
rlabel metal2 s 411810 159200 411866 160400 6 la_oenb[122]
port 350 nsew signal tristate
rlabel metal2 s 415214 159200 415270 160400 6 la_oenb[123]
port 351 nsew signal tristate
rlabel metal2 s 418526 159200 418582 160400 6 la_oenb[124]
port 352 nsew signal tristate
rlabel metal2 s 421930 159200 421986 160400 6 la_oenb[125]
port 353 nsew signal tristate
rlabel metal2 s 425242 159200 425298 160400 6 la_oenb[126]
port 354 nsew signal tristate
rlabel metal2 s 428646 159200 428702 160400 6 la_oenb[127]
port 355 nsew signal tristate
rlabel metal2 s 42338 159200 42394 160400 6 la_oenb[12]
port 356 nsew signal tristate
rlabel metal2 s 45650 159200 45706 160400 6 la_oenb[13]
port 357 nsew signal tristate
rlabel metal2 s 49054 159200 49110 160400 6 la_oenb[14]
port 358 nsew signal tristate
rlabel metal2 s 52366 159200 52422 160400 6 la_oenb[15]
port 359 nsew signal tristate
rlabel metal2 s 55770 159200 55826 160400 6 la_oenb[16]
port 360 nsew signal tristate
rlabel metal2 s 59082 159200 59138 160400 6 la_oenb[17]
port 361 nsew signal tristate
rlabel metal2 s 62486 159200 62542 160400 6 la_oenb[18]
port 362 nsew signal tristate
rlabel metal2 s 65890 159200 65946 160400 6 la_oenb[19]
port 363 nsew signal tristate
rlabel metal2 s 5354 159200 5410 160400 6 la_oenb[1]
port 364 nsew signal tristate
rlabel metal2 s 69202 159200 69258 160400 6 la_oenb[20]
port 365 nsew signal tristate
rlabel metal2 s 72606 159200 72662 160400 6 la_oenb[21]
port 366 nsew signal tristate
rlabel metal2 s 75918 159200 75974 160400 6 la_oenb[22]
port 367 nsew signal tristate
rlabel metal2 s 79322 159200 79378 160400 6 la_oenb[23]
port 368 nsew signal tristate
rlabel metal2 s 82634 159200 82690 160400 6 la_oenb[24]
port 369 nsew signal tristate
rlabel metal2 s 86038 159200 86094 160400 6 la_oenb[25]
port 370 nsew signal tristate
rlabel metal2 s 89350 159200 89406 160400 6 la_oenb[26]
port 371 nsew signal tristate
rlabel metal2 s 92754 159200 92810 160400 6 la_oenb[27]
port 372 nsew signal tristate
rlabel metal2 s 96066 159200 96122 160400 6 la_oenb[28]
port 373 nsew signal tristate
rlabel metal2 s 99470 159200 99526 160400 6 la_oenb[29]
port 374 nsew signal tristate
rlabel metal2 s 8758 159200 8814 160400 6 la_oenb[2]
port 375 nsew signal tristate
rlabel metal2 s 102782 159200 102838 160400 6 la_oenb[30]
port 376 nsew signal tristate
rlabel metal2 s 106186 159200 106242 160400 6 la_oenb[31]
port 377 nsew signal tristate
rlabel metal2 s 109498 159200 109554 160400 6 la_oenb[32]
port 378 nsew signal tristate
rlabel metal2 s 112902 159200 112958 160400 6 la_oenb[33]
port 379 nsew signal tristate
rlabel metal2 s 116214 159200 116270 160400 6 la_oenb[34]
port 380 nsew signal tristate
rlabel metal2 s 119618 159200 119674 160400 6 la_oenb[35]
port 381 nsew signal tristate
rlabel metal2 s 122930 159200 122986 160400 6 la_oenb[36]
port 382 nsew signal tristate
rlabel metal2 s 126334 159200 126390 160400 6 la_oenb[37]
port 383 nsew signal tristate
rlabel metal2 s 129646 159200 129702 160400 6 la_oenb[38]
port 384 nsew signal tristate
rlabel metal2 s 133050 159200 133106 160400 6 la_oenb[39]
port 385 nsew signal tristate
rlabel metal2 s 12070 159200 12126 160400 6 la_oenb[3]
port 386 nsew signal tristate
rlabel metal2 s 136362 159200 136418 160400 6 la_oenb[40]
port 387 nsew signal tristate
rlabel metal2 s 139766 159200 139822 160400 6 la_oenb[41]
port 388 nsew signal tristate
rlabel metal2 s 143078 159200 143134 160400 6 la_oenb[42]
port 389 nsew signal tristate
rlabel metal2 s 146482 159200 146538 160400 6 la_oenb[43]
port 390 nsew signal tristate
rlabel metal2 s 149794 159200 149850 160400 6 la_oenb[44]
port 391 nsew signal tristate
rlabel metal2 s 153198 159200 153254 160400 6 la_oenb[45]
port 392 nsew signal tristate
rlabel metal2 s 156510 159200 156566 160400 6 la_oenb[46]
port 393 nsew signal tristate
rlabel metal2 s 159914 159200 159970 160400 6 la_oenb[47]
port 394 nsew signal tristate
rlabel metal2 s 163226 159200 163282 160400 6 la_oenb[48]
port 395 nsew signal tristate
rlabel metal2 s 166630 159200 166686 160400 6 la_oenb[49]
port 396 nsew signal tristate
rlabel metal2 s 15474 159200 15530 160400 6 la_oenb[4]
port 397 nsew signal tristate
rlabel metal2 s 169942 159200 169998 160400 6 la_oenb[50]
port 398 nsew signal tristate
rlabel metal2 s 173346 159200 173402 160400 6 la_oenb[51]
port 399 nsew signal tristate
rlabel metal2 s 176658 159200 176714 160400 6 la_oenb[52]
port 400 nsew signal tristate
rlabel metal2 s 180062 159200 180118 160400 6 la_oenb[53]
port 401 nsew signal tristate
rlabel metal2 s 183374 159200 183430 160400 6 la_oenb[54]
port 402 nsew signal tristate
rlabel metal2 s 186778 159200 186834 160400 6 la_oenb[55]
port 403 nsew signal tristate
rlabel metal2 s 190090 159200 190146 160400 6 la_oenb[56]
port 404 nsew signal tristate
rlabel metal2 s 193494 159200 193550 160400 6 la_oenb[57]
port 405 nsew signal tristate
rlabel metal2 s 196898 159200 196954 160400 6 la_oenb[58]
port 406 nsew signal tristate
rlabel metal2 s 200210 159200 200266 160400 6 la_oenb[59]
port 407 nsew signal tristate
rlabel metal2 s 18786 159200 18842 160400 6 la_oenb[5]
port 408 nsew signal tristate
rlabel metal2 s 203614 159200 203670 160400 6 la_oenb[60]
port 409 nsew signal tristate
rlabel metal2 s 206926 159200 206982 160400 6 la_oenb[61]
port 410 nsew signal tristate
rlabel metal2 s 210330 159200 210386 160400 6 la_oenb[62]
port 411 nsew signal tristate
rlabel metal2 s 213642 159200 213698 160400 6 la_oenb[63]
port 412 nsew signal tristate
rlabel metal2 s 217046 159200 217102 160400 6 la_oenb[64]
port 413 nsew signal tristate
rlabel metal2 s 220358 159200 220414 160400 6 la_oenb[65]
port 414 nsew signal tristate
rlabel metal2 s 223762 159200 223818 160400 6 la_oenb[66]
port 415 nsew signal tristate
rlabel metal2 s 227074 159200 227130 160400 6 la_oenb[67]
port 416 nsew signal tristate
rlabel metal2 s 230478 159200 230534 160400 6 la_oenb[68]
port 417 nsew signal tristate
rlabel metal2 s 233790 159200 233846 160400 6 la_oenb[69]
port 418 nsew signal tristate
rlabel metal2 s 22190 159200 22246 160400 6 la_oenb[6]
port 419 nsew signal tristate
rlabel metal2 s 237194 159200 237250 160400 6 la_oenb[70]
port 420 nsew signal tristate
rlabel metal2 s 240506 159200 240562 160400 6 la_oenb[71]
port 421 nsew signal tristate
rlabel metal2 s 243910 159200 243966 160400 6 la_oenb[72]
port 422 nsew signal tristate
rlabel metal2 s 247222 159200 247278 160400 6 la_oenb[73]
port 423 nsew signal tristate
rlabel metal2 s 250626 159200 250682 160400 6 la_oenb[74]
port 424 nsew signal tristate
rlabel metal2 s 253938 159200 253994 160400 6 la_oenb[75]
port 425 nsew signal tristate
rlabel metal2 s 257342 159200 257398 160400 6 la_oenb[76]
port 426 nsew signal tristate
rlabel metal2 s 260654 159200 260710 160400 6 la_oenb[77]
port 427 nsew signal tristate
rlabel metal2 s 264058 159200 264114 160400 6 la_oenb[78]
port 428 nsew signal tristate
rlabel metal2 s 267370 159200 267426 160400 6 la_oenb[79]
port 429 nsew signal tristate
rlabel metal2 s 25502 159200 25558 160400 6 la_oenb[7]
port 430 nsew signal tristate
rlabel metal2 s 270774 159200 270830 160400 6 la_oenb[80]
port 431 nsew signal tristate
rlabel metal2 s 274086 159200 274142 160400 6 la_oenb[81]
port 432 nsew signal tristate
rlabel metal2 s 277490 159200 277546 160400 6 la_oenb[82]
port 433 nsew signal tristate
rlabel metal2 s 280802 159200 280858 160400 6 la_oenb[83]
port 434 nsew signal tristate
rlabel metal2 s 284206 159200 284262 160400 6 la_oenb[84]
port 435 nsew signal tristate
rlabel metal2 s 287518 159200 287574 160400 6 la_oenb[85]
port 436 nsew signal tristate
rlabel metal2 s 290922 159200 290978 160400 6 la_oenb[86]
port 437 nsew signal tristate
rlabel metal2 s 294234 159200 294290 160400 6 la_oenb[87]
port 438 nsew signal tristate
rlabel metal2 s 297638 159200 297694 160400 6 la_oenb[88]
port 439 nsew signal tristate
rlabel metal2 s 300950 159200 301006 160400 6 la_oenb[89]
port 440 nsew signal tristate
rlabel metal2 s 28906 159200 28962 160400 6 la_oenb[8]
port 441 nsew signal tristate
rlabel metal2 s 304354 159200 304410 160400 6 la_oenb[90]
port 442 nsew signal tristate
rlabel metal2 s 307666 159200 307722 160400 6 la_oenb[91]
port 443 nsew signal tristate
rlabel metal2 s 311070 159200 311126 160400 6 la_oenb[92]
port 444 nsew signal tristate
rlabel metal2 s 314382 159200 314438 160400 6 la_oenb[93]
port 445 nsew signal tristate
rlabel metal2 s 317786 159200 317842 160400 6 la_oenb[94]
port 446 nsew signal tristate
rlabel metal2 s 321098 159200 321154 160400 6 la_oenb[95]
port 447 nsew signal tristate
rlabel metal2 s 324502 159200 324558 160400 6 la_oenb[96]
port 448 nsew signal tristate
rlabel metal2 s 327906 159200 327962 160400 6 la_oenb[97]
port 449 nsew signal tristate
rlabel metal2 s 331218 159200 331274 160400 6 la_oenb[98]
port 450 nsew signal tristate
rlabel metal2 s 334622 159200 334678 160400 6 la_oenb[99]
port 451 nsew signal tristate
rlabel metal2 s 32218 159200 32274 160400 6 la_oenb[9]
port 452 nsew signal tristate
rlabel metal2 s 2870 159200 2926 160400 6 la_output[0]
port 453 nsew signal tristate
rlabel metal2 s 338762 159200 338818 160400 6 la_output[100]
port 454 nsew signal tristate
rlabel metal2 s 342166 159200 342222 160400 6 la_output[101]
port 455 nsew signal tristate
rlabel metal2 s 345478 159200 345534 160400 6 la_output[102]
port 456 nsew signal tristate
rlabel metal2 s 348882 159200 348938 160400 6 la_output[103]
port 457 nsew signal tristate
rlabel metal2 s 352194 159200 352250 160400 6 la_output[104]
port 458 nsew signal tristate
rlabel metal2 s 355598 159200 355654 160400 6 la_output[105]
port 459 nsew signal tristate
rlabel metal2 s 358910 159200 358966 160400 6 la_output[106]
port 460 nsew signal tristate
rlabel metal2 s 362314 159200 362370 160400 6 la_output[107]
port 461 nsew signal tristate
rlabel metal2 s 365626 159200 365682 160400 6 la_output[108]
port 462 nsew signal tristate
rlabel metal2 s 369030 159200 369086 160400 6 la_output[109]
port 463 nsew signal tristate
rlabel metal2 s 36450 159200 36506 160400 6 la_output[10]
port 464 nsew signal tristate
rlabel metal2 s 372342 159200 372398 160400 6 la_output[110]
port 465 nsew signal tristate
rlabel metal2 s 375746 159200 375802 160400 6 la_output[111]
port 466 nsew signal tristate
rlabel metal2 s 379058 159200 379114 160400 6 la_output[112]
port 467 nsew signal tristate
rlabel metal2 s 382462 159200 382518 160400 6 la_output[113]
port 468 nsew signal tristate
rlabel metal2 s 385774 159200 385830 160400 6 la_output[114]
port 469 nsew signal tristate
rlabel metal2 s 389178 159200 389234 160400 6 la_output[115]
port 470 nsew signal tristate
rlabel metal2 s 392490 159200 392546 160400 6 la_output[116]
port 471 nsew signal tristate
rlabel metal2 s 395894 159200 395950 160400 6 la_output[117]
port 472 nsew signal tristate
rlabel metal2 s 399206 159200 399262 160400 6 la_output[118]
port 473 nsew signal tristate
rlabel metal2 s 402610 159200 402666 160400 6 la_output[119]
port 474 nsew signal tristate
rlabel metal2 s 39854 159200 39910 160400 6 la_output[11]
port 475 nsew signal tristate
rlabel metal2 s 405922 159200 405978 160400 6 la_output[120]
port 476 nsew signal tristate
rlabel metal2 s 409326 159200 409382 160400 6 la_output[121]
port 477 nsew signal tristate
rlabel metal2 s 412638 159200 412694 160400 6 la_output[122]
port 478 nsew signal tristate
rlabel metal2 s 416042 159200 416098 160400 6 la_output[123]
port 479 nsew signal tristate
rlabel metal2 s 419354 159200 419410 160400 6 la_output[124]
port 480 nsew signal tristate
rlabel metal2 s 422758 159200 422814 160400 6 la_output[125]
port 481 nsew signal tristate
rlabel metal2 s 426162 159200 426218 160400 6 la_output[126]
port 482 nsew signal tristate
rlabel metal2 s 429474 159200 429530 160400 6 la_output[127]
port 483 nsew signal tristate
rlabel metal2 s 43166 159200 43222 160400 6 la_output[12]
port 484 nsew signal tristate
rlabel metal2 s 46570 159200 46626 160400 6 la_output[13]
port 485 nsew signal tristate
rlabel metal2 s 49882 159200 49938 160400 6 la_output[14]
port 486 nsew signal tristate
rlabel metal2 s 53286 159200 53342 160400 6 la_output[15]
port 487 nsew signal tristate
rlabel metal2 s 56598 159200 56654 160400 6 la_output[16]
port 488 nsew signal tristate
rlabel metal2 s 60002 159200 60058 160400 6 la_output[17]
port 489 nsew signal tristate
rlabel metal2 s 63314 159200 63370 160400 6 la_output[18]
port 490 nsew signal tristate
rlabel metal2 s 66718 159200 66774 160400 6 la_output[19]
port 491 nsew signal tristate
rlabel metal2 s 6182 159200 6238 160400 6 la_output[1]
port 492 nsew signal tristate
rlabel metal2 s 70030 159200 70086 160400 6 la_output[20]
port 493 nsew signal tristate
rlabel metal2 s 73434 159200 73490 160400 6 la_output[21]
port 494 nsew signal tristate
rlabel metal2 s 76746 159200 76802 160400 6 la_output[22]
port 495 nsew signal tristate
rlabel metal2 s 80150 159200 80206 160400 6 la_output[23]
port 496 nsew signal tristate
rlabel metal2 s 83462 159200 83518 160400 6 la_output[24]
port 497 nsew signal tristate
rlabel metal2 s 86866 159200 86922 160400 6 la_output[25]
port 498 nsew signal tristate
rlabel metal2 s 90178 159200 90234 160400 6 la_output[26]
port 499 nsew signal tristate
rlabel metal2 s 93582 159200 93638 160400 6 la_output[27]
port 500 nsew signal tristate
rlabel metal2 s 96894 159200 96950 160400 6 la_output[28]
port 501 nsew signal tristate
rlabel metal2 s 100298 159200 100354 160400 6 la_output[29]
port 502 nsew signal tristate
rlabel metal2 s 9586 159200 9642 160400 6 la_output[2]
port 503 nsew signal tristate
rlabel metal2 s 103610 159200 103666 160400 6 la_output[30]
port 504 nsew signal tristate
rlabel metal2 s 107014 159200 107070 160400 6 la_output[31]
port 505 nsew signal tristate
rlabel metal2 s 110326 159200 110382 160400 6 la_output[32]
port 506 nsew signal tristate
rlabel metal2 s 113730 159200 113786 160400 6 la_output[33]
port 507 nsew signal tristate
rlabel metal2 s 117042 159200 117098 160400 6 la_output[34]
port 508 nsew signal tristate
rlabel metal2 s 120446 159200 120502 160400 6 la_output[35]
port 509 nsew signal tristate
rlabel metal2 s 123758 159200 123814 160400 6 la_output[36]
port 510 nsew signal tristate
rlabel metal2 s 127162 159200 127218 160400 6 la_output[37]
port 511 nsew signal tristate
rlabel metal2 s 130474 159200 130530 160400 6 la_output[38]
port 512 nsew signal tristate
rlabel metal2 s 133878 159200 133934 160400 6 la_output[39]
port 513 nsew signal tristate
rlabel metal2 s 12898 159200 12954 160400 6 la_output[3]
port 514 nsew signal tristate
rlabel metal2 s 137190 159200 137246 160400 6 la_output[40]
port 515 nsew signal tristate
rlabel metal2 s 140594 159200 140650 160400 6 la_output[41]
port 516 nsew signal tristate
rlabel metal2 s 143906 159200 143962 160400 6 la_output[42]
port 517 nsew signal tristate
rlabel metal2 s 147310 159200 147366 160400 6 la_output[43]
port 518 nsew signal tristate
rlabel metal2 s 150622 159200 150678 160400 6 la_output[44]
port 519 nsew signal tristate
rlabel metal2 s 154026 159200 154082 160400 6 la_output[45]
port 520 nsew signal tristate
rlabel metal2 s 157338 159200 157394 160400 6 la_output[46]
port 521 nsew signal tristate
rlabel metal2 s 160742 159200 160798 160400 6 la_output[47]
port 522 nsew signal tristate
rlabel metal2 s 164146 159200 164202 160400 6 la_output[48]
port 523 nsew signal tristate
rlabel metal2 s 167458 159200 167514 160400 6 la_output[49]
port 524 nsew signal tristate
rlabel metal2 s 16302 159200 16358 160400 6 la_output[4]
port 525 nsew signal tristate
rlabel metal2 s 170862 159200 170918 160400 6 la_output[50]
port 526 nsew signal tristate
rlabel metal2 s 174174 159200 174230 160400 6 la_output[51]
port 527 nsew signal tristate
rlabel metal2 s 177578 159200 177634 160400 6 la_output[52]
port 528 nsew signal tristate
rlabel metal2 s 180890 159200 180946 160400 6 la_output[53]
port 529 nsew signal tristate
rlabel metal2 s 184294 159200 184350 160400 6 la_output[54]
port 530 nsew signal tristate
rlabel metal2 s 187606 159200 187662 160400 6 la_output[55]
port 531 nsew signal tristate
rlabel metal2 s 191010 159200 191066 160400 6 la_output[56]
port 532 nsew signal tristate
rlabel metal2 s 194322 159200 194378 160400 6 la_output[57]
port 533 nsew signal tristate
rlabel metal2 s 197726 159200 197782 160400 6 la_output[58]
port 534 nsew signal tristate
rlabel metal2 s 201038 159200 201094 160400 6 la_output[59]
port 535 nsew signal tristate
rlabel metal2 s 19614 159200 19670 160400 6 la_output[5]
port 536 nsew signal tristate
rlabel metal2 s 204442 159200 204498 160400 6 la_output[60]
port 537 nsew signal tristate
rlabel metal2 s 207754 159200 207810 160400 6 la_output[61]
port 538 nsew signal tristate
rlabel metal2 s 211158 159200 211214 160400 6 la_output[62]
port 539 nsew signal tristate
rlabel metal2 s 214470 159200 214526 160400 6 la_output[63]
port 540 nsew signal tristate
rlabel metal2 s 217874 159200 217930 160400 6 la_output[64]
port 541 nsew signal tristate
rlabel metal2 s 221186 159200 221242 160400 6 la_output[65]
port 542 nsew signal tristate
rlabel metal2 s 224590 159200 224646 160400 6 la_output[66]
port 543 nsew signal tristate
rlabel metal2 s 227902 159200 227958 160400 6 la_output[67]
port 544 nsew signal tristate
rlabel metal2 s 231306 159200 231362 160400 6 la_output[68]
port 545 nsew signal tristate
rlabel metal2 s 234618 159200 234674 160400 6 la_output[69]
port 546 nsew signal tristate
rlabel metal2 s 23018 159200 23074 160400 6 la_output[6]
port 547 nsew signal tristate
rlabel metal2 s 238022 159200 238078 160400 6 la_output[70]
port 548 nsew signal tristate
rlabel metal2 s 241334 159200 241390 160400 6 la_output[71]
port 549 nsew signal tristate
rlabel metal2 s 244738 159200 244794 160400 6 la_output[72]
port 550 nsew signal tristate
rlabel metal2 s 248050 159200 248106 160400 6 la_output[73]
port 551 nsew signal tristate
rlabel metal2 s 251454 159200 251510 160400 6 la_output[74]
port 552 nsew signal tristate
rlabel metal2 s 254766 159200 254822 160400 6 la_output[75]
port 553 nsew signal tristate
rlabel metal2 s 258170 159200 258226 160400 6 la_output[76]
port 554 nsew signal tristate
rlabel metal2 s 261482 159200 261538 160400 6 la_output[77]
port 555 nsew signal tristate
rlabel metal2 s 264886 159200 264942 160400 6 la_output[78]
port 556 nsew signal tristate
rlabel metal2 s 268198 159200 268254 160400 6 la_output[79]
port 557 nsew signal tristate
rlabel metal2 s 26330 159200 26386 160400 6 la_output[7]
port 558 nsew signal tristate
rlabel metal2 s 271602 159200 271658 160400 6 la_output[80]
port 559 nsew signal tristate
rlabel metal2 s 274914 159200 274970 160400 6 la_output[81]
port 560 nsew signal tristate
rlabel metal2 s 278318 159200 278374 160400 6 la_output[82]
port 561 nsew signal tristate
rlabel metal2 s 281630 159200 281686 160400 6 la_output[83]
port 562 nsew signal tristate
rlabel metal2 s 285034 159200 285090 160400 6 la_output[84]
port 563 nsew signal tristate
rlabel metal2 s 288346 159200 288402 160400 6 la_output[85]
port 564 nsew signal tristate
rlabel metal2 s 291750 159200 291806 160400 6 la_output[86]
port 565 nsew signal tristate
rlabel metal2 s 295154 159200 295210 160400 6 la_output[87]
port 566 nsew signal tristate
rlabel metal2 s 298466 159200 298522 160400 6 la_output[88]
port 567 nsew signal tristate
rlabel metal2 s 301870 159200 301926 160400 6 la_output[89]
port 568 nsew signal tristate
rlabel metal2 s 29734 159200 29790 160400 6 la_output[8]
port 569 nsew signal tristate
rlabel metal2 s 305182 159200 305238 160400 6 la_output[90]
port 570 nsew signal tristate
rlabel metal2 s 308586 159200 308642 160400 6 la_output[91]
port 571 nsew signal tristate
rlabel metal2 s 311898 159200 311954 160400 6 la_output[92]
port 572 nsew signal tristate
rlabel metal2 s 315302 159200 315358 160400 6 la_output[93]
port 573 nsew signal tristate
rlabel metal2 s 318614 159200 318670 160400 6 la_output[94]
port 574 nsew signal tristate
rlabel metal2 s 322018 159200 322074 160400 6 la_output[95]
port 575 nsew signal tristate
rlabel metal2 s 325330 159200 325386 160400 6 la_output[96]
port 576 nsew signal tristate
rlabel metal2 s 328734 159200 328790 160400 6 la_output[97]
port 577 nsew signal tristate
rlabel metal2 s 332046 159200 332102 160400 6 la_output[98]
port 578 nsew signal tristate
rlabel metal2 s 335450 159200 335506 160400 6 la_output[99]
port 579 nsew signal tristate
rlabel metal2 s 33138 159200 33194 160400 6 la_output[9]
port 580 nsew signal tristate
rlabel metal2 s 430302 159200 430358 160400 6 mprj_ack_i
port 581 nsew signal input
rlabel metal2 s 434534 159200 434590 160400 6 mprj_adr_o[0]
port 582 nsew signal tristate
rlabel metal2 s 463054 159200 463110 160400 6 mprj_adr_o[10]
port 583 nsew signal tristate
rlabel metal2 s 465630 159200 465686 160400 6 mprj_adr_o[11]
port 584 nsew signal tristate
rlabel metal2 s 468114 159200 468170 160400 6 mprj_adr_o[12]
port 585 nsew signal tristate
rlabel metal2 s 470598 159200 470654 160400 6 mprj_adr_o[13]
port 586 nsew signal tristate
rlabel metal2 s 473174 159200 473230 160400 6 mprj_adr_o[14]
port 587 nsew signal tristate
rlabel metal2 s 475658 159200 475714 160400 6 mprj_adr_o[15]
port 588 nsew signal tristate
rlabel metal2 s 478142 159200 478198 160400 6 mprj_adr_o[16]
port 589 nsew signal tristate
rlabel metal2 s 480718 159200 480774 160400 6 mprj_adr_o[17]
port 590 nsew signal tristate
rlabel metal2 s 483202 159200 483258 160400 6 mprj_adr_o[18]
port 591 nsew signal tristate
rlabel metal2 s 485778 159200 485834 160400 6 mprj_adr_o[19]
port 592 nsew signal tristate
rlabel metal2 s 437846 159200 437902 160400 6 mprj_adr_o[1]
port 593 nsew signal tristate
rlabel metal2 s 488262 159200 488318 160400 6 mprj_adr_o[20]
port 594 nsew signal tristate
rlabel metal2 s 490746 159200 490802 160400 6 mprj_adr_o[21]
port 595 nsew signal tristate
rlabel metal2 s 493322 159200 493378 160400 6 mprj_adr_o[22]
port 596 nsew signal tristate
rlabel metal2 s 495806 159200 495862 160400 6 mprj_adr_o[23]
port 597 nsew signal tristate
rlabel metal2 s 498382 159200 498438 160400 6 mprj_adr_o[24]
port 598 nsew signal tristate
rlabel metal2 s 500866 159200 500922 160400 6 mprj_adr_o[25]
port 599 nsew signal tristate
rlabel metal2 s 503350 159200 503406 160400 6 mprj_adr_o[26]
port 600 nsew signal tristate
rlabel metal2 s 505926 159200 505982 160400 6 mprj_adr_o[27]
port 601 nsew signal tristate
rlabel metal2 s 508410 159200 508466 160400 6 mprj_adr_o[28]
port 602 nsew signal tristate
rlabel metal2 s 510894 159200 510950 160400 6 mprj_adr_o[29]
port 603 nsew signal tristate
rlabel metal2 s 441250 159200 441306 160400 6 mprj_adr_o[2]
port 604 nsew signal tristate
rlabel metal2 s 513470 159200 513526 160400 6 mprj_adr_o[30]
port 605 nsew signal tristate
rlabel metal2 s 515954 159200 516010 160400 6 mprj_adr_o[31]
port 606 nsew signal tristate
rlabel metal2 s 444562 159200 444618 160400 6 mprj_adr_o[3]
port 607 nsew signal tristate
rlabel metal2 s 447966 159200 448022 160400 6 mprj_adr_o[4]
port 608 nsew signal tristate
rlabel metal2 s 450450 159200 450506 160400 6 mprj_adr_o[5]
port 609 nsew signal tristate
rlabel metal2 s 453026 159200 453082 160400 6 mprj_adr_o[6]
port 610 nsew signal tristate
rlabel metal2 s 455510 159200 455566 160400 6 mprj_adr_o[7]
port 611 nsew signal tristate
rlabel metal2 s 457994 159200 458050 160400 6 mprj_adr_o[8]
port 612 nsew signal tristate
rlabel metal2 s 460570 159200 460626 160400 6 mprj_adr_o[9]
port 613 nsew signal tristate
rlabel metal2 s 431130 159200 431186 160400 6 mprj_cyc_o
port 614 nsew signal tristate
rlabel metal2 s 435362 159200 435418 160400 6 mprj_dat_i[0]
port 615 nsew signal input
rlabel metal2 s 463882 159200 463938 160400 6 mprj_dat_i[10]
port 616 nsew signal input
rlabel metal2 s 466458 159200 466514 160400 6 mprj_dat_i[11]
port 617 nsew signal input
rlabel metal2 s 468942 159200 468998 160400 6 mprj_dat_i[12]
port 618 nsew signal input
rlabel metal2 s 471426 159200 471482 160400 6 mprj_dat_i[13]
port 619 nsew signal input
rlabel metal2 s 474002 159200 474058 160400 6 mprj_dat_i[14]
port 620 nsew signal input
rlabel metal2 s 476486 159200 476542 160400 6 mprj_dat_i[15]
port 621 nsew signal input
rlabel metal2 s 479062 159200 479118 160400 6 mprj_dat_i[16]
port 622 nsew signal input
rlabel metal2 s 481546 159200 481602 160400 6 mprj_dat_i[17]
port 623 nsew signal input
rlabel metal2 s 484030 159200 484086 160400 6 mprj_dat_i[18]
port 624 nsew signal input
rlabel metal2 s 486606 159200 486662 160400 6 mprj_dat_i[19]
port 625 nsew signal input
rlabel metal2 s 438674 159200 438730 160400 6 mprj_dat_i[1]
port 626 nsew signal input
rlabel metal2 s 489090 159200 489146 160400 6 mprj_dat_i[20]
port 627 nsew signal input
rlabel metal2 s 491666 159200 491722 160400 6 mprj_dat_i[21]
port 628 nsew signal input
rlabel metal2 s 494150 159200 494206 160400 6 mprj_dat_i[22]
port 629 nsew signal input
rlabel metal2 s 496634 159200 496690 160400 6 mprj_dat_i[23]
port 630 nsew signal input
rlabel metal2 s 499210 159200 499266 160400 6 mprj_dat_i[24]
port 631 nsew signal input
rlabel metal2 s 501694 159200 501750 160400 6 mprj_dat_i[25]
port 632 nsew signal input
rlabel metal2 s 504178 159200 504234 160400 6 mprj_dat_i[26]
port 633 nsew signal input
rlabel metal2 s 506754 159200 506810 160400 6 mprj_dat_i[27]
port 634 nsew signal input
rlabel metal2 s 509238 159200 509294 160400 6 mprj_dat_i[28]
port 635 nsew signal input
rlabel metal2 s 511814 159200 511870 160400 6 mprj_dat_i[29]
port 636 nsew signal input
rlabel metal2 s 442078 159200 442134 160400 6 mprj_dat_i[2]
port 637 nsew signal input
rlabel metal2 s 514298 159200 514354 160400 6 mprj_dat_i[30]
port 638 nsew signal input
rlabel metal2 s 516782 159200 516838 160400 6 mprj_dat_i[31]
port 639 nsew signal input
rlabel metal2 s 445390 159200 445446 160400 6 mprj_dat_i[3]
port 640 nsew signal input
rlabel metal2 s 448794 159200 448850 160400 6 mprj_dat_i[4]
port 641 nsew signal input
rlabel metal2 s 451278 159200 451334 160400 6 mprj_dat_i[5]
port 642 nsew signal input
rlabel metal2 s 453854 159200 453910 160400 6 mprj_dat_i[6]
port 643 nsew signal input
rlabel metal2 s 456338 159200 456394 160400 6 mprj_dat_i[7]
port 644 nsew signal input
rlabel metal2 s 458914 159200 458970 160400 6 mprj_dat_i[8]
port 645 nsew signal input
rlabel metal2 s 461398 159200 461454 160400 6 mprj_dat_i[9]
port 646 nsew signal input
rlabel metal2 s 436190 159200 436246 160400 6 mprj_dat_o[0]
port 647 nsew signal tristate
rlabel metal2 s 464710 159200 464766 160400 6 mprj_dat_o[10]
port 648 nsew signal tristate
rlabel metal2 s 467286 159200 467342 160400 6 mprj_dat_o[11]
port 649 nsew signal tristate
rlabel metal2 s 469770 159200 469826 160400 6 mprj_dat_o[12]
port 650 nsew signal tristate
rlabel metal2 s 472346 159200 472402 160400 6 mprj_dat_o[13]
port 651 nsew signal tristate
rlabel metal2 s 474830 159200 474886 160400 6 mprj_dat_o[14]
port 652 nsew signal tristate
rlabel metal2 s 477314 159200 477370 160400 6 mprj_dat_o[15]
port 653 nsew signal tristate
rlabel metal2 s 479890 159200 479946 160400 6 mprj_dat_o[16]
port 654 nsew signal tristate
rlabel metal2 s 482374 159200 482430 160400 6 mprj_dat_o[17]
port 655 nsew signal tristate
rlabel metal2 s 484858 159200 484914 160400 6 mprj_dat_o[18]
port 656 nsew signal tristate
rlabel metal2 s 487434 159200 487490 160400 6 mprj_dat_o[19]
port 657 nsew signal tristate
rlabel metal2 s 439594 159200 439650 160400 6 mprj_dat_o[1]
port 658 nsew signal tristate
rlabel metal2 s 489918 159200 489974 160400 6 mprj_dat_o[20]
port 659 nsew signal tristate
rlabel metal2 s 492494 159200 492550 160400 6 mprj_dat_o[21]
port 660 nsew signal tristate
rlabel metal2 s 494978 159200 495034 160400 6 mprj_dat_o[22]
port 661 nsew signal tristate
rlabel metal2 s 497462 159200 497518 160400 6 mprj_dat_o[23]
port 662 nsew signal tristate
rlabel metal2 s 500038 159200 500094 160400 6 mprj_dat_o[24]
port 663 nsew signal tristate
rlabel metal2 s 502522 159200 502578 160400 6 mprj_dat_o[25]
port 664 nsew signal tristate
rlabel metal2 s 505098 159200 505154 160400 6 mprj_dat_o[26]
port 665 nsew signal tristate
rlabel metal2 s 507582 159200 507638 160400 6 mprj_dat_o[27]
port 666 nsew signal tristate
rlabel metal2 s 510066 159200 510122 160400 6 mprj_dat_o[28]
port 667 nsew signal tristate
rlabel metal2 s 512642 159200 512698 160400 6 mprj_dat_o[29]
port 668 nsew signal tristate
rlabel metal2 s 442906 159200 442962 160400 6 mprj_dat_o[2]
port 669 nsew signal tristate
rlabel metal2 s 515126 159200 515182 160400 6 mprj_dat_o[30]
port 670 nsew signal tristate
rlabel metal2 s 517610 159200 517666 160400 6 mprj_dat_o[31]
port 671 nsew signal tristate
rlabel metal2 s 446310 159200 446366 160400 6 mprj_dat_o[3]
port 672 nsew signal tristate
rlabel metal2 s 449622 159200 449678 160400 6 mprj_dat_o[4]
port 673 nsew signal tristate
rlabel metal2 s 452106 159200 452162 160400 6 mprj_dat_o[5]
port 674 nsew signal tristate
rlabel metal2 s 454682 159200 454738 160400 6 mprj_dat_o[6]
port 675 nsew signal tristate
rlabel metal2 s 457166 159200 457222 160400 6 mprj_dat_o[7]
port 676 nsew signal tristate
rlabel metal2 s 459742 159200 459798 160400 6 mprj_dat_o[8]
port 677 nsew signal tristate
rlabel metal2 s 462226 159200 462282 160400 6 mprj_dat_o[9]
port 678 nsew signal tristate
rlabel metal2 s 437018 159200 437074 160400 6 mprj_sel_o[0]
port 679 nsew signal tristate
rlabel metal2 s 440422 159200 440478 160400 6 mprj_sel_o[1]
port 680 nsew signal tristate
rlabel metal2 s 443734 159200 443790 160400 6 mprj_sel_o[2]
port 681 nsew signal tristate
rlabel metal2 s 447138 159200 447194 160400 6 mprj_sel_o[3]
port 682 nsew signal tristate
rlabel metal2 s 431958 159200 432014 160400 6 mprj_stb_o
port 683 nsew signal tristate
rlabel metal2 s 432878 159200 432934 160400 6 mprj_wb_iena
port 684 nsew signal tristate
rlabel metal2 s 433706 159200 433762 160400 6 mprj_we_o
port 685 nsew signal tristate
rlabel metal3 s 523200 88000 524400 88120 6 qspi_enabled
port 686 nsew signal tristate
rlabel metal3 s 523200 82016 524400 82136 6 ser_rx
port 687 nsew signal input
rlabel metal3 s 523200 83512 524400 83632 6 ser_tx
port 688 nsew signal tristate
rlabel metal3 s 523200 79160 524400 79280 6 spi_csb
port 689 nsew signal tristate
rlabel metal3 s 523200 85008 524400 85128 6 spi_enabled
port 690 nsew signal tristate
rlabel metal3 s 523200 77664 524400 77784 6 spi_sck
port 691 nsew signal tristate
rlabel metal3 s 523200 80656 524400 80776 6 spi_sdi
port 692 nsew signal input
rlabel metal3 s 523200 76168 524400 76288 6 spi_sdo
port 693 nsew signal tristate
rlabel metal3 s 523200 74672 524400 74792 6 spi_sdoenb
port 694 nsew signal tristate
rlabel metal3 s 523200 2048 524400 2168 6 sram_ro_addr[0]
port 695 nsew signal input
rlabel metal3 s 523200 3544 524400 3664 6 sram_ro_addr[1]
port 696 nsew signal input
rlabel metal3 s 523200 5040 524400 5160 6 sram_ro_addr[2]
port 697 nsew signal input
rlabel metal3 s 523200 6536 524400 6656 6 sram_ro_addr[3]
port 698 nsew signal input
rlabel metal3 s 523200 8032 524400 8152 6 sram_ro_addr[4]
port 699 nsew signal input
rlabel metal3 s 523200 9528 524400 9648 6 sram_ro_addr[5]
port 700 nsew signal input
rlabel metal3 s 523200 11024 524400 11144 6 sram_ro_addr[6]
port 701 nsew signal input
rlabel metal3 s 523200 12520 524400 12640 6 sram_ro_addr[7]
port 702 nsew signal input
rlabel metal3 s 523200 14016 524400 14136 6 sram_ro_clk
port 703 nsew signal input
rlabel metal3 s 523200 688 524400 808 6 sram_ro_csb
port 704 nsew signal input
rlabel metal3 s 523200 15376 524400 15496 6 sram_ro_data[0]
port 705 nsew signal tristate
rlabel metal3 s 523200 30200 524400 30320 6 sram_ro_data[10]
port 706 nsew signal tristate
rlabel metal3 s 523200 31696 524400 31816 6 sram_ro_data[11]
port 707 nsew signal tristate
rlabel metal3 s 523200 33192 524400 33312 6 sram_ro_data[12]
port 708 nsew signal tristate
rlabel metal3 s 523200 34688 524400 34808 6 sram_ro_data[13]
port 709 nsew signal tristate
rlabel metal3 s 523200 36184 524400 36304 6 sram_ro_data[14]
port 710 nsew signal tristate
rlabel metal3 s 523200 37680 524400 37800 6 sram_ro_data[15]
port 711 nsew signal tristate
rlabel metal3 s 523200 39176 524400 39296 6 sram_ro_data[16]
port 712 nsew signal tristate
rlabel metal3 s 523200 40672 524400 40792 6 sram_ro_data[17]
port 713 nsew signal tristate
rlabel metal3 s 523200 42032 524400 42152 6 sram_ro_data[18]
port 714 nsew signal tristate
rlabel metal3 s 523200 43528 524400 43648 6 sram_ro_data[19]
port 715 nsew signal tristate
rlabel metal3 s 523200 16872 524400 16992 6 sram_ro_data[1]
port 716 nsew signal tristate
rlabel metal3 s 523200 45024 524400 45144 6 sram_ro_data[20]
port 717 nsew signal tristate
rlabel metal3 s 523200 46520 524400 46640 6 sram_ro_data[21]
port 718 nsew signal tristate
rlabel metal3 s 523200 48016 524400 48136 6 sram_ro_data[22]
port 719 nsew signal tristate
rlabel metal3 s 523200 49512 524400 49632 6 sram_ro_data[23]
port 720 nsew signal tristate
rlabel metal3 s 523200 51008 524400 51128 6 sram_ro_data[24]
port 721 nsew signal tristate
rlabel metal3 s 523200 52504 524400 52624 6 sram_ro_data[25]
port 722 nsew signal tristate
rlabel metal3 s 523200 54000 524400 54120 6 sram_ro_data[26]
port 723 nsew signal tristate
rlabel metal3 s 523200 55360 524400 55480 6 sram_ro_data[27]
port 724 nsew signal tristate
rlabel metal3 s 523200 56856 524400 56976 6 sram_ro_data[28]
port 725 nsew signal tristate
rlabel metal3 s 523200 58352 524400 58472 6 sram_ro_data[29]
port 726 nsew signal tristate
rlabel metal3 s 523200 18368 524400 18488 6 sram_ro_data[2]
port 727 nsew signal tristate
rlabel metal3 s 523200 59848 524400 59968 6 sram_ro_data[30]
port 728 nsew signal tristate
rlabel metal3 s 523200 61344 524400 61464 6 sram_ro_data[31]
port 729 nsew signal tristate
rlabel metal3 s 523200 19864 524400 19984 6 sram_ro_data[3]
port 730 nsew signal tristate
rlabel metal3 s 523200 21360 524400 21480 6 sram_ro_data[4]
port 731 nsew signal tristate
rlabel metal3 s 523200 22856 524400 22976 6 sram_ro_data[5]
port 732 nsew signal tristate
rlabel metal3 s 523200 24352 524400 24472 6 sram_ro_data[6]
port 733 nsew signal tristate
rlabel metal3 s 523200 25848 524400 25968 6 sram_ro_data[7]
port 734 nsew signal tristate
rlabel metal3 s 523200 27344 524400 27464 6 sram_ro_data[8]
port 735 nsew signal tristate
rlabel metal3 s 523200 28704 524400 28824 6 sram_ro_data[9]
port 736 nsew signal tristate
rlabel metal3 s 523200 68688 524400 68808 6 trap
port 737 nsew signal tristate
rlabel metal3 s 523200 86504 524400 86624 6 uart_enabled
port 738 nsew signal tristate
rlabel metal2 s 518530 159200 518586 160400 6 user_irq_ena[0]
port 739 nsew signal tristate
rlabel metal2 s 519358 159200 519414 160400 6 user_irq_ena[1]
port 740 nsew signal tristate
rlabel metal2 s 520186 159200 520242 160400 6 user_irq_ena[2]
port 741 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 524000 160000
<< end >>
