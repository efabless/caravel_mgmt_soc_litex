magic
tech sky130A
magscale 1 2
timestamp 1668011404
<< obsli1 >>
rect 2024 2703 521916 161041
<< obsm1 >>
rect 2024 2672 521916 163804
<< metal2 >>
rect 3606 163200 3662 164000
rect 4434 163200 4490 164000
rect 5262 163200 5318 164000
rect 6090 163200 6146 164000
rect 6918 163200 6974 164000
rect 7746 163200 7802 164000
rect 8574 163200 8630 164000
rect 9402 163200 9458 164000
rect 10230 163200 10286 164000
rect 11058 163200 11114 164000
rect 11886 163200 11942 164000
rect 12714 163200 12770 164000
rect 13542 163200 13598 164000
rect 14370 163200 14426 164000
rect 15198 163200 15254 164000
rect 16026 163200 16082 164000
rect 16854 163200 16910 164000
rect 17682 163200 17738 164000
rect 18510 163200 18566 164000
rect 19338 163200 19394 164000
rect 20166 163200 20222 164000
rect 20994 163200 21050 164000
rect 21822 163200 21878 164000
rect 22650 163200 22706 164000
rect 23478 163200 23534 164000
rect 24306 163200 24362 164000
rect 25134 163200 25190 164000
rect 25962 163200 26018 164000
rect 26790 163200 26846 164000
rect 27618 163200 27674 164000
rect 28446 163200 28502 164000
rect 29274 163200 29330 164000
rect 30102 163200 30158 164000
rect 30930 163200 30986 164000
rect 31758 163200 31814 164000
rect 32586 163200 32642 164000
rect 33414 163200 33470 164000
rect 34242 163200 34298 164000
rect 35070 163200 35126 164000
rect 35898 163200 35954 164000
rect 36726 163200 36782 164000
rect 37554 163200 37610 164000
rect 38382 163200 38438 164000
rect 39210 163200 39266 164000
rect 40038 163200 40094 164000
rect 40866 163200 40922 164000
rect 41694 163200 41750 164000
rect 42522 163200 42578 164000
rect 43350 163200 43406 164000
rect 44178 163200 44234 164000
rect 45006 163200 45062 164000
rect 45834 163200 45890 164000
rect 46662 163200 46718 164000
rect 47490 163200 47546 164000
rect 48318 163200 48374 164000
rect 49146 163200 49202 164000
rect 49974 163200 50030 164000
rect 50802 163200 50858 164000
rect 51630 163200 51686 164000
rect 52458 163200 52514 164000
rect 53286 163200 53342 164000
rect 54114 163200 54170 164000
rect 54942 163200 54998 164000
rect 55770 163200 55826 164000
rect 56598 163200 56654 164000
rect 57426 163200 57482 164000
rect 58254 163200 58310 164000
rect 59082 163200 59138 164000
rect 59910 163200 59966 164000
rect 60738 163200 60794 164000
rect 61566 163200 61622 164000
rect 62394 163200 62450 164000
rect 63222 163200 63278 164000
rect 64050 163200 64106 164000
rect 64878 163200 64934 164000
rect 65706 163200 65762 164000
rect 66534 163200 66590 164000
rect 67362 163200 67418 164000
rect 68190 163200 68246 164000
rect 69018 163200 69074 164000
rect 69846 163200 69902 164000
rect 70674 163200 70730 164000
rect 71502 163200 71558 164000
rect 72330 163200 72386 164000
rect 73158 163200 73214 164000
rect 73986 163200 74042 164000
rect 74814 163200 74870 164000
rect 75642 163200 75698 164000
rect 76470 163200 76526 164000
rect 77298 163200 77354 164000
rect 78126 163200 78182 164000
rect 78954 163200 79010 164000
rect 79782 163200 79838 164000
rect 80610 163200 80666 164000
rect 81438 163200 81494 164000
rect 82266 163200 82322 164000
rect 83094 163200 83150 164000
rect 83922 163200 83978 164000
rect 84750 163200 84806 164000
rect 85578 163200 85634 164000
rect 86406 163200 86462 164000
rect 87234 163200 87290 164000
rect 88062 163200 88118 164000
rect 88890 163200 88946 164000
rect 89718 163200 89774 164000
rect 90546 163200 90602 164000
rect 91374 163200 91430 164000
rect 92202 163200 92258 164000
rect 93030 163200 93086 164000
rect 93858 163200 93914 164000
rect 94686 163200 94742 164000
rect 95514 163200 95570 164000
rect 96342 163200 96398 164000
rect 97170 163200 97226 164000
rect 97998 163200 98054 164000
rect 98826 163200 98882 164000
rect 99654 163200 99710 164000
rect 100482 163200 100538 164000
rect 101310 163200 101366 164000
rect 102138 163200 102194 164000
rect 102966 163200 103022 164000
rect 103794 163200 103850 164000
rect 104622 163200 104678 164000
rect 105450 163200 105506 164000
rect 106278 163200 106334 164000
rect 107106 163200 107162 164000
rect 107934 163200 107990 164000
rect 108762 163200 108818 164000
rect 109590 163200 109646 164000
rect 110418 163200 110474 164000
rect 111246 163200 111302 164000
rect 112074 163200 112130 164000
rect 112902 163200 112958 164000
rect 113730 163200 113786 164000
rect 114558 163200 114614 164000
rect 115386 163200 115442 164000
rect 116214 163200 116270 164000
rect 117042 163200 117098 164000
rect 117870 163200 117926 164000
rect 118698 163200 118754 164000
rect 119526 163200 119582 164000
rect 120354 163200 120410 164000
rect 121182 163200 121238 164000
rect 122010 163200 122066 164000
rect 122838 163200 122894 164000
rect 123666 163200 123722 164000
rect 124494 163200 124550 164000
rect 125322 163200 125378 164000
rect 126150 163200 126206 164000
rect 126978 163200 127034 164000
rect 127806 163200 127862 164000
rect 128634 163200 128690 164000
rect 129462 163200 129518 164000
rect 130290 163200 130346 164000
rect 131118 163200 131174 164000
rect 131946 163200 132002 164000
rect 132774 163200 132830 164000
rect 133602 163200 133658 164000
rect 134430 163200 134486 164000
rect 135258 163200 135314 164000
rect 136086 163200 136142 164000
rect 136914 163200 136970 164000
rect 137742 163200 137798 164000
rect 138570 163200 138626 164000
rect 139398 163200 139454 164000
rect 140226 163200 140282 164000
rect 141054 163200 141110 164000
rect 141882 163200 141938 164000
rect 142710 163200 142766 164000
rect 143538 163200 143594 164000
rect 144366 163200 144422 164000
rect 145194 163200 145250 164000
rect 146022 163200 146078 164000
rect 146850 163200 146906 164000
rect 147678 163200 147734 164000
rect 148506 163200 148562 164000
rect 149334 163200 149390 164000
rect 150162 163200 150218 164000
rect 150990 163200 151046 164000
rect 151818 163200 151874 164000
rect 152646 163200 152702 164000
rect 153474 163200 153530 164000
rect 154302 163200 154358 164000
rect 155130 163200 155186 164000
rect 155958 163200 156014 164000
rect 156786 163200 156842 164000
rect 157614 163200 157670 164000
rect 158442 163200 158498 164000
rect 159270 163200 159326 164000
rect 160098 163200 160154 164000
rect 160926 163200 160982 164000
rect 161754 163200 161810 164000
rect 162582 163200 162638 164000
rect 163410 163200 163466 164000
rect 164238 163200 164294 164000
rect 165066 163200 165122 164000
rect 165894 163200 165950 164000
rect 166722 163200 166778 164000
rect 167550 163200 167606 164000
rect 168378 163200 168434 164000
rect 169206 163200 169262 164000
rect 170034 163200 170090 164000
rect 170862 163200 170918 164000
rect 171690 163200 171746 164000
rect 172518 163200 172574 164000
rect 173346 163200 173402 164000
rect 174174 163200 174230 164000
rect 175002 163200 175058 164000
rect 175830 163200 175886 164000
rect 176658 163200 176714 164000
rect 177486 163200 177542 164000
rect 178314 163200 178370 164000
rect 179142 163200 179198 164000
rect 179970 163200 180026 164000
rect 180798 163200 180854 164000
rect 181626 163200 181682 164000
rect 182454 163200 182510 164000
rect 183282 163200 183338 164000
rect 184110 163200 184166 164000
rect 184938 163200 184994 164000
rect 185766 163200 185822 164000
rect 186594 163200 186650 164000
rect 187422 163200 187478 164000
rect 188250 163200 188306 164000
rect 189078 163200 189134 164000
rect 189906 163200 189962 164000
rect 190734 163200 190790 164000
rect 191562 163200 191618 164000
rect 192390 163200 192446 164000
rect 193218 163200 193274 164000
rect 194046 163200 194102 164000
rect 194874 163200 194930 164000
rect 195702 163200 195758 164000
rect 196530 163200 196586 164000
rect 197358 163200 197414 164000
rect 198186 163200 198242 164000
rect 199014 163200 199070 164000
rect 199842 163200 199898 164000
rect 200670 163200 200726 164000
rect 201498 163200 201554 164000
rect 202326 163200 202382 164000
rect 203154 163200 203210 164000
rect 203982 163200 204038 164000
rect 204810 163200 204866 164000
rect 205638 163200 205694 164000
rect 206466 163200 206522 164000
rect 207294 163200 207350 164000
rect 208122 163200 208178 164000
rect 208950 163200 209006 164000
rect 209778 163200 209834 164000
rect 210606 163200 210662 164000
rect 211434 163200 211490 164000
rect 212262 163200 212318 164000
rect 213090 163200 213146 164000
rect 213918 163200 213974 164000
rect 214746 163200 214802 164000
rect 215574 163200 215630 164000
rect 216402 163200 216458 164000
rect 217230 163200 217286 164000
rect 218058 163200 218114 164000
rect 218886 163200 218942 164000
rect 219714 163200 219770 164000
rect 220542 163200 220598 164000
rect 221370 163200 221426 164000
rect 222198 163200 222254 164000
rect 223026 163200 223082 164000
rect 223854 163200 223910 164000
rect 224682 163200 224738 164000
rect 225510 163200 225566 164000
rect 226338 163200 226394 164000
rect 227166 163200 227222 164000
rect 227994 163200 228050 164000
rect 228822 163200 228878 164000
rect 229650 163200 229706 164000
rect 230478 163200 230534 164000
rect 231306 163200 231362 164000
rect 232134 163200 232190 164000
rect 232962 163200 233018 164000
rect 233790 163200 233846 164000
rect 234618 163200 234674 164000
rect 235446 163200 235502 164000
rect 236274 163200 236330 164000
rect 237102 163200 237158 164000
rect 237930 163200 237986 164000
rect 238758 163200 238814 164000
rect 239586 163200 239642 164000
rect 240414 163200 240470 164000
rect 241242 163200 241298 164000
rect 242070 163200 242126 164000
rect 242898 163200 242954 164000
rect 243726 163200 243782 164000
rect 244554 163200 244610 164000
rect 245382 163200 245438 164000
rect 246210 163200 246266 164000
rect 247038 163200 247094 164000
rect 247866 163200 247922 164000
rect 248694 163200 248750 164000
rect 249522 163200 249578 164000
rect 250350 163200 250406 164000
rect 251178 163200 251234 164000
rect 252006 163200 252062 164000
rect 252834 163200 252890 164000
rect 253662 163200 253718 164000
rect 254490 163200 254546 164000
rect 255318 163200 255374 164000
rect 256146 163200 256202 164000
rect 256974 163200 257030 164000
rect 257802 163200 257858 164000
rect 258630 163200 258686 164000
rect 259458 163200 259514 164000
rect 260286 163200 260342 164000
rect 261114 163200 261170 164000
rect 261942 163200 261998 164000
rect 262770 163200 262826 164000
rect 263598 163200 263654 164000
rect 264426 163200 264482 164000
rect 265254 163200 265310 164000
rect 266082 163200 266138 164000
rect 266910 163200 266966 164000
rect 267738 163200 267794 164000
rect 268566 163200 268622 164000
rect 269394 163200 269450 164000
rect 270222 163200 270278 164000
rect 271050 163200 271106 164000
rect 271878 163200 271934 164000
rect 272706 163200 272762 164000
rect 273534 163200 273590 164000
rect 274362 163200 274418 164000
rect 275190 163200 275246 164000
rect 276018 163200 276074 164000
rect 276846 163200 276902 164000
rect 277674 163200 277730 164000
rect 278502 163200 278558 164000
rect 279330 163200 279386 164000
rect 280158 163200 280214 164000
rect 280986 163200 281042 164000
rect 281814 163200 281870 164000
rect 282642 163200 282698 164000
rect 283470 163200 283526 164000
rect 284298 163200 284354 164000
rect 285126 163200 285182 164000
rect 285954 163200 286010 164000
rect 286782 163200 286838 164000
rect 287610 163200 287666 164000
rect 288438 163200 288494 164000
rect 289266 163200 289322 164000
rect 290094 163200 290150 164000
rect 290922 163200 290978 164000
rect 291750 163200 291806 164000
rect 292578 163200 292634 164000
rect 293406 163200 293462 164000
rect 294234 163200 294290 164000
rect 295062 163200 295118 164000
rect 295890 163200 295946 164000
rect 296718 163200 296774 164000
rect 297546 163200 297602 164000
rect 298374 163200 298430 164000
rect 299202 163200 299258 164000
rect 300030 163200 300086 164000
rect 300858 163200 300914 164000
rect 301686 163200 301742 164000
rect 302514 163200 302570 164000
rect 303342 163200 303398 164000
rect 304170 163200 304226 164000
rect 304998 163200 305054 164000
rect 305826 163200 305882 164000
rect 306654 163200 306710 164000
rect 307482 163200 307538 164000
rect 308310 163200 308366 164000
rect 309138 163200 309194 164000
rect 309966 163200 310022 164000
rect 310794 163200 310850 164000
rect 311622 163200 311678 164000
rect 312450 163200 312506 164000
rect 313278 163200 313334 164000
rect 314106 163200 314162 164000
rect 314934 163200 314990 164000
rect 315762 163200 315818 164000
rect 316590 163200 316646 164000
rect 317418 163200 317474 164000
rect 318246 163200 318302 164000
rect 319074 163200 319130 164000
rect 319902 163200 319958 164000
rect 320730 163200 320786 164000
rect 321558 163200 321614 164000
rect 322386 163200 322442 164000
rect 323214 163200 323270 164000
rect 324042 163200 324098 164000
rect 324870 163200 324926 164000
rect 325698 163200 325754 164000
rect 326526 163200 326582 164000
rect 327354 163200 327410 164000
rect 328182 163200 328238 164000
rect 329010 163200 329066 164000
rect 329838 163200 329894 164000
rect 330666 163200 330722 164000
rect 331494 163200 331550 164000
rect 332322 163200 332378 164000
rect 333150 163200 333206 164000
rect 333978 163200 334034 164000
rect 334806 163200 334862 164000
rect 335634 163200 335690 164000
rect 336462 163200 336518 164000
rect 337290 163200 337346 164000
rect 338118 163200 338174 164000
rect 338946 163200 339002 164000
rect 339774 163200 339830 164000
rect 340602 163200 340658 164000
rect 341430 163200 341486 164000
rect 342258 163200 342314 164000
rect 343086 163200 343142 164000
rect 343914 163200 343970 164000
rect 344742 163200 344798 164000
rect 345570 163200 345626 164000
rect 346398 163200 346454 164000
rect 347226 163200 347282 164000
rect 348054 163200 348110 164000
rect 348882 163200 348938 164000
rect 349710 163200 349766 164000
rect 350538 163200 350594 164000
rect 351366 163200 351422 164000
rect 352194 163200 352250 164000
rect 353022 163200 353078 164000
rect 353850 163200 353906 164000
rect 354678 163200 354734 164000
rect 355506 163200 355562 164000
rect 356334 163200 356390 164000
rect 357162 163200 357218 164000
rect 357990 163200 358046 164000
rect 358818 163200 358874 164000
rect 359646 163200 359702 164000
rect 360474 163200 360530 164000
rect 361302 163200 361358 164000
rect 362130 163200 362186 164000
rect 362958 163200 363014 164000
rect 363786 163200 363842 164000
rect 364614 163200 364670 164000
rect 365442 163200 365498 164000
rect 366270 163200 366326 164000
rect 367098 163200 367154 164000
rect 367926 163200 367982 164000
rect 368754 163200 368810 164000
rect 369582 163200 369638 164000
rect 370410 163200 370466 164000
rect 371238 163200 371294 164000
rect 372066 163200 372122 164000
rect 372894 163200 372950 164000
rect 373722 163200 373778 164000
rect 374550 163200 374606 164000
rect 375378 163200 375434 164000
rect 376206 163200 376262 164000
rect 377034 163200 377090 164000
rect 377862 163200 377918 164000
rect 378690 163200 378746 164000
rect 379518 163200 379574 164000
rect 380346 163200 380402 164000
rect 381174 163200 381230 164000
rect 382002 163200 382058 164000
rect 382830 163200 382886 164000
rect 383658 163200 383714 164000
rect 384486 163200 384542 164000
rect 385314 163200 385370 164000
rect 386142 163200 386198 164000
rect 386970 163200 387026 164000
rect 387798 163200 387854 164000
rect 388626 163200 388682 164000
rect 389454 163200 389510 164000
rect 390282 163200 390338 164000
rect 391110 163200 391166 164000
rect 391938 163200 391994 164000
rect 392766 163200 392822 164000
rect 393594 163200 393650 164000
rect 394422 163200 394478 164000
rect 395250 163200 395306 164000
rect 396078 163200 396134 164000
rect 396906 163200 396962 164000
rect 397734 163200 397790 164000
rect 398562 163200 398618 164000
rect 399390 163200 399446 164000
rect 400218 163200 400274 164000
rect 401046 163200 401102 164000
rect 401874 163200 401930 164000
rect 402702 163200 402758 164000
rect 403530 163200 403586 164000
rect 404358 163200 404414 164000
rect 405186 163200 405242 164000
rect 406014 163200 406070 164000
rect 406842 163200 406898 164000
rect 407670 163200 407726 164000
rect 408498 163200 408554 164000
rect 409326 163200 409382 164000
rect 410154 163200 410210 164000
rect 410982 163200 411038 164000
rect 411810 163200 411866 164000
rect 412638 163200 412694 164000
rect 413466 163200 413522 164000
rect 414294 163200 414350 164000
rect 415122 163200 415178 164000
rect 415950 163200 416006 164000
rect 416778 163200 416834 164000
rect 417606 163200 417662 164000
rect 418434 163200 418490 164000
rect 419262 163200 419318 164000
rect 420090 163200 420146 164000
rect 420918 163200 420974 164000
rect 421746 163200 421802 164000
rect 422574 163200 422630 164000
rect 423402 163200 423458 164000
rect 424230 163200 424286 164000
rect 425058 163200 425114 164000
rect 425886 163200 425942 164000
rect 426714 163200 426770 164000
rect 427542 163200 427598 164000
rect 428370 163200 428426 164000
rect 429198 163200 429254 164000
rect 430026 163200 430082 164000
rect 430854 163200 430910 164000
rect 431682 163200 431738 164000
rect 432510 163200 432566 164000
rect 433338 163200 433394 164000
rect 434166 163200 434222 164000
rect 434994 163200 435050 164000
rect 435822 163200 435878 164000
rect 436650 163200 436706 164000
rect 437478 163200 437534 164000
rect 438306 163200 438362 164000
rect 439134 163200 439190 164000
rect 439962 163200 440018 164000
rect 440790 163200 440846 164000
rect 441618 163200 441674 164000
rect 442446 163200 442502 164000
rect 443274 163200 443330 164000
rect 444102 163200 444158 164000
rect 444930 163200 444986 164000
rect 445758 163200 445814 164000
rect 446586 163200 446642 164000
rect 447414 163200 447470 164000
rect 448242 163200 448298 164000
rect 449070 163200 449126 164000
rect 449898 163200 449954 164000
rect 450726 163200 450782 164000
rect 451554 163200 451610 164000
rect 452382 163200 452438 164000
rect 453210 163200 453266 164000
rect 454038 163200 454094 164000
rect 454866 163200 454922 164000
rect 455694 163200 455750 164000
rect 456522 163200 456578 164000
rect 457350 163200 457406 164000
rect 458178 163200 458234 164000
rect 459006 163200 459062 164000
rect 459834 163200 459890 164000
rect 460662 163200 460718 164000
rect 461490 163200 461546 164000
rect 462318 163200 462374 164000
rect 463146 163200 463202 164000
rect 463974 163200 464030 164000
rect 464802 163200 464858 164000
rect 465630 163200 465686 164000
rect 466458 163200 466514 164000
rect 467286 163200 467342 164000
rect 468114 163200 468170 164000
rect 468942 163200 468998 164000
rect 469770 163200 469826 164000
rect 470598 163200 470654 164000
rect 471426 163200 471482 164000
rect 472254 163200 472310 164000
rect 473082 163200 473138 164000
rect 473910 163200 473966 164000
rect 474738 163200 474794 164000
rect 475566 163200 475622 164000
rect 476394 163200 476450 164000
rect 477222 163200 477278 164000
rect 478050 163200 478106 164000
rect 478878 163200 478934 164000
rect 479706 163200 479762 164000
rect 480534 163200 480590 164000
rect 481362 163200 481418 164000
rect 482190 163200 482246 164000
rect 483018 163200 483074 164000
rect 483846 163200 483902 164000
rect 484674 163200 484730 164000
rect 485502 163200 485558 164000
rect 486330 163200 486386 164000
rect 487158 163200 487214 164000
rect 487986 163200 488042 164000
rect 488814 163200 488870 164000
rect 489642 163200 489698 164000
rect 490470 163200 490526 164000
rect 491298 163200 491354 164000
rect 492126 163200 492182 164000
rect 492954 163200 493010 164000
rect 493782 163200 493838 164000
rect 494610 163200 494666 164000
rect 495438 163200 495494 164000
rect 496266 163200 496322 164000
rect 497094 163200 497150 164000
rect 497922 163200 497978 164000
rect 498750 163200 498806 164000
rect 499578 163200 499634 164000
rect 500406 163200 500462 164000
rect 501234 163200 501290 164000
rect 502062 163200 502118 164000
rect 502890 163200 502946 164000
rect 503718 163200 503774 164000
rect 504546 163200 504602 164000
rect 505374 163200 505430 164000
rect 506202 163200 506258 164000
rect 507030 163200 507086 164000
rect 507858 163200 507914 164000
rect 508686 163200 508742 164000
rect 509514 163200 509570 164000
rect 510342 163200 510398 164000
rect 511170 163200 511226 164000
rect 511998 163200 512054 164000
rect 512826 163200 512882 164000
rect 513654 163200 513710 164000
rect 514482 163200 514538 164000
rect 515310 163200 515366 164000
rect 516138 163200 516194 164000
rect 516966 163200 517022 164000
rect 517794 163200 517850 164000
rect 518622 163200 518678 164000
rect 519450 163200 519506 164000
rect 520278 163200 520334 164000
rect 253972 0 254028 800
rect 255972 0 256028 800
rect 257972 0 258028 800
rect 259972 0 260028 800
rect 261972 0 262028 800
rect 263972 0 264028 800
rect 265972 0 266028 800
rect 491972 0 492028 800
rect 493972 0 494028 800
rect 495972 0 496028 800
rect 497972 0 498028 800
rect 499972 0 500028 800
rect 501972 0 502028 800
<< obsm2 >>
rect 2870 163144 3550 163810
rect 3718 163144 4378 163810
rect 4546 163144 5206 163810
rect 5374 163144 6034 163810
rect 6202 163144 6862 163810
rect 7030 163144 7690 163810
rect 7858 163144 8518 163810
rect 8686 163144 9346 163810
rect 9514 163144 10174 163810
rect 10342 163144 11002 163810
rect 11170 163144 11830 163810
rect 11998 163144 12658 163810
rect 12826 163144 13486 163810
rect 13654 163144 14314 163810
rect 14482 163144 15142 163810
rect 15310 163144 15970 163810
rect 16138 163144 16798 163810
rect 16966 163144 17626 163810
rect 17794 163144 18454 163810
rect 18622 163144 19282 163810
rect 19450 163144 20110 163810
rect 20278 163144 20938 163810
rect 21106 163144 21766 163810
rect 21934 163144 22594 163810
rect 22762 163144 23422 163810
rect 23590 163144 24250 163810
rect 24418 163144 25078 163810
rect 25246 163144 25906 163810
rect 26074 163144 26734 163810
rect 26902 163144 27562 163810
rect 27730 163144 28390 163810
rect 28558 163144 29218 163810
rect 29386 163144 30046 163810
rect 30214 163144 30874 163810
rect 31042 163144 31702 163810
rect 31870 163144 32530 163810
rect 32698 163144 33358 163810
rect 33526 163144 34186 163810
rect 34354 163144 35014 163810
rect 35182 163144 35842 163810
rect 36010 163144 36670 163810
rect 36838 163144 37498 163810
rect 37666 163144 38326 163810
rect 38494 163144 39154 163810
rect 39322 163144 39982 163810
rect 40150 163144 40810 163810
rect 40978 163144 41638 163810
rect 41806 163144 42466 163810
rect 42634 163144 43294 163810
rect 43462 163144 44122 163810
rect 44290 163144 44950 163810
rect 45118 163144 45778 163810
rect 45946 163144 46606 163810
rect 46774 163144 47434 163810
rect 47602 163144 48262 163810
rect 48430 163144 49090 163810
rect 49258 163144 49918 163810
rect 50086 163144 50746 163810
rect 50914 163144 51574 163810
rect 51742 163144 52402 163810
rect 52570 163144 53230 163810
rect 53398 163144 54058 163810
rect 54226 163144 54886 163810
rect 55054 163144 55714 163810
rect 55882 163144 56542 163810
rect 56710 163144 57370 163810
rect 57538 163144 58198 163810
rect 58366 163144 59026 163810
rect 59194 163144 59854 163810
rect 60022 163144 60682 163810
rect 60850 163144 61510 163810
rect 61678 163144 62338 163810
rect 62506 163144 63166 163810
rect 63334 163144 63994 163810
rect 64162 163144 64822 163810
rect 64990 163144 65650 163810
rect 65818 163144 66478 163810
rect 66646 163144 67306 163810
rect 67474 163144 68134 163810
rect 68302 163144 68962 163810
rect 69130 163144 69790 163810
rect 69958 163144 70618 163810
rect 70786 163144 71446 163810
rect 71614 163144 72274 163810
rect 72442 163144 73102 163810
rect 73270 163144 73930 163810
rect 74098 163144 74758 163810
rect 74926 163144 75586 163810
rect 75754 163144 76414 163810
rect 76582 163144 77242 163810
rect 77410 163144 78070 163810
rect 78238 163144 78898 163810
rect 79066 163144 79726 163810
rect 79894 163144 80554 163810
rect 80722 163144 81382 163810
rect 81550 163144 82210 163810
rect 82378 163144 83038 163810
rect 83206 163144 83866 163810
rect 84034 163144 84694 163810
rect 84862 163144 85522 163810
rect 85690 163144 86350 163810
rect 86518 163144 87178 163810
rect 87346 163144 88006 163810
rect 88174 163144 88834 163810
rect 89002 163144 89662 163810
rect 89830 163144 90490 163810
rect 90658 163144 91318 163810
rect 91486 163144 92146 163810
rect 92314 163144 92974 163810
rect 93142 163144 93802 163810
rect 93970 163144 94630 163810
rect 94798 163144 95458 163810
rect 95626 163144 96286 163810
rect 96454 163144 97114 163810
rect 97282 163144 97942 163810
rect 98110 163144 98770 163810
rect 98938 163144 99598 163810
rect 99766 163144 100426 163810
rect 100594 163144 101254 163810
rect 101422 163144 102082 163810
rect 102250 163144 102910 163810
rect 103078 163144 103738 163810
rect 103906 163144 104566 163810
rect 104734 163144 105394 163810
rect 105562 163144 106222 163810
rect 106390 163144 107050 163810
rect 107218 163144 107878 163810
rect 108046 163144 108706 163810
rect 108874 163144 109534 163810
rect 109702 163144 110362 163810
rect 110530 163144 111190 163810
rect 111358 163144 112018 163810
rect 112186 163144 112846 163810
rect 113014 163144 113674 163810
rect 113842 163144 114502 163810
rect 114670 163144 115330 163810
rect 115498 163144 116158 163810
rect 116326 163144 116986 163810
rect 117154 163144 117814 163810
rect 117982 163144 118642 163810
rect 118810 163144 119470 163810
rect 119638 163144 120298 163810
rect 120466 163144 121126 163810
rect 121294 163144 121954 163810
rect 122122 163144 122782 163810
rect 122950 163144 123610 163810
rect 123778 163144 124438 163810
rect 124606 163144 125266 163810
rect 125434 163144 126094 163810
rect 126262 163144 126922 163810
rect 127090 163144 127750 163810
rect 127918 163144 128578 163810
rect 128746 163144 129406 163810
rect 129574 163144 130234 163810
rect 130402 163144 131062 163810
rect 131230 163144 131890 163810
rect 132058 163144 132718 163810
rect 132886 163144 133546 163810
rect 133714 163144 134374 163810
rect 134542 163144 135202 163810
rect 135370 163144 136030 163810
rect 136198 163144 136858 163810
rect 137026 163144 137686 163810
rect 137854 163144 138514 163810
rect 138682 163144 139342 163810
rect 139510 163144 140170 163810
rect 140338 163144 140998 163810
rect 141166 163144 141826 163810
rect 141994 163144 142654 163810
rect 142822 163144 143482 163810
rect 143650 163144 144310 163810
rect 144478 163144 145138 163810
rect 145306 163144 145966 163810
rect 146134 163144 146794 163810
rect 146962 163144 147622 163810
rect 147790 163144 148450 163810
rect 148618 163144 149278 163810
rect 149446 163144 150106 163810
rect 150274 163144 150934 163810
rect 151102 163144 151762 163810
rect 151930 163144 152590 163810
rect 152758 163144 153418 163810
rect 153586 163144 154246 163810
rect 154414 163144 155074 163810
rect 155242 163144 155902 163810
rect 156070 163144 156730 163810
rect 156898 163144 157558 163810
rect 157726 163144 158386 163810
rect 158554 163144 159214 163810
rect 159382 163144 160042 163810
rect 160210 163144 160870 163810
rect 161038 163144 161698 163810
rect 161866 163144 162526 163810
rect 162694 163144 163354 163810
rect 163522 163144 164182 163810
rect 164350 163144 165010 163810
rect 165178 163144 165838 163810
rect 166006 163144 166666 163810
rect 166834 163144 167494 163810
rect 167662 163144 168322 163810
rect 168490 163144 169150 163810
rect 169318 163144 169978 163810
rect 170146 163144 170806 163810
rect 170974 163144 171634 163810
rect 171802 163144 172462 163810
rect 172630 163144 173290 163810
rect 173458 163144 174118 163810
rect 174286 163144 174946 163810
rect 175114 163144 175774 163810
rect 175942 163144 176602 163810
rect 176770 163144 177430 163810
rect 177598 163144 178258 163810
rect 178426 163144 179086 163810
rect 179254 163144 179914 163810
rect 180082 163144 180742 163810
rect 180910 163144 181570 163810
rect 181738 163144 182398 163810
rect 182566 163144 183226 163810
rect 183394 163144 184054 163810
rect 184222 163144 184882 163810
rect 185050 163144 185710 163810
rect 185878 163144 186538 163810
rect 186706 163144 187366 163810
rect 187534 163144 188194 163810
rect 188362 163144 189022 163810
rect 189190 163144 189850 163810
rect 190018 163144 190678 163810
rect 190846 163144 191506 163810
rect 191674 163144 192334 163810
rect 192502 163144 193162 163810
rect 193330 163144 193990 163810
rect 194158 163144 194818 163810
rect 194986 163144 195646 163810
rect 195814 163144 196474 163810
rect 196642 163144 197302 163810
rect 197470 163144 198130 163810
rect 198298 163144 198958 163810
rect 199126 163144 199786 163810
rect 199954 163144 200614 163810
rect 200782 163144 201442 163810
rect 201610 163144 202270 163810
rect 202438 163144 203098 163810
rect 203266 163144 203926 163810
rect 204094 163144 204754 163810
rect 204922 163144 205582 163810
rect 205750 163144 206410 163810
rect 206578 163144 207238 163810
rect 207406 163144 208066 163810
rect 208234 163144 208894 163810
rect 209062 163144 209722 163810
rect 209890 163144 210550 163810
rect 210718 163144 211378 163810
rect 211546 163144 212206 163810
rect 212374 163144 213034 163810
rect 213202 163144 213862 163810
rect 214030 163144 214690 163810
rect 214858 163144 215518 163810
rect 215686 163144 216346 163810
rect 216514 163144 217174 163810
rect 217342 163144 218002 163810
rect 218170 163144 218830 163810
rect 218998 163144 219658 163810
rect 219826 163144 220486 163810
rect 220654 163144 221314 163810
rect 221482 163144 222142 163810
rect 222310 163144 222970 163810
rect 223138 163144 223798 163810
rect 223966 163144 224626 163810
rect 224794 163144 225454 163810
rect 225622 163144 226282 163810
rect 226450 163144 227110 163810
rect 227278 163144 227938 163810
rect 228106 163144 228766 163810
rect 228934 163144 229594 163810
rect 229762 163144 230422 163810
rect 230590 163144 231250 163810
rect 231418 163144 232078 163810
rect 232246 163144 232906 163810
rect 233074 163144 233734 163810
rect 233902 163144 234562 163810
rect 234730 163144 235390 163810
rect 235558 163144 236218 163810
rect 236386 163144 237046 163810
rect 237214 163144 237874 163810
rect 238042 163144 238702 163810
rect 238870 163144 239530 163810
rect 239698 163144 240358 163810
rect 240526 163144 241186 163810
rect 241354 163144 242014 163810
rect 242182 163144 242842 163810
rect 243010 163144 243670 163810
rect 243838 163144 244498 163810
rect 244666 163144 245326 163810
rect 245494 163144 246154 163810
rect 246322 163144 246982 163810
rect 247150 163144 247810 163810
rect 247978 163144 248638 163810
rect 248806 163144 249466 163810
rect 249634 163144 250294 163810
rect 250462 163144 251122 163810
rect 251290 163144 251950 163810
rect 252118 163144 252778 163810
rect 252946 163144 253606 163810
rect 253774 163144 254434 163810
rect 254602 163144 255262 163810
rect 255430 163144 256090 163810
rect 256258 163144 256918 163810
rect 257086 163144 257746 163810
rect 257914 163144 258574 163810
rect 258742 163144 259402 163810
rect 259570 163144 260230 163810
rect 260398 163144 261058 163810
rect 261226 163144 261886 163810
rect 262054 163144 262714 163810
rect 262882 163144 263542 163810
rect 263710 163144 264370 163810
rect 264538 163144 265198 163810
rect 265366 163144 266026 163810
rect 266194 163144 266854 163810
rect 267022 163144 267682 163810
rect 267850 163144 268510 163810
rect 268678 163144 269338 163810
rect 269506 163144 270166 163810
rect 270334 163144 270994 163810
rect 271162 163144 271822 163810
rect 271990 163144 272650 163810
rect 272818 163144 273478 163810
rect 273646 163144 274306 163810
rect 274474 163144 275134 163810
rect 275302 163144 275962 163810
rect 276130 163144 276790 163810
rect 276958 163144 277618 163810
rect 277786 163144 278446 163810
rect 278614 163144 279274 163810
rect 279442 163144 280102 163810
rect 280270 163144 280930 163810
rect 281098 163144 281758 163810
rect 281926 163144 282586 163810
rect 282754 163144 283414 163810
rect 283582 163144 284242 163810
rect 284410 163144 285070 163810
rect 285238 163144 285898 163810
rect 286066 163144 286726 163810
rect 286894 163144 287554 163810
rect 287722 163144 288382 163810
rect 288550 163144 289210 163810
rect 289378 163144 290038 163810
rect 290206 163144 290866 163810
rect 291034 163144 291694 163810
rect 291862 163144 292522 163810
rect 292690 163144 293350 163810
rect 293518 163144 294178 163810
rect 294346 163144 295006 163810
rect 295174 163144 295834 163810
rect 296002 163144 296662 163810
rect 296830 163144 297490 163810
rect 297658 163144 298318 163810
rect 298486 163144 299146 163810
rect 299314 163144 299974 163810
rect 300142 163144 300802 163810
rect 300970 163144 301630 163810
rect 301798 163144 302458 163810
rect 302626 163144 303286 163810
rect 303454 163144 304114 163810
rect 304282 163144 304942 163810
rect 305110 163144 305770 163810
rect 305938 163144 306598 163810
rect 306766 163144 307426 163810
rect 307594 163144 308254 163810
rect 308422 163144 309082 163810
rect 309250 163144 309910 163810
rect 310078 163144 310738 163810
rect 310906 163144 311566 163810
rect 311734 163144 312394 163810
rect 312562 163144 313222 163810
rect 313390 163144 314050 163810
rect 314218 163144 314878 163810
rect 315046 163144 315706 163810
rect 315874 163144 316534 163810
rect 316702 163144 317362 163810
rect 317530 163144 318190 163810
rect 318358 163144 319018 163810
rect 319186 163144 319846 163810
rect 320014 163144 320674 163810
rect 320842 163144 321502 163810
rect 321670 163144 322330 163810
rect 322498 163144 323158 163810
rect 323326 163144 323986 163810
rect 324154 163144 324814 163810
rect 324982 163144 325642 163810
rect 325810 163144 326470 163810
rect 326638 163144 327298 163810
rect 327466 163144 328126 163810
rect 328294 163144 328954 163810
rect 329122 163144 329782 163810
rect 329950 163144 330610 163810
rect 330778 163144 331438 163810
rect 331606 163144 332266 163810
rect 332434 163144 333094 163810
rect 333262 163144 333922 163810
rect 334090 163144 334750 163810
rect 334918 163144 335578 163810
rect 335746 163144 336406 163810
rect 336574 163144 337234 163810
rect 337402 163144 338062 163810
rect 338230 163144 338890 163810
rect 339058 163144 339718 163810
rect 339886 163144 340546 163810
rect 340714 163144 341374 163810
rect 341542 163144 342202 163810
rect 342370 163144 343030 163810
rect 343198 163144 343858 163810
rect 344026 163144 344686 163810
rect 344854 163144 345514 163810
rect 345682 163144 346342 163810
rect 346510 163144 347170 163810
rect 347338 163144 347998 163810
rect 348166 163144 348826 163810
rect 348994 163144 349654 163810
rect 349822 163144 350482 163810
rect 350650 163144 351310 163810
rect 351478 163144 352138 163810
rect 352306 163144 352966 163810
rect 353134 163144 353794 163810
rect 353962 163144 354622 163810
rect 354790 163144 355450 163810
rect 355618 163144 356278 163810
rect 356446 163144 357106 163810
rect 357274 163144 357934 163810
rect 358102 163144 358762 163810
rect 358930 163144 359590 163810
rect 359758 163144 360418 163810
rect 360586 163144 361246 163810
rect 361414 163144 362074 163810
rect 362242 163144 362902 163810
rect 363070 163144 363730 163810
rect 363898 163144 364558 163810
rect 364726 163144 365386 163810
rect 365554 163144 366214 163810
rect 366382 163144 367042 163810
rect 367210 163144 367870 163810
rect 368038 163144 368698 163810
rect 368866 163144 369526 163810
rect 369694 163144 370354 163810
rect 370522 163144 371182 163810
rect 371350 163144 372010 163810
rect 372178 163144 372838 163810
rect 373006 163144 373666 163810
rect 373834 163144 374494 163810
rect 374662 163144 375322 163810
rect 375490 163144 376150 163810
rect 376318 163144 376978 163810
rect 377146 163144 377806 163810
rect 377974 163144 378634 163810
rect 378802 163144 379462 163810
rect 379630 163144 380290 163810
rect 380458 163144 381118 163810
rect 381286 163144 381946 163810
rect 382114 163144 382774 163810
rect 382942 163144 383602 163810
rect 383770 163144 384430 163810
rect 384598 163144 385258 163810
rect 385426 163144 386086 163810
rect 386254 163144 386914 163810
rect 387082 163144 387742 163810
rect 387910 163144 388570 163810
rect 388738 163144 389398 163810
rect 389566 163144 390226 163810
rect 390394 163144 391054 163810
rect 391222 163144 391882 163810
rect 392050 163144 392710 163810
rect 392878 163144 393538 163810
rect 393706 163144 394366 163810
rect 394534 163144 395194 163810
rect 395362 163144 396022 163810
rect 396190 163144 396850 163810
rect 397018 163144 397678 163810
rect 397846 163144 398506 163810
rect 398674 163144 399334 163810
rect 399502 163144 400162 163810
rect 400330 163144 400990 163810
rect 401158 163144 401818 163810
rect 401986 163144 402646 163810
rect 402814 163144 403474 163810
rect 403642 163144 404302 163810
rect 404470 163144 405130 163810
rect 405298 163144 405958 163810
rect 406126 163144 406786 163810
rect 406954 163144 407614 163810
rect 407782 163144 408442 163810
rect 408610 163144 409270 163810
rect 409438 163144 410098 163810
rect 410266 163144 410926 163810
rect 411094 163144 411754 163810
rect 411922 163144 412582 163810
rect 412750 163144 413410 163810
rect 413578 163144 414238 163810
rect 414406 163144 415066 163810
rect 415234 163144 415894 163810
rect 416062 163144 416722 163810
rect 416890 163144 417550 163810
rect 417718 163144 418378 163810
rect 418546 163144 419206 163810
rect 419374 163144 420034 163810
rect 420202 163144 420862 163810
rect 421030 163144 421690 163810
rect 421858 163144 422518 163810
rect 422686 163144 423346 163810
rect 423514 163144 424174 163810
rect 424342 163144 425002 163810
rect 425170 163144 425830 163810
rect 425998 163144 426658 163810
rect 426826 163144 427486 163810
rect 427654 163144 428314 163810
rect 428482 163144 429142 163810
rect 429310 163144 429970 163810
rect 430138 163144 430798 163810
rect 430966 163144 431626 163810
rect 431794 163144 432454 163810
rect 432622 163144 433282 163810
rect 433450 163144 434110 163810
rect 434278 163144 434938 163810
rect 435106 163144 435766 163810
rect 435934 163144 436594 163810
rect 436762 163144 437422 163810
rect 437590 163144 438250 163810
rect 438418 163144 439078 163810
rect 439246 163144 439906 163810
rect 440074 163144 440734 163810
rect 440902 163144 441562 163810
rect 441730 163144 442390 163810
rect 442558 163144 443218 163810
rect 443386 163144 444046 163810
rect 444214 163144 444874 163810
rect 445042 163144 445702 163810
rect 445870 163144 446530 163810
rect 446698 163144 447358 163810
rect 447526 163144 448186 163810
rect 448354 163144 449014 163810
rect 449182 163144 449842 163810
rect 450010 163144 450670 163810
rect 450838 163144 451498 163810
rect 451666 163144 452326 163810
rect 452494 163144 453154 163810
rect 453322 163144 453982 163810
rect 454150 163144 454810 163810
rect 454978 163144 455638 163810
rect 455806 163144 456466 163810
rect 456634 163144 457294 163810
rect 457462 163144 458122 163810
rect 458290 163144 458950 163810
rect 459118 163144 459778 163810
rect 459946 163144 460606 163810
rect 460774 163144 461434 163810
rect 461602 163144 462262 163810
rect 462430 163144 463090 163810
rect 463258 163144 463918 163810
rect 464086 163144 464746 163810
rect 464914 163144 465574 163810
rect 465742 163144 466402 163810
rect 466570 163144 467230 163810
rect 467398 163144 468058 163810
rect 468226 163144 468886 163810
rect 469054 163144 469714 163810
rect 469882 163144 470542 163810
rect 470710 163144 471370 163810
rect 471538 163144 472198 163810
rect 472366 163144 473026 163810
rect 473194 163144 473854 163810
rect 474022 163144 474682 163810
rect 474850 163144 475510 163810
rect 475678 163144 476338 163810
rect 476506 163144 477166 163810
rect 477334 163144 477994 163810
rect 478162 163144 478822 163810
rect 478990 163144 479650 163810
rect 479818 163144 480478 163810
rect 480646 163144 481306 163810
rect 481474 163144 482134 163810
rect 482302 163144 482962 163810
rect 483130 163144 483790 163810
rect 483958 163144 484618 163810
rect 484786 163144 485446 163810
rect 485614 163144 486274 163810
rect 486442 163144 487102 163810
rect 487270 163144 487930 163810
rect 488098 163144 488758 163810
rect 488926 163144 489586 163810
rect 489754 163144 490414 163810
rect 490582 163144 491242 163810
rect 491410 163144 492070 163810
rect 492238 163144 492898 163810
rect 493066 163144 493726 163810
rect 493894 163144 494554 163810
rect 494722 163144 495382 163810
rect 495550 163144 496210 163810
rect 496378 163144 497038 163810
rect 497206 163144 497866 163810
rect 498034 163144 498694 163810
rect 498862 163144 499522 163810
rect 499690 163144 500350 163810
rect 500518 163144 501178 163810
rect 501346 163144 502006 163810
rect 502174 163144 502834 163810
rect 503002 163144 503662 163810
rect 503830 163144 504490 163810
rect 504658 163144 505318 163810
rect 505486 163144 506146 163810
rect 506314 163144 506974 163810
rect 507142 163144 507802 163810
rect 507970 163144 508630 163810
rect 508798 163144 509458 163810
rect 509626 163144 510286 163810
rect 510454 163144 511114 163810
rect 511282 163144 511942 163810
rect 512110 163144 512770 163810
rect 512938 163144 513598 163810
rect 513766 163144 514426 163810
rect 514594 163144 515254 163810
rect 515422 163144 516082 163810
rect 516250 163144 516910 163810
rect 517078 163144 517738 163810
rect 517906 163144 518566 163810
rect 518734 163144 519394 163810
rect 519562 163144 520222 163810
rect 520390 163144 521622 163810
rect 2870 856 521622 163144
rect 2870 748 253916 856
rect 254084 748 255916 856
rect 256084 748 257916 856
rect 258084 748 259916 856
rect 260084 748 261916 856
rect 262084 748 263916 856
rect 264084 748 265916 856
rect 266084 748 491916 856
rect 492084 748 493916 856
rect 494084 748 495916 856
rect 496084 748 497916 856
rect 498084 748 499916 856
rect 500084 748 501916 856
rect 502084 748 521622 856
<< metal3 >>
rect 523200 161304 524000 161424
rect 523200 159128 524000 159248
rect 523200 156952 524000 157072
rect 523200 154776 524000 154896
rect 523200 152600 524000 152720
rect 523200 150424 524000 150544
rect 523200 148248 524000 148368
rect 523200 146072 524000 146192
rect 523200 143896 524000 144016
rect 0 143352 800 143472
rect 523200 141720 524000 141840
rect 0 141352 800 141472
rect 0 139352 800 139472
rect 523200 139544 524000 139664
rect 0 137352 800 137472
rect 523200 137368 524000 137488
rect 523200 135192 524000 135312
rect 523200 133016 524000 133136
rect 523200 130840 524000 130960
rect 523200 128664 524000 128784
rect 523200 126488 524000 126608
rect 523200 124312 524000 124432
rect 523200 122136 524000 122256
rect 523200 119960 524000 120080
rect 523200 117784 524000 117904
rect 523200 115608 524000 115728
rect 523200 113432 524000 113552
rect 523200 111256 524000 111376
rect 523200 109080 524000 109200
rect 523200 106904 524000 107024
rect 523200 104728 524000 104848
rect 523200 102552 524000 102672
rect 523200 100376 524000 100496
rect 523200 98200 524000 98320
rect 523200 96024 524000 96144
rect 523200 93848 524000 93968
rect 523200 91672 524000 91792
rect 523200 89496 524000 89616
rect 523200 87320 524000 87440
rect 523200 85144 524000 85264
rect 523200 82968 524000 83088
rect 523200 80792 524000 80912
rect 523200 78616 524000 78736
rect 523200 76440 524000 76560
rect 523200 74264 524000 74384
rect 523200 72088 524000 72208
rect 523200 69912 524000 70032
rect 523200 67736 524000 67856
rect 523200 65560 524000 65680
rect 523200 63384 524000 63504
rect 523200 61208 524000 61328
rect 523200 59032 524000 59152
rect 523200 56856 524000 56976
rect 523200 54680 524000 54800
rect 523200 52504 524000 52624
rect 523200 50328 524000 50448
rect 523200 48152 524000 48272
rect 523200 45976 524000 46096
rect 523200 43800 524000 43920
rect 523200 41624 524000 41744
rect 523200 39448 524000 39568
rect 523200 37272 524000 37392
rect 523200 35096 524000 35216
rect 523200 32920 524000 33040
rect 523200 30744 524000 30864
rect 523200 28568 524000 28688
rect 523200 26392 524000 26512
rect 523200 24216 524000 24336
rect 523200 22040 524000 22160
rect 523200 19864 524000 19984
rect 523200 17688 524000 17808
rect 523200 15512 524000 15632
rect 523200 13336 524000 13456
rect 523200 11160 524000 11280
rect 523200 8984 524000 9104
rect 523200 6808 524000 6928
rect 523200 4632 524000 4752
rect 523200 2456 524000 2576
<< obsm3 >>
rect 644 161504 523200 163709
rect 644 161224 523120 161504
rect 644 159328 523200 161224
rect 644 159048 523120 159328
rect 644 157152 523200 159048
rect 644 156872 523120 157152
rect 644 154976 523200 156872
rect 644 154696 523120 154976
rect 644 152800 523200 154696
rect 644 152520 523120 152800
rect 644 150624 523200 152520
rect 644 150344 523120 150624
rect 644 148448 523200 150344
rect 644 148168 523120 148448
rect 644 146272 523200 148168
rect 644 145992 523120 146272
rect 644 144096 523200 145992
rect 644 143816 523120 144096
rect 644 143552 523200 143816
rect 880 143272 523200 143552
rect 644 141920 523200 143272
rect 644 141640 523120 141920
rect 644 141552 523200 141640
rect 880 141272 523200 141552
rect 644 139744 523200 141272
rect 644 139552 523120 139744
rect 880 139464 523120 139552
rect 880 139272 523200 139464
rect 644 137568 523200 139272
rect 644 137552 523120 137568
rect 880 137288 523120 137552
rect 880 137272 523200 137288
rect 644 135392 523200 137272
rect 644 135112 523120 135392
rect 644 133216 523200 135112
rect 644 132936 523120 133216
rect 644 131040 523200 132936
rect 644 130760 523120 131040
rect 644 128864 523200 130760
rect 644 128584 523120 128864
rect 644 126688 523200 128584
rect 644 126408 523120 126688
rect 644 124512 523200 126408
rect 644 124232 523120 124512
rect 644 122336 523200 124232
rect 644 122056 523120 122336
rect 644 120160 523200 122056
rect 644 119880 523120 120160
rect 644 117984 523200 119880
rect 644 117704 523120 117984
rect 644 115808 523200 117704
rect 644 115528 523120 115808
rect 644 113632 523200 115528
rect 644 113352 523120 113632
rect 644 111456 523200 113352
rect 644 111176 523120 111456
rect 644 109280 523200 111176
rect 644 109000 523120 109280
rect 644 107104 523200 109000
rect 644 106824 523120 107104
rect 644 104928 523200 106824
rect 644 104648 523120 104928
rect 644 102752 523200 104648
rect 644 102472 523120 102752
rect 644 100576 523200 102472
rect 644 100296 523120 100576
rect 644 98400 523200 100296
rect 644 98120 523120 98400
rect 644 96224 523200 98120
rect 644 95944 523120 96224
rect 644 94048 523200 95944
rect 644 93768 523120 94048
rect 644 91872 523200 93768
rect 644 91592 523120 91872
rect 644 89696 523200 91592
rect 644 89416 523120 89696
rect 644 87520 523200 89416
rect 644 87240 523120 87520
rect 644 85344 523200 87240
rect 644 85064 523120 85344
rect 644 83168 523200 85064
rect 644 82888 523120 83168
rect 644 80992 523200 82888
rect 644 80712 523120 80992
rect 644 78816 523200 80712
rect 644 78536 523120 78816
rect 644 76640 523200 78536
rect 644 76360 523120 76640
rect 644 74464 523200 76360
rect 644 74184 523120 74464
rect 644 72288 523200 74184
rect 644 72008 523120 72288
rect 644 70112 523200 72008
rect 644 69832 523120 70112
rect 644 67936 523200 69832
rect 644 67656 523120 67936
rect 644 65760 523200 67656
rect 644 65480 523120 65760
rect 644 63584 523200 65480
rect 644 63304 523120 63584
rect 644 61408 523200 63304
rect 644 61128 523120 61408
rect 644 59232 523200 61128
rect 644 58952 523120 59232
rect 644 57056 523200 58952
rect 644 56776 523120 57056
rect 644 54880 523200 56776
rect 644 54600 523120 54880
rect 644 52704 523200 54600
rect 644 52424 523120 52704
rect 644 50528 523200 52424
rect 644 50248 523120 50528
rect 644 48352 523200 50248
rect 644 48072 523120 48352
rect 644 46176 523200 48072
rect 644 45896 523120 46176
rect 644 44000 523200 45896
rect 644 43720 523120 44000
rect 644 41824 523200 43720
rect 644 41544 523120 41824
rect 644 39648 523200 41544
rect 644 39368 523120 39648
rect 644 37472 523200 39368
rect 644 37192 523120 37472
rect 644 35296 523200 37192
rect 644 35016 523120 35296
rect 644 33120 523200 35016
rect 644 32840 523120 33120
rect 644 30944 523200 32840
rect 644 30664 523120 30944
rect 644 28768 523200 30664
rect 644 28488 523120 28768
rect 644 26592 523200 28488
rect 644 26312 523120 26592
rect 644 24416 523200 26312
rect 644 24136 523120 24416
rect 644 22240 523200 24136
rect 644 21960 523120 22240
rect 644 20064 523200 21960
rect 644 19784 523120 20064
rect 644 17888 523200 19784
rect 644 17608 523120 17888
rect 644 15712 523200 17608
rect 644 15432 523120 15712
rect 644 13536 523200 15432
rect 644 13256 523120 13536
rect 644 11360 523200 13256
rect 644 11080 523120 11360
rect 644 9184 523200 11080
rect 644 8904 523120 9184
rect 644 7008 523200 8904
rect 644 6728 523120 7008
rect 644 4832 523200 6728
rect 644 4552 523120 4832
rect 644 2656 523200 4552
rect 644 2483 523120 2656
<< metal4 >>
rect -156 540 164 163204
rect 504 1200 824 162544
rect 5128 540 5448 163204
rect 7448 540 7768 163204
rect 15128 117017 15448 163204
rect 17448 117017 17768 163204
rect 25128 117017 25448 163204
rect 27448 117017 27768 163204
rect 35128 117017 35448 163204
rect 37448 117017 37768 163204
rect 45128 119820 45448 163204
rect 47448 117017 47768 163204
rect 55128 117017 55448 163204
rect 57448 117017 57768 163204
rect 65128 117017 65448 163204
rect 67448 117017 67768 163204
rect 75128 119820 75448 163204
rect 77448 117017 77768 163204
rect 85128 117017 85448 163204
rect 87448 117017 87768 163204
rect 95128 117017 95448 163204
rect 97448 117017 97768 163204
rect 105128 117017 105448 163204
rect 107448 117017 107768 163204
rect 115128 117017 115448 163204
rect 117448 117017 117768 163204
rect 125128 117017 125448 163204
rect 127448 117017 127768 163204
rect 135128 117017 135448 163204
rect 137448 117017 137768 163204
rect 145128 117017 145448 163204
rect 147448 117017 147768 163204
rect 15128 540 15448 14367
rect 17448 540 17768 14367
rect 25128 540 25448 14367
rect 27448 540 27768 14367
rect 35128 540 35448 14367
rect 37448 540 37768 14367
rect 45128 540 45448 10068
rect 47448 540 47768 14367
rect 55128 540 55448 14367
rect 57448 540 57768 14367
rect 65128 540 65448 14367
rect 67448 540 67768 14367
rect 75128 540 75448 10068
rect 77448 540 77768 14367
rect 85128 540 85448 14367
rect 87448 540 87768 14367
rect 95128 540 95448 14367
rect 97448 540 97768 14367
rect 105128 540 105448 14367
rect 107448 540 107768 14367
rect 115128 540 115448 14367
rect 117448 540 117768 14367
rect 125128 540 125448 14367
rect 127448 540 127768 14367
rect 135128 540 135448 14367
rect 137448 540 137768 14367
rect 145128 540 145448 14367
rect 147448 540 147768 14367
rect 155128 540 155448 163204
rect 157448 540 157768 163204
rect 165128 540 165448 163204
rect 167448 119820 167768 163204
rect 167448 540 167768 10068
rect 175128 540 175448 163204
rect 177448 540 177768 163204
rect 185128 540 185448 163204
rect 187448 540 187768 163204
rect 195128 540 195448 163204
rect 197448 540 197768 163204
rect 205128 540 205448 163204
rect 207448 540 207768 163204
rect 215128 540 215448 163204
rect 217448 540 217768 163204
rect 225128 540 225448 163204
rect 227448 540 227768 163204
rect 235128 540 235448 163204
rect 237448 540 237768 163204
rect 245128 540 245448 163204
rect 247448 540 247768 163204
rect 255128 540 255448 163204
rect 257448 540 257768 163204
rect 265128 540 265448 163204
rect 267448 540 267768 163204
rect 275128 540 275448 163204
rect 277448 540 277768 163204
rect 285128 540 285448 163204
rect 287448 540 287768 163204
rect 295128 540 295448 163204
rect 297448 540 297768 163204
rect 305128 540 305448 163204
rect 307448 540 307768 163204
rect 315128 540 315448 163204
rect 317448 540 317768 163204
rect 325128 540 325448 163204
rect 327448 540 327768 163204
rect 335128 540 335448 163204
rect 337448 540 337768 163204
rect 345128 540 345448 163204
rect 347448 540 347768 163204
rect 355128 540 355448 163204
rect 357448 540 357768 163204
rect 365128 540 365448 163204
rect 367448 540 367768 163204
rect 375128 540 375448 163204
rect 377448 540 377768 163204
rect 385128 540 385448 163204
rect 387448 540 387768 163204
rect 395128 540 395448 163204
rect 397448 540 397768 163204
rect 405128 540 405448 163204
rect 407448 540 407768 163204
rect 415128 98793 415448 163204
rect 417448 98793 417768 163204
rect 425128 99692 425448 163204
rect 427448 98793 427768 163204
rect 435128 98793 435448 163204
rect 437448 98793 437768 163204
rect 445128 98793 445448 163204
rect 447448 98793 447768 163204
rect 455128 98793 455448 163204
rect 457448 98793 457768 163204
rect 465128 98793 465448 163204
rect 467448 98793 467768 163204
rect 475128 98793 475448 163204
rect 477448 98793 477768 163204
rect 485128 98793 485448 163204
rect 487448 98793 487768 163204
rect 495128 98793 495448 163204
rect 497448 98793 497768 163204
rect 415128 540 415448 14775
rect 417448 540 417768 14775
rect 425128 540 425448 10068
rect 427448 540 427768 14775
rect 435128 540 435448 14775
rect 437448 540 437768 14775
rect 445128 540 445448 14775
rect 447448 540 447768 14775
rect 455128 540 455448 14775
rect 457448 540 457768 14775
rect 465128 540 465448 14775
rect 467448 540 467768 14775
rect 475128 540 475448 14775
rect 477448 540 477768 14775
rect 485128 540 485448 14775
rect 487448 540 487768 14775
rect 495128 540 495448 14775
rect 497448 540 497768 14775
rect 505128 540 505448 163204
rect 507448 540 507768 163204
rect 515128 540 515448 163204
rect 517448 540 517768 163204
rect 523116 1200 523436 162544
rect 523776 540 524096 163204
<< obsm4 >>
rect 13675 163284 514122 163709
rect 13675 116937 15048 163284
rect 15528 116937 17368 163284
rect 17848 116937 25048 163284
rect 25528 116937 27368 163284
rect 27848 116937 35048 163284
rect 35528 116937 37368 163284
rect 37848 119740 45048 163284
rect 45528 119740 47368 163284
rect 37848 116937 47368 119740
rect 47848 116937 55048 163284
rect 55528 116937 57368 163284
rect 57848 116937 65048 163284
rect 65528 116937 67368 163284
rect 67848 119740 75048 163284
rect 75528 119740 77368 163284
rect 67848 116937 77368 119740
rect 77848 116937 85048 163284
rect 85528 116937 87368 163284
rect 87848 116937 95048 163284
rect 95528 116937 97368 163284
rect 97848 116937 105048 163284
rect 105528 116937 107368 163284
rect 107848 116937 115048 163284
rect 115528 116937 117368 163284
rect 117848 116937 125048 163284
rect 125528 116937 127368 163284
rect 127848 116937 135048 163284
rect 135528 116937 137368 163284
rect 137848 116937 145048 163284
rect 145528 116937 147368 163284
rect 147848 116937 155048 163284
rect 13675 14447 155048 116937
rect 13675 5203 15048 14447
rect 15528 5203 17368 14447
rect 17848 5203 25048 14447
rect 25528 5203 27368 14447
rect 27848 5203 35048 14447
rect 35528 5203 37368 14447
rect 37848 10148 47368 14447
rect 37848 5203 45048 10148
rect 45528 5203 47368 10148
rect 47848 5203 55048 14447
rect 55528 5203 57368 14447
rect 57848 5203 65048 14447
rect 65528 5203 67368 14447
rect 67848 10148 77368 14447
rect 67848 5203 75048 10148
rect 75528 5203 77368 10148
rect 77848 5203 85048 14447
rect 85528 5203 87368 14447
rect 87848 5203 95048 14447
rect 95528 5203 97368 14447
rect 97848 5203 105048 14447
rect 105528 5203 107368 14447
rect 107848 5203 115048 14447
rect 115528 5203 117368 14447
rect 117848 5203 125048 14447
rect 125528 5203 127368 14447
rect 127848 5203 135048 14447
rect 135528 5203 137368 14447
rect 137848 5203 145048 14447
rect 145528 5203 147368 14447
rect 147848 5203 155048 14447
rect 155528 5203 157368 163284
rect 157848 5203 165048 163284
rect 165528 119740 167368 163284
rect 167848 119740 175048 163284
rect 165528 10148 175048 119740
rect 165528 5203 167368 10148
rect 167848 5203 175048 10148
rect 175528 5203 177368 163284
rect 177848 5203 185048 163284
rect 185528 5203 187368 163284
rect 187848 5203 195048 163284
rect 195528 5203 197368 163284
rect 197848 5203 205048 163284
rect 205528 5203 207368 163284
rect 207848 5203 215048 163284
rect 215528 5203 217368 163284
rect 217848 5203 225048 163284
rect 225528 5203 227368 163284
rect 227848 5203 235048 163284
rect 235528 5203 237368 163284
rect 237848 5203 245048 163284
rect 245528 5203 247368 163284
rect 247848 5203 255048 163284
rect 255528 5203 257368 163284
rect 257848 5203 265048 163284
rect 265528 5203 267368 163284
rect 267848 5203 275048 163284
rect 275528 5203 277368 163284
rect 277848 5203 285048 163284
rect 285528 5203 287368 163284
rect 287848 5203 295048 163284
rect 295528 5203 297368 163284
rect 297848 5203 305048 163284
rect 305528 5203 307368 163284
rect 307848 5203 315048 163284
rect 315528 5203 317368 163284
rect 317848 5203 325048 163284
rect 325528 5203 327368 163284
rect 327848 5203 335048 163284
rect 335528 5203 337368 163284
rect 337848 5203 345048 163284
rect 345528 5203 347368 163284
rect 347848 5203 355048 163284
rect 355528 5203 357368 163284
rect 357848 5203 365048 163284
rect 365528 5203 367368 163284
rect 367848 5203 375048 163284
rect 375528 5203 377368 163284
rect 377848 5203 385048 163284
rect 385528 5203 387368 163284
rect 387848 5203 395048 163284
rect 395528 5203 397368 163284
rect 397848 5203 405048 163284
rect 405528 5203 407368 163284
rect 407848 98713 415048 163284
rect 415528 98713 417368 163284
rect 417848 99612 425048 163284
rect 425528 99612 427368 163284
rect 417848 98713 427368 99612
rect 427848 98713 435048 163284
rect 435528 98713 437368 163284
rect 437848 98713 445048 163284
rect 445528 98713 447368 163284
rect 447848 98713 455048 163284
rect 455528 98713 457368 163284
rect 457848 98713 465048 163284
rect 465528 98713 467368 163284
rect 467848 98713 475048 163284
rect 475528 98713 477368 163284
rect 477848 98713 485048 163284
rect 485528 98713 487368 163284
rect 487848 98713 495048 163284
rect 495528 98713 497368 163284
rect 497848 98713 505048 163284
rect 407848 14855 505048 98713
rect 407848 5203 415048 14855
rect 415528 5203 417368 14855
rect 417848 10148 427368 14855
rect 417848 5203 425048 10148
rect 425528 5203 427368 10148
rect 427848 5203 435048 14855
rect 435528 5203 437368 14855
rect 437848 5203 445048 14855
rect 445528 5203 447368 14855
rect 447848 5203 455048 14855
rect 455528 5203 457368 14855
rect 457848 5203 465048 14855
rect 465528 5203 467368 14855
rect 467848 5203 475048 14855
rect 475528 5203 477368 14855
rect 477848 5203 485048 14855
rect 485528 5203 487368 14855
rect 487848 5203 495048 14855
rect 495528 5203 497368 14855
rect 497848 5203 505048 14855
rect 505528 5203 507368 163284
rect 507848 5203 514122 163284
<< metal5 >>
rect -156 162884 524096 163204
rect 504 162224 523436 162544
rect -156 158210 524096 158530
rect -156 155890 524096 156210
rect -156 148210 524096 148530
rect -156 145890 524096 146210
rect -156 138210 524096 138530
rect -156 135890 524096 136210
rect -156 128210 524096 128530
rect -156 125890 524096 126210
rect -156 118210 524096 118530
rect -156 115890 524096 116210
rect -156 108210 524096 108530
rect -156 105890 524096 106210
rect -156 98210 524096 98530
rect -156 95890 524096 96210
rect -156 88210 524096 88530
rect -156 85890 524096 86210
rect -156 78210 524096 78530
rect -156 75890 524096 76210
rect -156 68210 524096 68530
rect -156 65890 524096 66210
rect -156 58210 524096 58530
rect -156 55890 524096 56210
rect -156 48210 524096 48530
rect -156 45890 524096 46210
rect -156 38210 524096 38530
rect -156 35890 524096 36210
rect -156 28210 524096 28530
rect -156 25890 524096 26210
rect -156 18210 524096 18530
rect -156 15890 524096 16210
rect -156 8210 524096 8530
rect -156 5890 524096 6210
rect 504 1200 523436 1520
rect -156 540 524096 860
<< obsm5 >>
rect 88620 158850 514164 161660
rect 88620 156530 514164 157890
rect 88620 148850 514164 155570
rect 88620 146530 514164 147890
rect 88620 138850 514164 145570
rect 88620 136530 514164 137890
rect 88620 128850 514164 135570
rect 88620 126530 514164 127890
rect 88620 118850 514164 125570
rect 88620 116530 514164 117890
rect 88620 108850 514164 115570
rect 88620 106530 514164 107890
rect 88620 98850 514164 105570
rect 88620 96530 514164 97890
rect 88620 88850 514164 95570
rect 88620 86530 514164 87890
rect 88620 78850 514164 85570
rect 88620 76530 514164 77890
rect 88620 68850 514164 75570
rect 88620 66530 514164 67890
rect 88620 58850 514164 65570
rect 88620 56530 514164 57890
rect 88620 49820 514164 55570
<< labels >>
rlabel metal4 s -156 540 164 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -156 540 524096 860 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -156 162884 524096 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 523776 540 524096 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 7448 540 7768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 17448 540 17768 14367 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 17448 117017 17768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 27448 540 27768 14367 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 27448 117017 27768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 37448 540 37768 14367 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 37448 117017 37768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47448 540 47768 14367 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47448 117017 47768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 57448 540 57768 14367 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 57448 117017 57768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 67448 540 67768 14367 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 67448 117017 67768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 77448 540 77768 14367 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 77448 117017 77768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 87448 540 87768 14367 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 87448 117017 87768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 97448 540 97768 14367 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 97448 117017 97768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 107448 540 107768 14367 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 107448 117017 107768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 117448 540 117768 14367 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 117448 117017 117768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127448 540 127768 14367 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127448 117017 127768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 137448 540 137768 14367 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 137448 117017 137768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 147448 540 147768 14367 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 147448 117017 147768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 157448 540 157768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 167448 540 167768 10068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 167448 119820 167768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 177448 540 177768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 187448 540 187768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 197448 540 197768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 207448 540 207768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 217448 540 217768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 227448 540 227768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 237448 540 237768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 247448 540 247768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 257448 540 257768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 267448 540 267768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 277448 540 277768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 287448 540 287768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 297448 540 297768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 307448 540 307768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 317448 540 317768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 327448 540 327768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 337448 540 337768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 347448 540 347768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 357448 540 357768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 367448 540 367768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 377448 540 377768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 387448 540 387768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 397448 540 397768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 407448 540 407768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 417448 540 417768 14775 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 417448 98793 417768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 427448 540 427768 14775 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 427448 98793 427768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 437448 540 437768 14775 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 437448 98793 437768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 447448 540 447768 14775 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 447448 98793 447768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 457448 540 457768 14775 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 457448 98793 457768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 467448 540 467768 14775 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 467448 98793 467768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 477448 540 477768 14775 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 477448 98793 477768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 487448 540 487768 14775 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 487448 98793 487768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 497448 540 497768 14775 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 497448 98793 497768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 507448 540 507768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 517448 540 517768 163204 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -156 8210 524096 8530 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -156 18210 524096 18530 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -156 28210 524096 28530 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -156 38210 524096 38530 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -156 48210 524096 48530 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -156 58210 524096 58530 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -156 68210 524096 68530 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -156 78210 524096 78530 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -156 88210 524096 88530 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -156 98210 524096 98530 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -156 108210 524096 108530 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -156 118210 524096 118530 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -156 128210 524096 128530 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -156 138210 524096 138530 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -156 148210 524096 148530 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -156 158210 524096 158530 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 504 1200 824 162544 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 504 1200 523436 1520 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 504 162224 523436 162544 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 523116 1200 523436 162544 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 5128 540 5448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 15128 540 15448 14367 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 15128 117017 15448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 25128 540 25448 14367 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 25128 117017 25448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 35128 540 35448 14367 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 35128 117017 35448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 45128 540 45448 10068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 45128 119820 45448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 55128 540 55448 14367 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 55128 117017 55448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 65128 540 65448 14367 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 65128 117017 65448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 75128 540 75448 10068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 75128 119820 75448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 85128 540 85448 14367 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 85128 117017 85448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 95128 540 95448 14367 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 95128 117017 95448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 105128 540 105448 14367 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 105128 117017 105448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 115128 540 115448 14367 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 115128 117017 115448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 125128 540 125448 14367 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 125128 117017 125448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 135128 540 135448 14367 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 135128 117017 135448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 145128 540 145448 14367 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 145128 117017 145448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 155128 540 155448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 165128 540 165448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 175128 540 175448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 185128 540 185448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 195128 540 195448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 205128 540 205448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 215128 540 215448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 225128 540 225448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 235128 540 235448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 245128 540 245448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 255128 540 255448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 265128 540 265448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 275128 540 275448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 285128 540 285448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 295128 540 295448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 305128 540 305448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 315128 540 315448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 325128 540 325448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 335128 540 335448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 345128 540 345448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 355128 540 355448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 365128 540 365448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 375128 540 375448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 385128 540 385448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 395128 540 395448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 405128 540 405448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 415128 540 415448 14775 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 415128 98793 415448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 425128 540 425448 10068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 425128 99692 425448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 435128 540 435448 14775 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 435128 98793 435448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 445128 540 445448 14775 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 445128 98793 445448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 455128 540 455448 14775 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 455128 98793 455448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 465128 540 465448 14775 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 465128 98793 465448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 475128 540 475448 14775 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 475128 98793 475448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 485128 540 485448 14775 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 485128 98793 485448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 495128 540 495448 14775 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 495128 98793 495448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 505128 540 505448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 515128 540 515448 163204 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -156 5890 524096 6210 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -156 15890 524096 16210 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -156 25890 524096 26210 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -156 35890 524096 36210 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -156 45890 524096 46210 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -156 55890 524096 56210 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -156 65890 524096 66210 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -156 75890 524096 76210 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -156 85890 524096 86210 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -156 95890 524096 96210 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -156 105890 524096 106210 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -156 115890 524096 116210 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -156 125890 524096 126210 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -156 135890 524096 136210 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -156 145890 524096 146210 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -156 155890 524096 156210 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 261972 0 262028 800 6 clk_in
port 3 nsew signal input
rlabel metal2 s 238758 163200 238814 164000 6 clk_out
port 4 nsew signal output
rlabel metal2 s 259972 0 260028 800 6 core_clk
port 5 nsew signal input
rlabel metal2 s 263972 0 264028 800 6 core_rstn
port 6 nsew signal input
rlabel metal3 s 523200 17688 524000 17808 6 debug_in
port 7 nsew signal input
rlabel metal3 s 523200 19864 524000 19984 6 debug_mode
port 8 nsew signal output
rlabel metal3 s 523200 22040 524000 22160 6 debug_oeb
port 9 nsew signal output
rlabel metal3 s 523200 24216 524000 24336 6 debug_out
port 10 nsew signal output
rlabel metal3 s 523200 135192 524000 135312 6 flash_clk
port 11 nsew signal output
rlabel metal3 s 523200 133016 524000 133136 6 flash_csb
port 12 nsew signal output
rlabel metal3 s 523200 137368 524000 137488 6 flash_io0_di
port 13 nsew signal input
rlabel metal3 s 523200 139544 524000 139664 6 flash_io0_do
port 14 nsew signal output
rlabel metal3 s 523200 141720 524000 141840 6 flash_io0_oeb
port 15 nsew signal output
rlabel metal3 s 523200 143896 524000 144016 6 flash_io1_di
port 16 nsew signal input
rlabel metal3 s 523200 146072 524000 146192 6 flash_io1_do
port 17 nsew signal output
rlabel metal3 s 523200 148248 524000 148368 6 flash_io1_oeb
port 18 nsew signal output
rlabel metal3 s 523200 150424 524000 150544 6 flash_io2_di
port 19 nsew signal input
rlabel metal3 s 523200 152600 524000 152720 6 flash_io2_do
port 20 nsew signal output
rlabel metal3 s 523200 154776 524000 154896 6 flash_io2_oeb
port 21 nsew signal output
rlabel metal3 s 523200 156952 524000 157072 6 flash_io3_di
port 22 nsew signal input
rlabel metal3 s 523200 159128 524000 159248 6 flash_io3_do
port 23 nsew signal output
rlabel metal3 s 523200 161304 524000 161424 6 flash_io3_oeb
port 24 nsew signal output
rlabel metal2 s 491972 0 492028 800 6 gpio_in_pad
port 25 nsew signal input
rlabel metal2 s 493972 0 494028 800 6 gpio_inenb_pad
port 26 nsew signal output
rlabel metal2 s 495972 0 496028 800 6 gpio_mode0_pad
port 27 nsew signal output
rlabel metal2 s 497972 0 498028 800 6 gpio_mode1_pad
port 28 nsew signal output
rlabel metal2 s 499972 0 500028 800 6 gpio_out_pad
port 29 nsew signal output
rlabel metal2 s 501972 0 502028 800 6 gpio_outenb_pad
port 30 nsew signal output
rlabel metal3 s 523200 56856 524000 56976 6 hk_ack_i
port 31 nsew signal input
rlabel metal3 s 523200 61208 524000 61328 6 hk_cyc_o
port 32 nsew signal output
rlabel metal3 s 523200 63384 524000 63504 6 hk_dat_i[0]
port 33 nsew signal input
rlabel metal3 s 523200 85144 524000 85264 6 hk_dat_i[10]
port 34 nsew signal input
rlabel metal3 s 523200 87320 524000 87440 6 hk_dat_i[11]
port 35 nsew signal input
rlabel metal3 s 523200 89496 524000 89616 6 hk_dat_i[12]
port 36 nsew signal input
rlabel metal3 s 523200 91672 524000 91792 6 hk_dat_i[13]
port 37 nsew signal input
rlabel metal3 s 523200 93848 524000 93968 6 hk_dat_i[14]
port 38 nsew signal input
rlabel metal3 s 523200 96024 524000 96144 6 hk_dat_i[15]
port 39 nsew signal input
rlabel metal3 s 523200 98200 524000 98320 6 hk_dat_i[16]
port 40 nsew signal input
rlabel metal3 s 523200 100376 524000 100496 6 hk_dat_i[17]
port 41 nsew signal input
rlabel metal3 s 523200 102552 524000 102672 6 hk_dat_i[18]
port 42 nsew signal input
rlabel metal3 s 523200 104728 524000 104848 6 hk_dat_i[19]
port 43 nsew signal input
rlabel metal3 s 523200 65560 524000 65680 6 hk_dat_i[1]
port 44 nsew signal input
rlabel metal3 s 523200 106904 524000 107024 6 hk_dat_i[20]
port 45 nsew signal input
rlabel metal3 s 523200 109080 524000 109200 6 hk_dat_i[21]
port 46 nsew signal input
rlabel metal3 s 523200 111256 524000 111376 6 hk_dat_i[22]
port 47 nsew signal input
rlabel metal3 s 523200 113432 524000 113552 6 hk_dat_i[23]
port 48 nsew signal input
rlabel metal3 s 523200 115608 524000 115728 6 hk_dat_i[24]
port 49 nsew signal input
rlabel metal3 s 523200 117784 524000 117904 6 hk_dat_i[25]
port 50 nsew signal input
rlabel metal3 s 523200 119960 524000 120080 6 hk_dat_i[26]
port 51 nsew signal input
rlabel metal3 s 523200 122136 524000 122256 6 hk_dat_i[27]
port 52 nsew signal input
rlabel metal3 s 523200 124312 524000 124432 6 hk_dat_i[28]
port 53 nsew signal input
rlabel metal3 s 523200 126488 524000 126608 6 hk_dat_i[29]
port 54 nsew signal input
rlabel metal3 s 523200 67736 524000 67856 6 hk_dat_i[2]
port 55 nsew signal input
rlabel metal3 s 523200 128664 524000 128784 6 hk_dat_i[30]
port 56 nsew signal input
rlabel metal3 s 523200 130840 524000 130960 6 hk_dat_i[31]
port 57 nsew signal input
rlabel metal3 s 523200 69912 524000 70032 6 hk_dat_i[3]
port 58 nsew signal input
rlabel metal3 s 523200 72088 524000 72208 6 hk_dat_i[4]
port 59 nsew signal input
rlabel metal3 s 523200 74264 524000 74384 6 hk_dat_i[5]
port 60 nsew signal input
rlabel metal3 s 523200 76440 524000 76560 6 hk_dat_i[6]
port 61 nsew signal input
rlabel metal3 s 523200 78616 524000 78736 6 hk_dat_i[7]
port 62 nsew signal input
rlabel metal3 s 523200 80792 524000 80912 6 hk_dat_i[8]
port 63 nsew signal input
rlabel metal3 s 523200 82968 524000 83088 6 hk_dat_i[9]
port 64 nsew signal input
rlabel metal3 s 523200 59032 524000 59152 6 hk_stb_o
port 65 nsew signal output
rlabel metal2 s 518622 163200 518678 164000 6 irq[0]
port 66 nsew signal input
rlabel metal2 s 519450 163200 519506 164000 6 irq[1]
port 67 nsew signal input
rlabel metal2 s 520278 163200 520334 164000 6 irq[2]
port 68 nsew signal input
rlabel metal3 s 523200 32920 524000 33040 6 irq[3]
port 69 nsew signal input
rlabel metal3 s 523200 30744 524000 30864 6 irq[4]
port 70 nsew signal input
rlabel metal3 s 523200 28568 524000 28688 6 irq[5]
port 71 nsew signal input
rlabel metal2 s 3606 163200 3662 164000 6 la_iena[0]
port 72 nsew signal output
rlabel metal2 s 336462 163200 336518 164000 6 la_iena[100]
port 73 nsew signal output
rlabel metal2 s 339774 163200 339830 164000 6 la_iena[101]
port 74 nsew signal output
rlabel metal2 s 343086 163200 343142 164000 6 la_iena[102]
port 75 nsew signal output
rlabel metal2 s 346398 163200 346454 164000 6 la_iena[103]
port 76 nsew signal output
rlabel metal2 s 349710 163200 349766 164000 6 la_iena[104]
port 77 nsew signal output
rlabel metal2 s 353022 163200 353078 164000 6 la_iena[105]
port 78 nsew signal output
rlabel metal2 s 356334 163200 356390 164000 6 la_iena[106]
port 79 nsew signal output
rlabel metal2 s 359646 163200 359702 164000 6 la_iena[107]
port 80 nsew signal output
rlabel metal2 s 362958 163200 363014 164000 6 la_iena[108]
port 81 nsew signal output
rlabel metal2 s 366270 163200 366326 164000 6 la_iena[109]
port 82 nsew signal output
rlabel metal2 s 36726 163200 36782 164000 6 la_iena[10]
port 83 nsew signal output
rlabel metal2 s 369582 163200 369638 164000 6 la_iena[110]
port 84 nsew signal output
rlabel metal2 s 372894 163200 372950 164000 6 la_iena[111]
port 85 nsew signal output
rlabel metal2 s 376206 163200 376262 164000 6 la_iena[112]
port 86 nsew signal output
rlabel metal2 s 379518 163200 379574 164000 6 la_iena[113]
port 87 nsew signal output
rlabel metal2 s 382830 163200 382886 164000 6 la_iena[114]
port 88 nsew signal output
rlabel metal2 s 386142 163200 386198 164000 6 la_iena[115]
port 89 nsew signal output
rlabel metal2 s 389454 163200 389510 164000 6 la_iena[116]
port 90 nsew signal output
rlabel metal2 s 392766 163200 392822 164000 6 la_iena[117]
port 91 nsew signal output
rlabel metal2 s 396078 163200 396134 164000 6 la_iena[118]
port 92 nsew signal output
rlabel metal2 s 399390 163200 399446 164000 6 la_iena[119]
port 93 nsew signal output
rlabel metal2 s 40038 163200 40094 164000 6 la_iena[11]
port 94 nsew signal output
rlabel metal2 s 402702 163200 402758 164000 6 la_iena[120]
port 95 nsew signal output
rlabel metal2 s 406014 163200 406070 164000 6 la_iena[121]
port 96 nsew signal output
rlabel metal2 s 409326 163200 409382 164000 6 la_iena[122]
port 97 nsew signal output
rlabel metal2 s 412638 163200 412694 164000 6 la_iena[123]
port 98 nsew signal output
rlabel metal2 s 415950 163200 416006 164000 6 la_iena[124]
port 99 nsew signal output
rlabel metal2 s 419262 163200 419318 164000 6 la_iena[125]
port 100 nsew signal output
rlabel metal2 s 422574 163200 422630 164000 6 la_iena[126]
port 101 nsew signal output
rlabel metal2 s 425886 163200 425942 164000 6 la_iena[127]
port 102 nsew signal output
rlabel metal2 s 43350 163200 43406 164000 6 la_iena[12]
port 103 nsew signal output
rlabel metal2 s 46662 163200 46718 164000 6 la_iena[13]
port 104 nsew signal output
rlabel metal2 s 49974 163200 50030 164000 6 la_iena[14]
port 105 nsew signal output
rlabel metal2 s 53286 163200 53342 164000 6 la_iena[15]
port 106 nsew signal output
rlabel metal2 s 56598 163200 56654 164000 6 la_iena[16]
port 107 nsew signal output
rlabel metal2 s 59910 163200 59966 164000 6 la_iena[17]
port 108 nsew signal output
rlabel metal2 s 63222 163200 63278 164000 6 la_iena[18]
port 109 nsew signal output
rlabel metal2 s 66534 163200 66590 164000 6 la_iena[19]
port 110 nsew signal output
rlabel metal2 s 6918 163200 6974 164000 6 la_iena[1]
port 111 nsew signal output
rlabel metal2 s 69846 163200 69902 164000 6 la_iena[20]
port 112 nsew signal output
rlabel metal2 s 73158 163200 73214 164000 6 la_iena[21]
port 113 nsew signal output
rlabel metal2 s 76470 163200 76526 164000 6 la_iena[22]
port 114 nsew signal output
rlabel metal2 s 79782 163200 79838 164000 6 la_iena[23]
port 115 nsew signal output
rlabel metal2 s 83094 163200 83150 164000 6 la_iena[24]
port 116 nsew signal output
rlabel metal2 s 86406 163200 86462 164000 6 la_iena[25]
port 117 nsew signal output
rlabel metal2 s 89718 163200 89774 164000 6 la_iena[26]
port 118 nsew signal output
rlabel metal2 s 93030 163200 93086 164000 6 la_iena[27]
port 119 nsew signal output
rlabel metal2 s 96342 163200 96398 164000 6 la_iena[28]
port 120 nsew signal output
rlabel metal2 s 99654 163200 99710 164000 6 la_iena[29]
port 121 nsew signal output
rlabel metal2 s 10230 163200 10286 164000 6 la_iena[2]
port 122 nsew signal output
rlabel metal2 s 102966 163200 103022 164000 6 la_iena[30]
port 123 nsew signal output
rlabel metal2 s 106278 163200 106334 164000 6 la_iena[31]
port 124 nsew signal output
rlabel metal2 s 109590 163200 109646 164000 6 la_iena[32]
port 125 nsew signal output
rlabel metal2 s 112902 163200 112958 164000 6 la_iena[33]
port 126 nsew signal output
rlabel metal2 s 116214 163200 116270 164000 6 la_iena[34]
port 127 nsew signal output
rlabel metal2 s 119526 163200 119582 164000 6 la_iena[35]
port 128 nsew signal output
rlabel metal2 s 122838 163200 122894 164000 6 la_iena[36]
port 129 nsew signal output
rlabel metal2 s 126150 163200 126206 164000 6 la_iena[37]
port 130 nsew signal output
rlabel metal2 s 129462 163200 129518 164000 6 la_iena[38]
port 131 nsew signal output
rlabel metal2 s 132774 163200 132830 164000 6 la_iena[39]
port 132 nsew signal output
rlabel metal2 s 13542 163200 13598 164000 6 la_iena[3]
port 133 nsew signal output
rlabel metal2 s 136086 163200 136142 164000 6 la_iena[40]
port 134 nsew signal output
rlabel metal2 s 139398 163200 139454 164000 6 la_iena[41]
port 135 nsew signal output
rlabel metal2 s 142710 163200 142766 164000 6 la_iena[42]
port 136 nsew signal output
rlabel metal2 s 146022 163200 146078 164000 6 la_iena[43]
port 137 nsew signal output
rlabel metal2 s 149334 163200 149390 164000 6 la_iena[44]
port 138 nsew signal output
rlabel metal2 s 152646 163200 152702 164000 6 la_iena[45]
port 139 nsew signal output
rlabel metal2 s 155958 163200 156014 164000 6 la_iena[46]
port 140 nsew signal output
rlabel metal2 s 159270 163200 159326 164000 6 la_iena[47]
port 141 nsew signal output
rlabel metal2 s 162582 163200 162638 164000 6 la_iena[48]
port 142 nsew signal output
rlabel metal2 s 165894 163200 165950 164000 6 la_iena[49]
port 143 nsew signal output
rlabel metal2 s 16854 163200 16910 164000 6 la_iena[4]
port 144 nsew signal output
rlabel metal2 s 169206 163200 169262 164000 6 la_iena[50]
port 145 nsew signal output
rlabel metal2 s 172518 163200 172574 164000 6 la_iena[51]
port 146 nsew signal output
rlabel metal2 s 175830 163200 175886 164000 6 la_iena[52]
port 147 nsew signal output
rlabel metal2 s 179142 163200 179198 164000 6 la_iena[53]
port 148 nsew signal output
rlabel metal2 s 182454 163200 182510 164000 6 la_iena[54]
port 149 nsew signal output
rlabel metal2 s 185766 163200 185822 164000 6 la_iena[55]
port 150 nsew signal output
rlabel metal2 s 189078 163200 189134 164000 6 la_iena[56]
port 151 nsew signal output
rlabel metal2 s 192390 163200 192446 164000 6 la_iena[57]
port 152 nsew signal output
rlabel metal2 s 195702 163200 195758 164000 6 la_iena[58]
port 153 nsew signal output
rlabel metal2 s 199014 163200 199070 164000 6 la_iena[59]
port 154 nsew signal output
rlabel metal2 s 20166 163200 20222 164000 6 la_iena[5]
port 155 nsew signal output
rlabel metal2 s 202326 163200 202382 164000 6 la_iena[60]
port 156 nsew signal output
rlabel metal2 s 205638 163200 205694 164000 6 la_iena[61]
port 157 nsew signal output
rlabel metal2 s 208950 163200 209006 164000 6 la_iena[62]
port 158 nsew signal output
rlabel metal2 s 212262 163200 212318 164000 6 la_iena[63]
port 159 nsew signal output
rlabel metal2 s 215574 163200 215630 164000 6 la_iena[64]
port 160 nsew signal output
rlabel metal2 s 218886 163200 218942 164000 6 la_iena[65]
port 161 nsew signal output
rlabel metal2 s 222198 163200 222254 164000 6 la_iena[66]
port 162 nsew signal output
rlabel metal2 s 225510 163200 225566 164000 6 la_iena[67]
port 163 nsew signal output
rlabel metal2 s 228822 163200 228878 164000 6 la_iena[68]
port 164 nsew signal output
rlabel metal2 s 232134 163200 232190 164000 6 la_iena[69]
port 165 nsew signal output
rlabel metal2 s 23478 163200 23534 164000 6 la_iena[6]
port 166 nsew signal output
rlabel metal2 s 235446 163200 235502 164000 6 la_iena[70]
port 167 nsew signal output
rlabel metal2 s 240414 163200 240470 164000 6 la_iena[71]
port 168 nsew signal output
rlabel metal2 s 243726 163200 243782 164000 6 la_iena[72]
port 169 nsew signal output
rlabel metal2 s 247038 163200 247094 164000 6 la_iena[73]
port 170 nsew signal output
rlabel metal2 s 250350 163200 250406 164000 6 la_iena[74]
port 171 nsew signal output
rlabel metal2 s 253662 163200 253718 164000 6 la_iena[75]
port 172 nsew signal output
rlabel metal2 s 256974 163200 257030 164000 6 la_iena[76]
port 173 nsew signal output
rlabel metal2 s 260286 163200 260342 164000 6 la_iena[77]
port 174 nsew signal output
rlabel metal2 s 263598 163200 263654 164000 6 la_iena[78]
port 175 nsew signal output
rlabel metal2 s 266910 163200 266966 164000 6 la_iena[79]
port 176 nsew signal output
rlabel metal2 s 26790 163200 26846 164000 6 la_iena[7]
port 177 nsew signal output
rlabel metal2 s 270222 163200 270278 164000 6 la_iena[80]
port 178 nsew signal output
rlabel metal2 s 273534 163200 273590 164000 6 la_iena[81]
port 179 nsew signal output
rlabel metal2 s 276846 163200 276902 164000 6 la_iena[82]
port 180 nsew signal output
rlabel metal2 s 280158 163200 280214 164000 6 la_iena[83]
port 181 nsew signal output
rlabel metal2 s 283470 163200 283526 164000 6 la_iena[84]
port 182 nsew signal output
rlabel metal2 s 286782 163200 286838 164000 6 la_iena[85]
port 183 nsew signal output
rlabel metal2 s 290094 163200 290150 164000 6 la_iena[86]
port 184 nsew signal output
rlabel metal2 s 293406 163200 293462 164000 6 la_iena[87]
port 185 nsew signal output
rlabel metal2 s 296718 163200 296774 164000 6 la_iena[88]
port 186 nsew signal output
rlabel metal2 s 300030 163200 300086 164000 6 la_iena[89]
port 187 nsew signal output
rlabel metal2 s 30102 163200 30158 164000 6 la_iena[8]
port 188 nsew signal output
rlabel metal2 s 303342 163200 303398 164000 6 la_iena[90]
port 189 nsew signal output
rlabel metal2 s 306654 163200 306710 164000 6 la_iena[91]
port 190 nsew signal output
rlabel metal2 s 309966 163200 310022 164000 6 la_iena[92]
port 191 nsew signal output
rlabel metal2 s 313278 163200 313334 164000 6 la_iena[93]
port 192 nsew signal output
rlabel metal2 s 316590 163200 316646 164000 6 la_iena[94]
port 193 nsew signal output
rlabel metal2 s 319902 163200 319958 164000 6 la_iena[95]
port 194 nsew signal output
rlabel metal2 s 323214 163200 323270 164000 6 la_iena[96]
port 195 nsew signal output
rlabel metal2 s 326526 163200 326582 164000 6 la_iena[97]
port 196 nsew signal output
rlabel metal2 s 329838 163200 329894 164000 6 la_iena[98]
port 197 nsew signal output
rlabel metal2 s 333150 163200 333206 164000 6 la_iena[99]
port 198 nsew signal output
rlabel metal2 s 33414 163200 33470 164000 6 la_iena[9]
port 199 nsew signal output
rlabel metal2 s 4434 163200 4490 164000 6 la_input[0]
port 200 nsew signal input
rlabel metal2 s 337290 163200 337346 164000 6 la_input[100]
port 201 nsew signal input
rlabel metal2 s 340602 163200 340658 164000 6 la_input[101]
port 202 nsew signal input
rlabel metal2 s 343914 163200 343970 164000 6 la_input[102]
port 203 nsew signal input
rlabel metal2 s 347226 163200 347282 164000 6 la_input[103]
port 204 nsew signal input
rlabel metal2 s 350538 163200 350594 164000 6 la_input[104]
port 205 nsew signal input
rlabel metal2 s 353850 163200 353906 164000 6 la_input[105]
port 206 nsew signal input
rlabel metal2 s 357162 163200 357218 164000 6 la_input[106]
port 207 nsew signal input
rlabel metal2 s 360474 163200 360530 164000 6 la_input[107]
port 208 nsew signal input
rlabel metal2 s 363786 163200 363842 164000 6 la_input[108]
port 209 nsew signal input
rlabel metal2 s 367098 163200 367154 164000 6 la_input[109]
port 210 nsew signal input
rlabel metal2 s 37554 163200 37610 164000 6 la_input[10]
port 211 nsew signal input
rlabel metal2 s 370410 163200 370466 164000 6 la_input[110]
port 212 nsew signal input
rlabel metal2 s 373722 163200 373778 164000 6 la_input[111]
port 213 nsew signal input
rlabel metal2 s 377034 163200 377090 164000 6 la_input[112]
port 214 nsew signal input
rlabel metal2 s 380346 163200 380402 164000 6 la_input[113]
port 215 nsew signal input
rlabel metal2 s 383658 163200 383714 164000 6 la_input[114]
port 216 nsew signal input
rlabel metal2 s 386970 163200 387026 164000 6 la_input[115]
port 217 nsew signal input
rlabel metal2 s 390282 163200 390338 164000 6 la_input[116]
port 218 nsew signal input
rlabel metal2 s 393594 163200 393650 164000 6 la_input[117]
port 219 nsew signal input
rlabel metal2 s 396906 163200 396962 164000 6 la_input[118]
port 220 nsew signal input
rlabel metal2 s 400218 163200 400274 164000 6 la_input[119]
port 221 nsew signal input
rlabel metal2 s 40866 163200 40922 164000 6 la_input[11]
port 222 nsew signal input
rlabel metal2 s 403530 163200 403586 164000 6 la_input[120]
port 223 nsew signal input
rlabel metal2 s 406842 163200 406898 164000 6 la_input[121]
port 224 nsew signal input
rlabel metal2 s 410154 163200 410210 164000 6 la_input[122]
port 225 nsew signal input
rlabel metal2 s 413466 163200 413522 164000 6 la_input[123]
port 226 nsew signal input
rlabel metal2 s 416778 163200 416834 164000 6 la_input[124]
port 227 nsew signal input
rlabel metal2 s 420090 163200 420146 164000 6 la_input[125]
port 228 nsew signal input
rlabel metal2 s 423402 163200 423458 164000 6 la_input[126]
port 229 nsew signal input
rlabel metal2 s 426714 163200 426770 164000 6 la_input[127]
port 230 nsew signal input
rlabel metal2 s 44178 163200 44234 164000 6 la_input[12]
port 231 nsew signal input
rlabel metal2 s 47490 163200 47546 164000 6 la_input[13]
port 232 nsew signal input
rlabel metal2 s 50802 163200 50858 164000 6 la_input[14]
port 233 nsew signal input
rlabel metal2 s 54114 163200 54170 164000 6 la_input[15]
port 234 nsew signal input
rlabel metal2 s 57426 163200 57482 164000 6 la_input[16]
port 235 nsew signal input
rlabel metal2 s 60738 163200 60794 164000 6 la_input[17]
port 236 nsew signal input
rlabel metal2 s 64050 163200 64106 164000 6 la_input[18]
port 237 nsew signal input
rlabel metal2 s 67362 163200 67418 164000 6 la_input[19]
port 238 nsew signal input
rlabel metal2 s 7746 163200 7802 164000 6 la_input[1]
port 239 nsew signal input
rlabel metal2 s 70674 163200 70730 164000 6 la_input[20]
port 240 nsew signal input
rlabel metal2 s 73986 163200 74042 164000 6 la_input[21]
port 241 nsew signal input
rlabel metal2 s 77298 163200 77354 164000 6 la_input[22]
port 242 nsew signal input
rlabel metal2 s 80610 163200 80666 164000 6 la_input[23]
port 243 nsew signal input
rlabel metal2 s 83922 163200 83978 164000 6 la_input[24]
port 244 nsew signal input
rlabel metal2 s 87234 163200 87290 164000 6 la_input[25]
port 245 nsew signal input
rlabel metal2 s 90546 163200 90602 164000 6 la_input[26]
port 246 nsew signal input
rlabel metal2 s 93858 163200 93914 164000 6 la_input[27]
port 247 nsew signal input
rlabel metal2 s 97170 163200 97226 164000 6 la_input[28]
port 248 nsew signal input
rlabel metal2 s 100482 163200 100538 164000 6 la_input[29]
port 249 nsew signal input
rlabel metal2 s 11058 163200 11114 164000 6 la_input[2]
port 250 nsew signal input
rlabel metal2 s 103794 163200 103850 164000 6 la_input[30]
port 251 nsew signal input
rlabel metal2 s 107106 163200 107162 164000 6 la_input[31]
port 252 nsew signal input
rlabel metal2 s 110418 163200 110474 164000 6 la_input[32]
port 253 nsew signal input
rlabel metal2 s 113730 163200 113786 164000 6 la_input[33]
port 254 nsew signal input
rlabel metal2 s 117042 163200 117098 164000 6 la_input[34]
port 255 nsew signal input
rlabel metal2 s 120354 163200 120410 164000 6 la_input[35]
port 256 nsew signal input
rlabel metal2 s 123666 163200 123722 164000 6 la_input[36]
port 257 nsew signal input
rlabel metal2 s 126978 163200 127034 164000 6 la_input[37]
port 258 nsew signal input
rlabel metal2 s 130290 163200 130346 164000 6 la_input[38]
port 259 nsew signal input
rlabel metal2 s 133602 163200 133658 164000 6 la_input[39]
port 260 nsew signal input
rlabel metal2 s 14370 163200 14426 164000 6 la_input[3]
port 261 nsew signal input
rlabel metal2 s 136914 163200 136970 164000 6 la_input[40]
port 262 nsew signal input
rlabel metal2 s 140226 163200 140282 164000 6 la_input[41]
port 263 nsew signal input
rlabel metal2 s 143538 163200 143594 164000 6 la_input[42]
port 264 nsew signal input
rlabel metal2 s 146850 163200 146906 164000 6 la_input[43]
port 265 nsew signal input
rlabel metal2 s 150162 163200 150218 164000 6 la_input[44]
port 266 nsew signal input
rlabel metal2 s 153474 163200 153530 164000 6 la_input[45]
port 267 nsew signal input
rlabel metal2 s 156786 163200 156842 164000 6 la_input[46]
port 268 nsew signal input
rlabel metal2 s 160098 163200 160154 164000 6 la_input[47]
port 269 nsew signal input
rlabel metal2 s 163410 163200 163466 164000 6 la_input[48]
port 270 nsew signal input
rlabel metal2 s 166722 163200 166778 164000 6 la_input[49]
port 271 nsew signal input
rlabel metal2 s 17682 163200 17738 164000 6 la_input[4]
port 272 nsew signal input
rlabel metal2 s 170034 163200 170090 164000 6 la_input[50]
port 273 nsew signal input
rlabel metal2 s 173346 163200 173402 164000 6 la_input[51]
port 274 nsew signal input
rlabel metal2 s 176658 163200 176714 164000 6 la_input[52]
port 275 nsew signal input
rlabel metal2 s 179970 163200 180026 164000 6 la_input[53]
port 276 nsew signal input
rlabel metal2 s 183282 163200 183338 164000 6 la_input[54]
port 277 nsew signal input
rlabel metal2 s 186594 163200 186650 164000 6 la_input[55]
port 278 nsew signal input
rlabel metal2 s 189906 163200 189962 164000 6 la_input[56]
port 279 nsew signal input
rlabel metal2 s 193218 163200 193274 164000 6 la_input[57]
port 280 nsew signal input
rlabel metal2 s 196530 163200 196586 164000 6 la_input[58]
port 281 nsew signal input
rlabel metal2 s 199842 163200 199898 164000 6 la_input[59]
port 282 nsew signal input
rlabel metal2 s 20994 163200 21050 164000 6 la_input[5]
port 283 nsew signal input
rlabel metal2 s 203154 163200 203210 164000 6 la_input[60]
port 284 nsew signal input
rlabel metal2 s 206466 163200 206522 164000 6 la_input[61]
port 285 nsew signal input
rlabel metal2 s 209778 163200 209834 164000 6 la_input[62]
port 286 nsew signal input
rlabel metal2 s 213090 163200 213146 164000 6 la_input[63]
port 287 nsew signal input
rlabel metal2 s 216402 163200 216458 164000 6 la_input[64]
port 288 nsew signal input
rlabel metal2 s 219714 163200 219770 164000 6 la_input[65]
port 289 nsew signal input
rlabel metal2 s 223026 163200 223082 164000 6 la_input[66]
port 290 nsew signal input
rlabel metal2 s 226338 163200 226394 164000 6 la_input[67]
port 291 nsew signal input
rlabel metal2 s 229650 163200 229706 164000 6 la_input[68]
port 292 nsew signal input
rlabel metal2 s 232962 163200 233018 164000 6 la_input[69]
port 293 nsew signal input
rlabel metal2 s 24306 163200 24362 164000 6 la_input[6]
port 294 nsew signal input
rlabel metal2 s 236274 163200 236330 164000 6 la_input[70]
port 295 nsew signal input
rlabel metal2 s 241242 163200 241298 164000 6 la_input[71]
port 296 nsew signal input
rlabel metal2 s 244554 163200 244610 164000 6 la_input[72]
port 297 nsew signal input
rlabel metal2 s 247866 163200 247922 164000 6 la_input[73]
port 298 nsew signal input
rlabel metal2 s 251178 163200 251234 164000 6 la_input[74]
port 299 nsew signal input
rlabel metal2 s 254490 163200 254546 164000 6 la_input[75]
port 300 nsew signal input
rlabel metal2 s 257802 163200 257858 164000 6 la_input[76]
port 301 nsew signal input
rlabel metal2 s 261114 163200 261170 164000 6 la_input[77]
port 302 nsew signal input
rlabel metal2 s 264426 163200 264482 164000 6 la_input[78]
port 303 nsew signal input
rlabel metal2 s 267738 163200 267794 164000 6 la_input[79]
port 304 nsew signal input
rlabel metal2 s 27618 163200 27674 164000 6 la_input[7]
port 305 nsew signal input
rlabel metal2 s 271050 163200 271106 164000 6 la_input[80]
port 306 nsew signal input
rlabel metal2 s 274362 163200 274418 164000 6 la_input[81]
port 307 nsew signal input
rlabel metal2 s 277674 163200 277730 164000 6 la_input[82]
port 308 nsew signal input
rlabel metal2 s 280986 163200 281042 164000 6 la_input[83]
port 309 nsew signal input
rlabel metal2 s 284298 163200 284354 164000 6 la_input[84]
port 310 nsew signal input
rlabel metal2 s 287610 163200 287666 164000 6 la_input[85]
port 311 nsew signal input
rlabel metal2 s 290922 163200 290978 164000 6 la_input[86]
port 312 nsew signal input
rlabel metal2 s 294234 163200 294290 164000 6 la_input[87]
port 313 nsew signal input
rlabel metal2 s 297546 163200 297602 164000 6 la_input[88]
port 314 nsew signal input
rlabel metal2 s 300858 163200 300914 164000 6 la_input[89]
port 315 nsew signal input
rlabel metal2 s 30930 163200 30986 164000 6 la_input[8]
port 316 nsew signal input
rlabel metal2 s 304170 163200 304226 164000 6 la_input[90]
port 317 nsew signal input
rlabel metal2 s 307482 163200 307538 164000 6 la_input[91]
port 318 nsew signal input
rlabel metal2 s 310794 163200 310850 164000 6 la_input[92]
port 319 nsew signal input
rlabel metal2 s 314106 163200 314162 164000 6 la_input[93]
port 320 nsew signal input
rlabel metal2 s 317418 163200 317474 164000 6 la_input[94]
port 321 nsew signal input
rlabel metal2 s 320730 163200 320786 164000 6 la_input[95]
port 322 nsew signal input
rlabel metal2 s 324042 163200 324098 164000 6 la_input[96]
port 323 nsew signal input
rlabel metal2 s 327354 163200 327410 164000 6 la_input[97]
port 324 nsew signal input
rlabel metal2 s 330666 163200 330722 164000 6 la_input[98]
port 325 nsew signal input
rlabel metal2 s 333978 163200 334034 164000 6 la_input[99]
port 326 nsew signal input
rlabel metal2 s 34242 163200 34298 164000 6 la_input[9]
port 327 nsew signal input
rlabel metal2 s 5262 163200 5318 164000 6 la_oenb[0]
port 328 nsew signal output
rlabel metal2 s 338118 163200 338174 164000 6 la_oenb[100]
port 329 nsew signal output
rlabel metal2 s 341430 163200 341486 164000 6 la_oenb[101]
port 330 nsew signal output
rlabel metal2 s 344742 163200 344798 164000 6 la_oenb[102]
port 331 nsew signal output
rlabel metal2 s 348054 163200 348110 164000 6 la_oenb[103]
port 332 nsew signal output
rlabel metal2 s 351366 163200 351422 164000 6 la_oenb[104]
port 333 nsew signal output
rlabel metal2 s 354678 163200 354734 164000 6 la_oenb[105]
port 334 nsew signal output
rlabel metal2 s 357990 163200 358046 164000 6 la_oenb[106]
port 335 nsew signal output
rlabel metal2 s 361302 163200 361358 164000 6 la_oenb[107]
port 336 nsew signal output
rlabel metal2 s 364614 163200 364670 164000 6 la_oenb[108]
port 337 nsew signal output
rlabel metal2 s 367926 163200 367982 164000 6 la_oenb[109]
port 338 nsew signal output
rlabel metal2 s 38382 163200 38438 164000 6 la_oenb[10]
port 339 nsew signal output
rlabel metal2 s 371238 163200 371294 164000 6 la_oenb[110]
port 340 nsew signal output
rlabel metal2 s 374550 163200 374606 164000 6 la_oenb[111]
port 341 nsew signal output
rlabel metal2 s 377862 163200 377918 164000 6 la_oenb[112]
port 342 nsew signal output
rlabel metal2 s 381174 163200 381230 164000 6 la_oenb[113]
port 343 nsew signal output
rlabel metal2 s 384486 163200 384542 164000 6 la_oenb[114]
port 344 nsew signal output
rlabel metal2 s 387798 163200 387854 164000 6 la_oenb[115]
port 345 nsew signal output
rlabel metal2 s 391110 163200 391166 164000 6 la_oenb[116]
port 346 nsew signal output
rlabel metal2 s 394422 163200 394478 164000 6 la_oenb[117]
port 347 nsew signal output
rlabel metal2 s 397734 163200 397790 164000 6 la_oenb[118]
port 348 nsew signal output
rlabel metal2 s 401046 163200 401102 164000 6 la_oenb[119]
port 349 nsew signal output
rlabel metal2 s 41694 163200 41750 164000 6 la_oenb[11]
port 350 nsew signal output
rlabel metal2 s 404358 163200 404414 164000 6 la_oenb[120]
port 351 nsew signal output
rlabel metal2 s 407670 163200 407726 164000 6 la_oenb[121]
port 352 nsew signal output
rlabel metal2 s 410982 163200 411038 164000 6 la_oenb[122]
port 353 nsew signal output
rlabel metal2 s 414294 163200 414350 164000 6 la_oenb[123]
port 354 nsew signal output
rlabel metal2 s 417606 163200 417662 164000 6 la_oenb[124]
port 355 nsew signal output
rlabel metal2 s 420918 163200 420974 164000 6 la_oenb[125]
port 356 nsew signal output
rlabel metal2 s 424230 163200 424286 164000 6 la_oenb[126]
port 357 nsew signal output
rlabel metal2 s 427542 163200 427598 164000 6 la_oenb[127]
port 358 nsew signal output
rlabel metal2 s 45006 163200 45062 164000 6 la_oenb[12]
port 359 nsew signal output
rlabel metal2 s 48318 163200 48374 164000 6 la_oenb[13]
port 360 nsew signal output
rlabel metal2 s 51630 163200 51686 164000 6 la_oenb[14]
port 361 nsew signal output
rlabel metal2 s 54942 163200 54998 164000 6 la_oenb[15]
port 362 nsew signal output
rlabel metal2 s 58254 163200 58310 164000 6 la_oenb[16]
port 363 nsew signal output
rlabel metal2 s 61566 163200 61622 164000 6 la_oenb[17]
port 364 nsew signal output
rlabel metal2 s 64878 163200 64934 164000 6 la_oenb[18]
port 365 nsew signal output
rlabel metal2 s 68190 163200 68246 164000 6 la_oenb[19]
port 366 nsew signal output
rlabel metal2 s 8574 163200 8630 164000 6 la_oenb[1]
port 367 nsew signal output
rlabel metal2 s 71502 163200 71558 164000 6 la_oenb[20]
port 368 nsew signal output
rlabel metal2 s 74814 163200 74870 164000 6 la_oenb[21]
port 369 nsew signal output
rlabel metal2 s 78126 163200 78182 164000 6 la_oenb[22]
port 370 nsew signal output
rlabel metal2 s 81438 163200 81494 164000 6 la_oenb[23]
port 371 nsew signal output
rlabel metal2 s 84750 163200 84806 164000 6 la_oenb[24]
port 372 nsew signal output
rlabel metal2 s 88062 163200 88118 164000 6 la_oenb[25]
port 373 nsew signal output
rlabel metal2 s 91374 163200 91430 164000 6 la_oenb[26]
port 374 nsew signal output
rlabel metal2 s 94686 163200 94742 164000 6 la_oenb[27]
port 375 nsew signal output
rlabel metal2 s 97998 163200 98054 164000 6 la_oenb[28]
port 376 nsew signal output
rlabel metal2 s 101310 163200 101366 164000 6 la_oenb[29]
port 377 nsew signal output
rlabel metal2 s 11886 163200 11942 164000 6 la_oenb[2]
port 378 nsew signal output
rlabel metal2 s 104622 163200 104678 164000 6 la_oenb[30]
port 379 nsew signal output
rlabel metal2 s 107934 163200 107990 164000 6 la_oenb[31]
port 380 nsew signal output
rlabel metal2 s 111246 163200 111302 164000 6 la_oenb[32]
port 381 nsew signal output
rlabel metal2 s 114558 163200 114614 164000 6 la_oenb[33]
port 382 nsew signal output
rlabel metal2 s 117870 163200 117926 164000 6 la_oenb[34]
port 383 nsew signal output
rlabel metal2 s 121182 163200 121238 164000 6 la_oenb[35]
port 384 nsew signal output
rlabel metal2 s 124494 163200 124550 164000 6 la_oenb[36]
port 385 nsew signal output
rlabel metal2 s 127806 163200 127862 164000 6 la_oenb[37]
port 386 nsew signal output
rlabel metal2 s 131118 163200 131174 164000 6 la_oenb[38]
port 387 nsew signal output
rlabel metal2 s 134430 163200 134486 164000 6 la_oenb[39]
port 388 nsew signal output
rlabel metal2 s 15198 163200 15254 164000 6 la_oenb[3]
port 389 nsew signal output
rlabel metal2 s 137742 163200 137798 164000 6 la_oenb[40]
port 390 nsew signal output
rlabel metal2 s 141054 163200 141110 164000 6 la_oenb[41]
port 391 nsew signal output
rlabel metal2 s 144366 163200 144422 164000 6 la_oenb[42]
port 392 nsew signal output
rlabel metal2 s 147678 163200 147734 164000 6 la_oenb[43]
port 393 nsew signal output
rlabel metal2 s 150990 163200 151046 164000 6 la_oenb[44]
port 394 nsew signal output
rlabel metal2 s 154302 163200 154358 164000 6 la_oenb[45]
port 395 nsew signal output
rlabel metal2 s 157614 163200 157670 164000 6 la_oenb[46]
port 396 nsew signal output
rlabel metal2 s 160926 163200 160982 164000 6 la_oenb[47]
port 397 nsew signal output
rlabel metal2 s 164238 163200 164294 164000 6 la_oenb[48]
port 398 nsew signal output
rlabel metal2 s 167550 163200 167606 164000 6 la_oenb[49]
port 399 nsew signal output
rlabel metal2 s 18510 163200 18566 164000 6 la_oenb[4]
port 400 nsew signal output
rlabel metal2 s 170862 163200 170918 164000 6 la_oenb[50]
port 401 nsew signal output
rlabel metal2 s 174174 163200 174230 164000 6 la_oenb[51]
port 402 nsew signal output
rlabel metal2 s 177486 163200 177542 164000 6 la_oenb[52]
port 403 nsew signal output
rlabel metal2 s 180798 163200 180854 164000 6 la_oenb[53]
port 404 nsew signal output
rlabel metal2 s 184110 163200 184166 164000 6 la_oenb[54]
port 405 nsew signal output
rlabel metal2 s 187422 163200 187478 164000 6 la_oenb[55]
port 406 nsew signal output
rlabel metal2 s 190734 163200 190790 164000 6 la_oenb[56]
port 407 nsew signal output
rlabel metal2 s 194046 163200 194102 164000 6 la_oenb[57]
port 408 nsew signal output
rlabel metal2 s 197358 163200 197414 164000 6 la_oenb[58]
port 409 nsew signal output
rlabel metal2 s 200670 163200 200726 164000 6 la_oenb[59]
port 410 nsew signal output
rlabel metal2 s 21822 163200 21878 164000 6 la_oenb[5]
port 411 nsew signal output
rlabel metal2 s 203982 163200 204038 164000 6 la_oenb[60]
port 412 nsew signal output
rlabel metal2 s 207294 163200 207350 164000 6 la_oenb[61]
port 413 nsew signal output
rlabel metal2 s 210606 163200 210662 164000 6 la_oenb[62]
port 414 nsew signal output
rlabel metal2 s 213918 163200 213974 164000 6 la_oenb[63]
port 415 nsew signal output
rlabel metal2 s 217230 163200 217286 164000 6 la_oenb[64]
port 416 nsew signal output
rlabel metal2 s 220542 163200 220598 164000 6 la_oenb[65]
port 417 nsew signal output
rlabel metal2 s 223854 163200 223910 164000 6 la_oenb[66]
port 418 nsew signal output
rlabel metal2 s 227166 163200 227222 164000 6 la_oenb[67]
port 419 nsew signal output
rlabel metal2 s 230478 163200 230534 164000 6 la_oenb[68]
port 420 nsew signal output
rlabel metal2 s 233790 163200 233846 164000 6 la_oenb[69]
port 421 nsew signal output
rlabel metal2 s 25134 163200 25190 164000 6 la_oenb[6]
port 422 nsew signal output
rlabel metal2 s 237102 163200 237158 164000 6 la_oenb[70]
port 423 nsew signal output
rlabel metal2 s 242070 163200 242126 164000 6 la_oenb[71]
port 424 nsew signal output
rlabel metal2 s 245382 163200 245438 164000 6 la_oenb[72]
port 425 nsew signal output
rlabel metal2 s 248694 163200 248750 164000 6 la_oenb[73]
port 426 nsew signal output
rlabel metal2 s 252006 163200 252062 164000 6 la_oenb[74]
port 427 nsew signal output
rlabel metal2 s 255318 163200 255374 164000 6 la_oenb[75]
port 428 nsew signal output
rlabel metal2 s 258630 163200 258686 164000 6 la_oenb[76]
port 429 nsew signal output
rlabel metal2 s 261942 163200 261998 164000 6 la_oenb[77]
port 430 nsew signal output
rlabel metal2 s 265254 163200 265310 164000 6 la_oenb[78]
port 431 nsew signal output
rlabel metal2 s 268566 163200 268622 164000 6 la_oenb[79]
port 432 nsew signal output
rlabel metal2 s 28446 163200 28502 164000 6 la_oenb[7]
port 433 nsew signal output
rlabel metal2 s 271878 163200 271934 164000 6 la_oenb[80]
port 434 nsew signal output
rlabel metal2 s 275190 163200 275246 164000 6 la_oenb[81]
port 435 nsew signal output
rlabel metal2 s 278502 163200 278558 164000 6 la_oenb[82]
port 436 nsew signal output
rlabel metal2 s 281814 163200 281870 164000 6 la_oenb[83]
port 437 nsew signal output
rlabel metal2 s 285126 163200 285182 164000 6 la_oenb[84]
port 438 nsew signal output
rlabel metal2 s 288438 163200 288494 164000 6 la_oenb[85]
port 439 nsew signal output
rlabel metal2 s 291750 163200 291806 164000 6 la_oenb[86]
port 440 nsew signal output
rlabel metal2 s 295062 163200 295118 164000 6 la_oenb[87]
port 441 nsew signal output
rlabel metal2 s 298374 163200 298430 164000 6 la_oenb[88]
port 442 nsew signal output
rlabel metal2 s 301686 163200 301742 164000 6 la_oenb[89]
port 443 nsew signal output
rlabel metal2 s 31758 163200 31814 164000 6 la_oenb[8]
port 444 nsew signal output
rlabel metal2 s 304998 163200 305054 164000 6 la_oenb[90]
port 445 nsew signal output
rlabel metal2 s 308310 163200 308366 164000 6 la_oenb[91]
port 446 nsew signal output
rlabel metal2 s 311622 163200 311678 164000 6 la_oenb[92]
port 447 nsew signal output
rlabel metal2 s 314934 163200 314990 164000 6 la_oenb[93]
port 448 nsew signal output
rlabel metal2 s 318246 163200 318302 164000 6 la_oenb[94]
port 449 nsew signal output
rlabel metal2 s 321558 163200 321614 164000 6 la_oenb[95]
port 450 nsew signal output
rlabel metal2 s 324870 163200 324926 164000 6 la_oenb[96]
port 451 nsew signal output
rlabel metal2 s 328182 163200 328238 164000 6 la_oenb[97]
port 452 nsew signal output
rlabel metal2 s 331494 163200 331550 164000 6 la_oenb[98]
port 453 nsew signal output
rlabel metal2 s 334806 163200 334862 164000 6 la_oenb[99]
port 454 nsew signal output
rlabel metal2 s 35070 163200 35126 164000 6 la_oenb[9]
port 455 nsew signal output
rlabel metal2 s 6090 163200 6146 164000 6 la_output[0]
port 456 nsew signal output
rlabel metal2 s 338946 163200 339002 164000 6 la_output[100]
port 457 nsew signal output
rlabel metal2 s 342258 163200 342314 164000 6 la_output[101]
port 458 nsew signal output
rlabel metal2 s 345570 163200 345626 164000 6 la_output[102]
port 459 nsew signal output
rlabel metal2 s 348882 163200 348938 164000 6 la_output[103]
port 460 nsew signal output
rlabel metal2 s 352194 163200 352250 164000 6 la_output[104]
port 461 nsew signal output
rlabel metal2 s 355506 163200 355562 164000 6 la_output[105]
port 462 nsew signal output
rlabel metal2 s 358818 163200 358874 164000 6 la_output[106]
port 463 nsew signal output
rlabel metal2 s 362130 163200 362186 164000 6 la_output[107]
port 464 nsew signal output
rlabel metal2 s 365442 163200 365498 164000 6 la_output[108]
port 465 nsew signal output
rlabel metal2 s 368754 163200 368810 164000 6 la_output[109]
port 466 nsew signal output
rlabel metal2 s 39210 163200 39266 164000 6 la_output[10]
port 467 nsew signal output
rlabel metal2 s 372066 163200 372122 164000 6 la_output[110]
port 468 nsew signal output
rlabel metal2 s 375378 163200 375434 164000 6 la_output[111]
port 469 nsew signal output
rlabel metal2 s 378690 163200 378746 164000 6 la_output[112]
port 470 nsew signal output
rlabel metal2 s 382002 163200 382058 164000 6 la_output[113]
port 471 nsew signal output
rlabel metal2 s 385314 163200 385370 164000 6 la_output[114]
port 472 nsew signal output
rlabel metal2 s 388626 163200 388682 164000 6 la_output[115]
port 473 nsew signal output
rlabel metal2 s 391938 163200 391994 164000 6 la_output[116]
port 474 nsew signal output
rlabel metal2 s 395250 163200 395306 164000 6 la_output[117]
port 475 nsew signal output
rlabel metal2 s 398562 163200 398618 164000 6 la_output[118]
port 476 nsew signal output
rlabel metal2 s 401874 163200 401930 164000 6 la_output[119]
port 477 nsew signal output
rlabel metal2 s 42522 163200 42578 164000 6 la_output[11]
port 478 nsew signal output
rlabel metal2 s 405186 163200 405242 164000 6 la_output[120]
port 479 nsew signal output
rlabel metal2 s 408498 163200 408554 164000 6 la_output[121]
port 480 nsew signal output
rlabel metal2 s 411810 163200 411866 164000 6 la_output[122]
port 481 nsew signal output
rlabel metal2 s 415122 163200 415178 164000 6 la_output[123]
port 482 nsew signal output
rlabel metal2 s 418434 163200 418490 164000 6 la_output[124]
port 483 nsew signal output
rlabel metal2 s 421746 163200 421802 164000 6 la_output[125]
port 484 nsew signal output
rlabel metal2 s 425058 163200 425114 164000 6 la_output[126]
port 485 nsew signal output
rlabel metal2 s 428370 163200 428426 164000 6 la_output[127]
port 486 nsew signal output
rlabel metal2 s 45834 163200 45890 164000 6 la_output[12]
port 487 nsew signal output
rlabel metal2 s 49146 163200 49202 164000 6 la_output[13]
port 488 nsew signal output
rlabel metal2 s 52458 163200 52514 164000 6 la_output[14]
port 489 nsew signal output
rlabel metal2 s 55770 163200 55826 164000 6 la_output[15]
port 490 nsew signal output
rlabel metal2 s 59082 163200 59138 164000 6 la_output[16]
port 491 nsew signal output
rlabel metal2 s 62394 163200 62450 164000 6 la_output[17]
port 492 nsew signal output
rlabel metal2 s 65706 163200 65762 164000 6 la_output[18]
port 493 nsew signal output
rlabel metal2 s 69018 163200 69074 164000 6 la_output[19]
port 494 nsew signal output
rlabel metal2 s 9402 163200 9458 164000 6 la_output[1]
port 495 nsew signal output
rlabel metal2 s 72330 163200 72386 164000 6 la_output[20]
port 496 nsew signal output
rlabel metal2 s 75642 163200 75698 164000 6 la_output[21]
port 497 nsew signal output
rlabel metal2 s 78954 163200 79010 164000 6 la_output[22]
port 498 nsew signal output
rlabel metal2 s 82266 163200 82322 164000 6 la_output[23]
port 499 nsew signal output
rlabel metal2 s 85578 163200 85634 164000 6 la_output[24]
port 500 nsew signal output
rlabel metal2 s 88890 163200 88946 164000 6 la_output[25]
port 501 nsew signal output
rlabel metal2 s 92202 163200 92258 164000 6 la_output[26]
port 502 nsew signal output
rlabel metal2 s 95514 163200 95570 164000 6 la_output[27]
port 503 nsew signal output
rlabel metal2 s 98826 163200 98882 164000 6 la_output[28]
port 504 nsew signal output
rlabel metal2 s 102138 163200 102194 164000 6 la_output[29]
port 505 nsew signal output
rlabel metal2 s 12714 163200 12770 164000 6 la_output[2]
port 506 nsew signal output
rlabel metal2 s 105450 163200 105506 164000 6 la_output[30]
port 507 nsew signal output
rlabel metal2 s 108762 163200 108818 164000 6 la_output[31]
port 508 nsew signal output
rlabel metal2 s 112074 163200 112130 164000 6 la_output[32]
port 509 nsew signal output
rlabel metal2 s 115386 163200 115442 164000 6 la_output[33]
port 510 nsew signal output
rlabel metal2 s 118698 163200 118754 164000 6 la_output[34]
port 511 nsew signal output
rlabel metal2 s 122010 163200 122066 164000 6 la_output[35]
port 512 nsew signal output
rlabel metal2 s 125322 163200 125378 164000 6 la_output[36]
port 513 nsew signal output
rlabel metal2 s 128634 163200 128690 164000 6 la_output[37]
port 514 nsew signal output
rlabel metal2 s 131946 163200 132002 164000 6 la_output[38]
port 515 nsew signal output
rlabel metal2 s 135258 163200 135314 164000 6 la_output[39]
port 516 nsew signal output
rlabel metal2 s 16026 163200 16082 164000 6 la_output[3]
port 517 nsew signal output
rlabel metal2 s 138570 163200 138626 164000 6 la_output[40]
port 518 nsew signal output
rlabel metal2 s 141882 163200 141938 164000 6 la_output[41]
port 519 nsew signal output
rlabel metal2 s 145194 163200 145250 164000 6 la_output[42]
port 520 nsew signal output
rlabel metal2 s 148506 163200 148562 164000 6 la_output[43]
port 521 nsew signal output
rlabel metal2 s 151818 163200 151874 164000 6 la_output[44]
port 522 nsew signal output
rlabel metal2 s 155130 163200 155186 164000 6 la_output[45]
port 523 nsew signal output
rlabel metal2 s 158442 163200 158498 164000 6 la_output[46]
port 524 nsew signal output
rlabel metal2 s 161754 163200 161810 164000 6 la_output[47]
port 525 nsew signal output
rlabel metal2 s 165066 163200 165122 164000 6 la_output[48]
port 526 nsew signal output
rlabel metal2 s 168378 163200 168434 164000 6 la_output[49]
port 527 nsew signal output
rlabel metal2 s 19338 163200 19394 164000 6 la_output[4]
port 528 nsew signal output
rlabel metal2 s 171690 163200 171746 164000 6 la_output[50]
port 529 nsew signal output
rlabel metal2 s 175002 163200 175058 164000 6 la_output[51]
port 530 nsew signal output
rlabel metal2 s 178314 163200 178370 164000 6 la_output[52]
port 531 nsew signal output
rlabel metal2 s 181626 163200 181682 164000 6 la_output[53]
port 532 nsew signal output
rlabel metal2 s 184938 163200 184994 164000 6 la_output[54]
port 533 nsew signal output
rlabel metal2 s 188250 163200 188306 164000 6 la_output[55]
port 534 nsew signal output
rlabel metal2 s 191562 163200 191618 164000 6 la_output[56]
port 535 nsew signal output
rlabel metal2 s 194874 163200 194930 164000 6 la_output[57]
port 536 nsew signal output
rlabel metal2 s 198186 163200 198242 164000 6 la_output[58]
port 537 nsew signal output
rlabel metal2 s 201498 163200 201554 164000 6 la_output[59]
port 538 nsew signal output
rlabel metal2 s 22650 163200 22706 164000 6 la_output[5]
port 539 nsew signal output
rlabel metal2 s 204810 163200 204866 164000 6 la_output[60]
port 540 nsew signal output
rlabel metal2 s 208122 163200 208178 164000 6 la_output[61]
port 541 nsew signal output
rlabel metal2 s 211434 163200 211490 164000 6 la_output[62]
port 542 nsew signal output
rlabel metal2 s 214746 163200 214802 164000 6 la_output[63]
port 543 nsew signal output
rlabel metal2 s 218058 163200 218114 164000 6 la_output[64]
port 544 nsew signal output
rlabel metal2 s 221370 163200 221426 164000 6 la_output[65]
port 545 nsew signal output
rlabel metal2 s 224682 163200 224738 164000 6 la_output[66]
port 546 nsew signal output
rlabel metal2 s 227994 163200 228050 164000 6 la_output[67]
port 547 nsew signal output
rlabel metal2 s 231306 163200 231362 164000 6 la_output[68]
port 548 nsew signal output
rlabel metal2 s 234618 163200 234674 164000 6 la_output[69]
port 549 nsew signal output
rlabel metal2 s 25962 163200 26018 164000 6 la_output[6]
port 550 nsew signal output
rlabel metal2 s 237930 163200 237986 164000 6 la_output[70]
port 551 nsew signal output
rlabel metal2 s 242898 163200 242954 164000 6 la_output[71]
port 552 nsew signal output
rlabel metal2 s 246210 163200 246266 164000 6 la_output[72]
port 553 nsew signal output
rlabel metal2 s 249522 163200 249578 164000 6 la_output[73]
port 554 nsew signal output
rlabel metal2 s 252834 163200 252890 164000 6 la_output[74]
port 555 nsew signal output
rlabel metal2 s 256146 163200 256202 164000 6 la_output[75]
port 556 nsew signal output
rlabel metal2 s 259458 163200 259514 164000 6 la_output[76]
port 557 nsew signal output
rlabel metal2 s 262770 163200 262826 164000 6 la_output[77]
port 558 nsew signal output
rlabel metal2 s 266082 163200 266138 164000 6 la_output[78]
port 559 nsew signal output
rlabel metal2 s 269394 163200 269450 164000 6 la_output[79]
port 560 nsew signal output
rlabel metal2 s 29274 163200 29330 164000 6 la_output[7]
port 561 nsew signal output
rlabel metal2 s 272706 163200 272762 164000 6 la_output[80]
port 562 nsew signal output
rlabel metal2 s 276018 163200 276074 164000 6 la_output[81]
port 563 nsew signal output
rlabel metal2 s 279330 163200 279386 164000 6 la_output[82]
port 564 nsew signal output
rlabel metal2 s 282642 163200 282698 164000 6 la_output[83]
port 565 nsew signal output
rlabel metal2 s 285954 163200 286010 164000 6 la_output[84]
port 566 nsew signal output
rlabel metal2 s 289266 163200 289322 164000 6 la_output[85]
port 567 nsew signal output
rlabel metal2 s 292578 163200 292634 164000 6 la_output[86]
port 568 nsew signal output
rlabel metal2 s 295890 163200 295946 164000 6 la_output[87]
port 569 nsew signal output
rlabel metal2 s 299202 163200 299258 164000 6 la_output[88]
port 570 nsew signal output
rlabel metal2 s 302514 163200 302570 164000 6 la_output[89]
port 571 nsew signal output
rlabel metal2 s 32586 163200 32642 164000 6 la_output[8]
port 572 nsew signal output
rlabel metal2 s 305826 163200 305882 164000 6 la_output[90]
port 573 nsew signal output
rlabel metal2 s 309138 163200 309194 164000 6 la_output[91]
port 574 nsew signal output
rlabel metal2 s 312450 163200 312506 164000 6 la_output[92]
port 575 nsew signal output
rlabel metal2 s 315762 163200 315818 164000 6 la_output[93]
port 576 nsew signal output
rlabel metal2 s 319074 163200 319130 164000 6 la_output[94]
port 577 nsew signal output
rlabel metal2 s 322386 163200 322442 164000 6 la_output[95]
port 578 nsew signal output
rlabel metal2 s 325698 163200 325754 164000 6 la_output[96]
port 579 nsew signal output
rlabel metal2 s 329010 163200 329066 164000 6 la_output[97]
port 580 nsew signal output
rlabel metal2 s 332322 163200 332378 164000 6 la_output[98]
port 581 nsew signal output
rlabel metal2 s 335634 163200 335690 164000 6 la_output[99]
port 582 nsew signal output
rlabel metal2 s 35898 163200 35954 164000 6 la_output[9]
port 583 nsew signal output
rlabel metal2 s 429198 163200 429254 164000 6 mprj_ack_i
port 584 nsew signal input
rlabel metal2 s 433338 163200 433394 164000 6 mprj_adr_o[0]
port 585 nsew signal output
rlabel metal2 s 461490 163200 461546 164000 6 mprj_adr_o[10]
port 586 nsew signal output
rlabel metal2 s 463974 163200 464030 164000 6 mprj_adr_o[11]
port 587 nsew signal output
rlabel metal2 s 466458 163200 466514 164000 6 mprj_adr_o[12]
port 588 nsew signal output
rlabel metal2 s 468942 163200 468998 164000 6 mprj_adr_o[13]
port 589 nsew signal output
rlabel metal2 s 471426 163200 471482 164000 6 mprj_adr_o[14]
port 590 nsew signal output
rlabel metal2 s 473910 163200 473966 164000 6 mprj_adr_o[15]
port 591 nsew signal output
rlabel metal2 s 476394 163200 476450 164000 6 mprj_adr_o[16]
port 592 nsew signal output
rlabel metal2 s 478878 163200 478934 164000 6 mprj_adr_o[17]
port 593 nsew signal output
rlabel metal2 s 481362 163200 481418 164000 6 mprj_adr_o[18]
port 594 nsew signal output
rlabel metal2 s 483846 163200 483902 164000 6 mprj_adr_o[19]
port 595 nsew signal output
rlabel metal2 s 436650 163200 436706 164000 6 mprj_adr_o[1]
port 596 nsew signal output
rlabel metal2 s 486330 163200 486386 164000 6 mprj_adr_o[20]
port 597 nsew signal output
rlabel metal2 s 488814 163200 488870 164000 6 mprj_adr_o[21]
port 598 nsew signal output
rlabel metal2 s 491298 163200 491354 164000 6 mprj_adr_o[22]
port 599 nsew signal output
rlabel metal2 s 493782 163200 493838 164000 6 mprj_adr_o[23]
port 600 nsew signal output
rlabel metal2 s 496266 163200 496322 164000 6 mprj_adr_o[24]
port 601 nsew signal output
rlabel metal2 s 498750 163200 498806 164000 6 mprj_adr_o[25]
port 602 nsew signal output
rlabel metal2 s 501234 163200 501290 164000 6 mprj_adr_o[26]
port 603 nsew signal output
rlabel metal2 s 503718 163200 503774 164000 6 mprj_adr_o[27]
port 604 nsew signal output
rlabel metal2 s 506202 163200 506258 164000 6 mprj_adr_o[28]
port 605 nsew signal output
rlabel metal2 s 508686 163200 508742 164000 6 mprj_adr_o[29]
port 606 nsew signal output
rlabel metal2 s 439962 163200 440018 164000 6 mprj_adr_o[2]
port 607 nsew signal output
rlabel metal2 s 511170 163200 511226 164000 6 mprj_adr_o[30]
port 608 nsew signal output
rlabel metal2 s 513654 163200 513710 164000 6 mprj_adr_o[31]
port 609 nsew signal output
rlabel metal2 s 443274 163200 443330 164000 6 mprj_adr_o[3]
port 610 nsew signal output
rlabel metal2 s 446586 163200 446642 164000 6 mprj_adr_o[4]
port 611 nsew signal output
rlabel metal2 s 449070 163200 449126 164000 6 mprj_adr_o[5]
port 612 nsew signal output
rlabel metal2 s 451554 163200 451610 164000 6 mprj_adr_o[6]
port 613 nsew signal output
rlabel metal2 s 454038 163200 454094 164000 6 mprj_adr_o[7]
port 614 nsew signal output
rlabel metal2 s 456522 163200 456578 164000 6 mprj_adr_o[8]
port 615 nsew signal output
rlabel metal2 s 459006 163200 459062 164000 6 mprj_adr_o[9]
port 616 nsew signal output
rlabel metal2 s 430026 163200 430082 164000 6 mprj_cyc_o
port 617 nsew signal output
rlabel metal2 s 434166 163200 434222 164000 6 mprj_dat_i[0]
port 618 nsew signal input
rlabel metal2 s 462318 163200 462374 164000 6 mprj_dat_i[10]
port 619 nsew signal input
rlabel metal2 s 464802 163200 464858 164000 6 mprj_dat_i[11]
port 620 nsew signal input
rlabel metal2 s 467286 163200 467342 164000 6 mprj_dat_i[12]
port 621 nsew signal input
rlabel metal2 s 469770 163200 469826 164000 6 mprj_dat_i[13]
port 622 nsew signal input
rlabel metal2 s 472254 163200 472310 164000 6 mprj_dat_i[14]
port 623 nsew signal input
rlabel metal2 s 474738 163200 474794 164000 6 mprj_dat_i[15]
port 624 nsew signal input
rlabel metal2 s 477222 163200 477278 164000 6 mprj_dat_i[16]
port 625 nsew signal input
rlabel metal2 s 479706 163200 479762 164000 6 mprj_dat_i[17]
port 626 nsew signal input
rlabel metal2 s 482190 163200 482246 164000 6 mprj_dat_i[18]
port 627 nsew signal input
rlabel metal2 s 484674 163200 484730 164000 6 mprj_dat_i[19]
port 628 nsew signal input
rlabel metal2 s 437478 163200 437534 164000 6 mprj_dat_i[1]
port 629 nsew signal input
rlabel metal2 s 487158 163200 487214 164000 6 mprj_dat_i[20]
port 630 nsew signal input
rlabel metal2 s 489642 163200 489698 164000 6 mprj_dat_i[21]
port 631 nsew signal input
rlabel metal2 s 492126 163200 492182 164000 6 mprj_dat_i[22]
port 632 nsew signal input
rlabel metal2 s 494610 163200 494666 164000 6 mprj_dat_i[23]
port 633 nsew signal input
rlabel metal2 s 497094 163200 497150 164000 6 mprj_dat_i[24]
port 634 nsew signal input
rlabel metal2 s 499578 163200 499634 164000 6 mprj_dat_i[25]
port 635 nsew signal input
rlabel metal2 s 502062 163200 502118 164000 6 mprj_dat_i[26]
port 636 nsew signal input
rlabel metal2 s 504546 163200 504602 164000 6 mprj_dat_i[27]
port 637 nsew signal input
rlabel metal2 s 507030 163200 507086 164000 6 mprj_dat_i[28]
port 638 nsew signal input
rlabel metal2 s 509514 163200 509570 164000 6 mprj_dat_i[29]
port 639 nsew signal input
rlabel metal2 s 440790 163200 440846 164000 6 mprj_dat_i[2]
port 640 nsew signal input
rlabel metal2 s 511998 163200 512054 164000 6 mprj_dat_i[30]
port 641 nsew signal input
rlabel metal2 s 514482 163200 514538 164000 6 mprj_dat_i[31]
port 642 nsew signal input
rlabel metal2 s 444102 163200 444158 164000 6 mprj_dat_i[3]
port 643 nsew signal input
rlabel metal2 s 447414 163200 447470 164000 6 mprj_dat_i[4]
port 644 nsew signal input
rlabel metal2 s 449898 163200 449954 164000 6 mprj_dat_i[5]
port 645 nsew signal input
rlabel metal2 s 452382 163200 452438 164000 6 mprj_dat_i[6]
port 646 nsew signal input
rlabel metal2 s 454866 163200 454922 164000 6 mprj_dat_i[7]
port 647 nsew signal input
rlabel metal2 s 457350 163200 457406 164000 6 mprj_dat_i[8]
port 648 nsew signal input
rlabel metal2 s 459834 163200 459890 164000 6 mprj_dat_i[9]
port 649 nsew signal input
rlabel metal2 s 434994 163200 435050 164000 6 mprj_dat_o[0]
port 650 nsew signal output
rlabel metal2 s 463146 163200 463202 164000 6 mprj_dat_o[10]
port 651 nsew signal output
rlabel metal2 s 465630 163200 465686 164000 6 mprj_dat_o[11]
port 652 nsew signal output
rlabel metal2 s 468114 163200 468170 164000 6 mprj_dat_o[12]
port 653 nsew signal output
rlabel metal2 s 470598 163200 470654 164000 6 mprj_dat_o[13]
port 654 nsew signal output
rlabel metal2 s 473082 163200 473138 164000 6 mprj_dat_o[14]
port 655 nsew signal output
rlabel metal2 s 475566 163200 475622 164000 6 mprj_dat_o[15]
port 656 nsew signal output
rlabel metal2 s 478050 163200 478106 164000 6 mprj_dat_o[16]
port 657 nsew signal output
rlabel metal2 s 480534 163200 480590 164000 6 mprj_dat_o[17]
port 658 nsew signal output
rlabel metal2 s 483018 163200 483074 164000 6 mprj_dat_o[18]
port 659 nsew signal output
rlabel metal2 s 485502 163200 485558 164000 6 mprj_dat_o[19]
port 660 nsew signal output
rlabel metal2 s 438306 163200 438362 164000 6 mprj_dat_o[1]
port 661 nsew signal output
rlabel metal2 s 487986 163200 488042 164000 6 mprj_dat_o[20]
port 662 nsew signal output
rlabel metal2 s 490470 163200 490526 164000 6 mprj_dat_o[21]
port 663 nsew signal output
rlabel metal2 s 492954 163200 493010 164000 6 mprj_dat_o[22]
port 664 nsew signal output
rlabel metal2 s 495438 163200 495494 164000 6 mprj_dat_o[23]
port 665 nsew signal output
rlabel metal2 s 497922 163200 497978 164000 6 mprj_dat_o[24]
port 666 nsew signal output
rlabel metal2 s 500406 163200 500462 164000 6 mprj_dat_o[25]
port 667 nsew signal output
rlabel metal2 s 502890 163200 502946 164000 6 mprj_dat_o[26]
port 668 nsew signal output
rlabel metal2 s 505374 163200 505430 164000 6 mprj_dat_o[27]
port 669 nsew signal output
rlabel metal2 s 507858 163200 507914 164000 6 mprj_dat_o[28]
port 670 nsew signal output
rlabel metal2 s 510342 163200 510398 164000 6 mprj_dat_o[29]
port 671 nsew signal output
rlabel metal2 s 441618 163200 441674 164000 6 mprj_dat_o[2]
port 672 nsew signal output
rlabel metal2 s 512826 163200 512882 164000 6 mprj_dat_o[30]
port 673 nsew signal output
rlabel metal2 s 515310 163200 515366 164000 6 mprj_dat_o[31]
port 674 nsew signal output
rlabel metal2 s 444930 163200 444986 164000 6 mprj_dat_o[3]
port 675 nsew signal output
rlabel metal2 s 448242 163200 448298 164000 6 mprj_dat_o[4]
port 676 nsew signal output
rlabel metal2 s 450726 163200 450782 164000 6 mprj_dat_o[5]
port 677 nsew signal output
rlabel metal2 s 453210 163200 453266 164000 6 mprj_dat_o[6]
port 678 nsew signal output
rlabel metal2 s 455694 163200 455750 164000 6 mprj_dat_o[7]
port 679 nsew signal output
rlabel metal2 s 458178 163200 458234 164000 6 mprj_dat_o[8]
port 680 nsew signal output
rlabel metal2 s 460662 163200 460718 164000 6 mprj_dat_o[9]
port 681 nsew signal output
rlabel metal2 s 435822 163200 435878 164000 6 mprj_sel_o[0]
port 682 nsew signal output
rlabel metal2 s 439134 163200 439190 164000 6 mprj_sel_o[1]
port 683 nsew signal output
rlabel metal2 s 442446 163200 442502 164000 6 mprj_sel_o[2]
port 684 nsew signal output
rlabel metal2 s 445758 163200 445814 164000 6 mprj_sel_o[3]
port 685 nsew signal output
rlabel metal2 s 430854 163200 430910 164000 6 mprj_stb_o
port 686 nsew signal output
rlabel metal2 s 431682 163200 431738 164000 6 mprj_wb_iena
port 687 nsew signal output
rlabel metal2 s 432510 163200 432566 164000 6 mprj_we_o
port 688 nsew signal output
rlabel metal3 s 523200 13336 524000 13456 6 por_l_in
port 689 nsew signal input
rlabel metal2 s 255972 0 256028 800 6 por_l_out
port 690 nsew signal output
rlabel metal3 s 523200 15512 524000 15632 6 porb_h_in
port 691 nsew signal input
rlabel metal2 s 257972 0 258028 800 6 porb_h_out
port 692 nsew signal output
rlabel metal3 s 523200 54680 524000 54800 6 qspi_enabled
port 693 nsew signal output
rlabel metal2 s 265972 0 266028 800 6 resetn_in
port 694 nsew signal input
rlabel metal2 s 239586 163200 239642 164000 6 resetn_out
port 695 nsew signal output
rlabel metal2 s 253972 0 254028 800 6 rstb_l_in
port 696 nsew signal input
rlabel metal3 s 523200 2456 524000 2576 6 rstb_l_out
port 697 nsew signal output
rlabel metal3 s 523200 45976 524000 46096 6 ser_rx
port 698 nsew signal input
rlabel metal3 s 523200 48152 524000 48272 6 ser_tx
port 699 nsew signal output
rlabel metal3 s 523200 11160 524000 11280 6 serial_clock_in
port 700 nsew signal input
rlabel metal3 s 0 143352 800 143472 6 serial_clock_out
port 701 nsew signal output
rlabel metal3 s 523200 6808 524000 6928 6 serial_data_2_in
port 702 nsew signal input
rlabel metal3 s 0 139352 800 139472 6 serial_data_2_out
port 703 nsew signal output
rlabel metal3 s 523200 4632 524000 4752 6 serial_load_in
port 704 nsew signal input
rlabel metal3 s 0 137352 800 137472 6 serial_load_out
port 705 nsew signal output
rlabel metal3 s 523200 8984 524000 9104 6 serial_resetn_in
port 706 nsew signal input
rlabel metal3 s 0 141352 800 141472 6 serial_resetn_out
port 707 nsew signal output
rlabel metal3 s 523200 41624 524000 41744 6 spi_csb
port 708 nsew signal output
rlabel metal3 s 523200 50328 524000 50448 6 spi_enabled
port 709 nsew signal output
rlabel metal3 s 523200 39448 524000 39568 6 spi_sck
port 710 nsew signal output
rlabel metal3 s 523200 43800 524000 43920 6 spi_sdi
port 711 nsew signal input
rlabel metal3 s 523200 37272 524000 37392 6 spi_sdo
port 712 nsew signal output
rlabel metal3 s 523200 35096 524000 35216 6 spi_sdoenb
port 713 nsew signal output
rlabel metal3 s 523200 26392 524000 26512 6 trap
port 714 nsew signal output
rlabel metal3 s 523200 52504 524000 52624 6 uart_enabled
port 715 nsew signal output
rlabel metal2 s 516138 163200 516194 164000 6 user_irq_ena[0]
port 716 nsew signal output
rlabel metal2 s 516966 163200 517022 164000 6 user_irq_ena[1]
port 717 nsew signal output
rlabel metal2 s 517794 163200 517850 164000 6 user_irq_ena[2]
port 718 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 524000 164000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 248498114
string GDS_FILE /home/hosni/mgmt_core_wrapper_hold_fix/caravel_mgmt_soc_litex/openlane/mgmt_core_wrapper/runs/RUN_2022.11.09_15.15.08/results/signoff/mgmt_core_wrapper.magic.gds
string GDS_START 93616930
<< end >>

