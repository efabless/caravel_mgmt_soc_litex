magic
tech sky130A
magscale 1 2
timestamp 1638138898
<< obsli1 >>
rect 5869 1785 578283 157335
<< obsm1 >>
rect 474 1096 578482 158976
<< metal2 >>
rect 478 159200 534 160000
rect 1398 159200 1454 160000
rect 2410 159200 2466 160000
rect 3330 159200 3386 160000
rect 4342 159200 4398 160000
rect 5262 159200 5318 160000
rect 6274 159200 6330 160000
rect 7286 159200 7342 160000
rect 8206 159200 8262 160000
rect 9218 159200 9274 160000
rect 10138 159200 10194 160000
rect 11150 159200 11206 160000
rect 12162 159200 12218 160000
rect 13082 159200 13138 160000
rect 14094 159200 14150 160000
rect 15014 159200 15070 160000
rect 16026 159200 16082 160000
rect 17038 159200 17094 160000
rect 17958 159200 18014 160000
rect 18970 159200 19026 160000
rect 19890 159200 19946 160000
rect 20902 159200 20958 160000
rect 21914 159200 21970 160000
rect 22834 159200 22890 160000
rect 23846 159200 23902 160000
rect 24766 159200 24822 160000
rect 25778 159200 25834 160000
rect 26790 159200 26846 160000
rect 27710 159200 27766 160000
rect 28722 159200 28778 160000
rect 29642 159200 29698 160000
rect 30654 159200 30710 160000
rect 31666 159200 31722 160000
rect 32586 159200 32642 160000
rect 33598 159200 33654 160000
rect 34518 159200 34574 160000
rect 35530 159200 35586 160000
rect 36542 159200 36598 160000
rect 37462 159200 37518 160000
rect 38474 159200 38530 160000
rect 39394 159200 39450 160000
rect 40406 159200 40462 160000
rect 41326 159200 41382 160000
rect 42338 159200 42394 160000
rect 43350 159200 43406 160000
rect 44270 159200 44326 160000
rect 45282 159200 45338 160000
rect 46202 159200 46258 160000
rect 47214 159200 47270 160000
rect 48226 159200 48282 160000
rect 49146 159200 49202 160000
rect 50158 159200 50214 160000
rect 51078 159200 51134 160000
rect 52090 159200 52146 160000
rect 53102 159200 53158 160000
rect 54022 159200 54078 160000
rect 55034 159200 55090 160000
rect 55954 159200 56010 160000
rect 56966 159200 57022 160000
rect 57978 159200 58034 160000
rect 58898 159200 58954 160000
rect 59910 159200 59966 160000
rect 60830 159200 60886 160000
rect 61842 159200 61898 160000
rect 62854 159200 62910 160000
rect 63774 159200 63830 160000
rect 64786 159200 64842 160000
rect 65706 159200 65762 160000
rect 66718 159200 66774 160000
rect 67730 159200 67786 160000
rect 68650 159200 68706 160000
rect 69662 159200 69718 160000
rect 70582 159200 70638 160000
rect 71594 159200 71650 160000
rect 72606 159200 72662 160000
rect 73526 159200 73582 160000
rect 74538 159200 74594 160000
rect 75458 159200 75514 160000
rect 76470 159200 76526 160000
rect 77482 159200 77538 160000
rect 78402 159200 78458 160000
rect 79414 159200 79470 160000
rect 80334 159200 80390 160000
rect 81346 159200 81402 160000
rect 82266 159200 82322 160000
rect 83278 159200 83334 160000
rect 84290 159200 84346 160000
rect 85210 159200 85266 160000
rect 86222 159200 86278 160000
rect 87142 159200 87198 160000
rect 88154 159200 88210 160000
rect 89166 159200 89222 160000
rect 90086 159200 90142 160000
rect 91098 159200 91154 160000
rect 92018 159200 92074 160000
rect 93030 159200 93086 160000
rect 94042 159200 94098 160000
rect 94962 159200 95018 160000
rect 95974 159200 96030 160000
rect 96894 159200 96950 160000
rect 97906 159200 97962 160000
rect 98918 159200 98974 160000
rect 99838 159200 99894 160000
rect 100850 159200 100906 160000
rect 101770 159200 101826 160000
rect 102782 159200 102838 160000
rect 103794 159200 103850 160000
rect 104714 159200 104770 160000
rect 105726 159200 105782 160000
rect 106646 159200 106702 160000
rect 107658 159200 107714 160000
rect 108670 159200 108726 160000
rect 109590 159200 109646 160000
rect 110602 159200 110658 160000
rect 111522 159200 111578 160000
rect 112534 159200 112590 160000
rect 113546 159200 113602 160000
rect 114466 159200 114522 160000
rect 115478 159200 115534 160000
rect 116398 159200 116454 160000
rect 117410 159200 117466 160000
rect 118330 159200 118386 160000
rect 119342 159200 119398 160000
rect 120354 159200 120410 160000
rect 121274 159200 121330 160000
rect 122286 159200 122342 160000
rect 123206 159200 123262 160000
rect 124218 159200 124274 160000
rect 125230 159200 125286 160000
rect 126150 159200 126206 160000
rect 127162 159200 127218 160000
rect 128082 159200 128138 160000
rect 129094 159200 129150 160000
rect 130106 159200 130162 160000
rect 131026 159200 131082 160000
rect 132038 159200 132094 160000
rect 132958 159200 133014 160000
rect 133970 159200 134026 160000
rect 134982 159200 135038 160000
rect 135902 159200 135958 160000
rect 136914 159200 136970 160000
rect 137834 159200 137890 160000
rect 138846 159200 138902 160000
rect 139858 159200 139914 160000
rect 140778 159200 140834 160000
rect 141790 159200 141846 160000
rect 142710 159200 142766 160000
rect 143722 159200 143778 160000
rect 144734 159200 144790 160000
rect 145654 159200 145710 160000
rect 146666 159200 146722 160000
rect 147586 159200 147642 160000
rect 148598 159200 148654 160000
rect 149610 159200 149666 160000
rect 150530 159200 150586 160000
rect 151542 159200 151598 160000
rect 152462 159200 152518 160000
rect 153474 159200 153530 160000
rect 154486 159200 154542 160000
rect 155406 159200 155462 160000
rect 156418 159200 156474 160000
rect 157338 159200 157394 160000
rect 158350 159200 158406 160000
rect 159270 159200 159326 160000
rect 160282 159200 160338 160000
rect 161294 159200 161350 160000
rect 162214 159200 162270 160000
rect 163226 159200 163282 160000
rect 164146 159200 164202 160000
rect 165158 159200 165214 160000
rect 166170 159200 166226 160000
rect 167090 159200 167146 160000
rect 168102 159200 168158 160000
rect 169022 159200 169078 160000
rect 170034 159200 170090 160000
rect 171046 159200 171102 160000
rect 171966 159200 172022 160000
rect 172978 159200 173034 160000
rect 173898 159200 173954 160000
rect 174910 159200 174966 160000
rect 175922 159200 175978 160000
rect 176842 159200 176898 160000
rect 177854 159200 177910 160000
rect 178774 159200 178830 160000
rect 179786 159200 179842 160000
rect 180798 159200 180854 160000
rect 181718 159200 181774 160000
rect 182730 159200 182786 160000
rect 183650 159200 183706 160000
rect 184662 159200 184718 160000
rect 185674 159200 185730 160000
rect 186594 159200 186650 160000
rect 187606 159200 187662 160000
rect 188526 159200 188582 160000
rect 189538 159200 189594 160000
rect 190550 159200 190606 160000
rect 191470 159200 191526 160000
rect 192482 159200 192538 160000
rect 193402 159200 193458 160000
rect 194414 159200 194470 160000
rect 195334 159200 195390 160000
rect 196346 159200 196402 160000
rect 197358 159200 197414 160000
rect 198278 159200 198334 160000
rect 199290 159200 199346 160000
rect 200210 159200 200266 160000
rect 201222 159200 201278 160000
rect 202234 159200 202290 160000
rect 203154 159200 203210 160000
rect 204166 159200 204222 160000
rect 205086 159200 205142 160000
rect 206098 159200 206154 160000
rect 207110 159200 207166 160000
rect 208030 159200 208086 160000
rect 209042 159200 209098 160000
rect 209962 159200 210018 160000
rect 210974 159200 211030 160000
rect 211986 159200 212042 160000
rect 212906 159200 212962 160000
rect 213918 159200 213974 160000
rect 214838 159200 214894 160000
rect 215850 159200 215906 160000
rect 216862 159200 216918 160000
rect 217782 159200 217838 160000
rect 218794 159200 218850 160000
rect 219714 159200 219770 160000
rect 220726 159200 220782 160000
rect 221738 159200 221794 160000
rect 222658 159200 222714 160000
rect 223670 159200 223726 160000
rect 224590 159200 224646 160000
rect 225602 159200 225658 160000
rect 226614 159200 226670 160000
rect 227534 159200 227590 160000
rect 228546 159200 228602 160000
rect 229466 159200 229522 160000
rect 230478 159200 230534 160000
rect 231490 159200 231546 160000
rect 232410 159200 232466 160000
rect 233422 159200 233478 160000
rect 234342 159200 234398 160000
rect 235354 159200 235410 160000
rect 236274 159200 236330 160000
rect 237286 159200 237342 160000
rect 238298 159200 238354 160000
rect 239218 159200 239274 160000
rect 240230 159200 240286 160000
rect 241150 159200 241206 160000
rect 242162 159200 242218 160000
rect 243174 159200 243230 160000
rect 244094 159200 244150 160000
rect 245106 159200 245162 160000
rect 246026 159200 246082 160000
rect 247038 159200 247094 160000
rect 248050 159200 248106 160000
rect 248970 159200 249026 160000
rect 249982 159200 250038 160000
rect 250902 159200 250958 160000
rect 251914 159200 251970 160000
rect 252926 159200 252982 160000
rect 253846 159200 253902 160000
rect 254858 159200 254914 160000
rect 255778 159200 255834 160000
rect 256790 159200 256846 160000
rect 257802 159200 257858 160000
rect 258722 159200 258778 160000
rect 259734 159200 259790 160000
rect 260654 159200 260710 160000
rect 261666 159200 261722 160000
rect 262678 159200 262734 160000
rect 263598 159200 263654 160000
rect 264610 159200 264666 160000
rect 265530 159200 265586 160000
rect 266542 159200 266598 160000
rect 267554 159200 267610 160000
rect 268474 159200 268530 160000
rect 269486 159200 269542 160000
rect 270406 159200 270462 160000
rect 271418 159200 271474 160000
rect 272338 159200 272394 160000
rect 273350 159200 273406 160000
rect 274362 159200 274418 160000
rect 275282 159200 275338 160000
rect 276294 159200 276350 160000
rect 277214 159200 277270 160000
rect 278226 159200 278282 160000
rect 279238 159200 279294 160000
rect 280158 159200 280214 160000
rect 281170 159200 281226 160000
rect 282090 159200 282146 160000
rect 283102 159200 283158 160000
rect 284114 159200 284170 160000
rect 285034 159200 285090 160000
rect 286046 159200 286102 160000
rect 286966 159200 287022 160000
rect 287978 159200 288034 160000
rect 288990 159200 289046 160000
rect 289910 159200 289966 160000
rect 290922 159200 290978 160000
rect 291842 159200 291898 160000
rect 292854 159200 292910 160000
rect 293866 159200 293922 160000
rect 294786 159200 294842 160000
rect 295798 159200 295854 160000
rect 296718 159200 296774 160000
rect 297730 159200 297786 160000
rect 298742 159200 298798 160000
rect 299662 159200 299718 160000
rect 300674 159200 300730 160000
rect 301594 159200 301650 160000
rect 302606 159200 302662 160000
rect 303618 159200 303674 160000
rect 304538 159200 304594 160000
rect 305550 159200 305606 160000
rect 306470 159200 306526 160000
rect 307482 159200 307538 160000
rect 308494 159200 308550 160000
rect 309414 159200 309470 160000
rect 310426 159200 310482 160000
rect 311346 159200 311402 160000
rect 312358 159200 312414 160000
rect 313278 159200 313334 160000
rect 314290 159200 314346 160000
rect 315302 159200 315358 160000
rect 316222 159200 316278 160000
rect 317234 159200 317290 160000
rect 318154 159200 318210 160000
rect 319166 159200 319222 160000
rect 320178 159200 320234 160000
rect 321098 159200 321154 160000
rect 322110 159200 322166 160000
rect 323030 159200 323086 160000
rect 324042 159200 324098 160000
rect 325054 159200 325110 160000
rect 325974 159200 326030 160000
rect 326986 159200 327042 160000
rect 327906 159200 327962 160000
rect 328918 159200 328974 160000
rect 329930 159200 329986 160000
rect 330850 159200 330906 160000
rect 331862 159200 331918 160000
rect 332782 159200 332838 160000
rect 333794 159200 333850 160000
rect 334806 159200 334862 160000
rect 335726 159200 335782 160000
rect 336738 159200 336794 160000
rect 337658 159200 337714 160000
rect 338670 159200 338726 160000
rect 339682 159200 339738 160000
rect 340602 159200 340658 160000
rect 341614 159200 341670 160000
rect 342534 159200 342590 160000
rect 343546 159200 343602 160000
rect 344558 159200 344614 160000
rect 345478 159200 345534 160000
rect 346490 159200 346546 160000
rect 347410 159200 347466 160000
rect 348422 159200 348478 160000
rect 349342 159200 349398 160000
rect 350354 159200 350410 160000
rect 351366 159200 351422 160000
rect 352286 159200 352342 160000
rect 353298 159200 353354 160000
rect 354218 159200 354274 160000
rect 355230 159200 355286 160000
rect 356242 159200 356298 160000
rect 357162 159200 357218 160000
rect 358174 159200 358230 160000
rect 359094 159200 359150 160000
rect 360106 159200 360162 160000
rect 361118 159200 361174 160000
rect 362038 159200 362094 160000
rect 363050 159200 363106 160000
rect 363970 159200 364026 160000
rect 364982 159200 365038 160000
rect 365994 159200 366050 160000
rect 366914 159200 366970 160000
rect 367926 159200 367982 160000
rect 368846 159200 368902 160000
rect 369858 159200 369914 160000
rect 370870 159200 370926 160000
rect 371790 159200 371846 160000
rect 372802 159200 372858 160000
rect 373722 159200 373778 160000
rect 374734 159200 374790 160000
rect 375746 159200 375802 160000
rect 376666 159200 376722 160000
rect 377678 159200 377734 160000
rect 378598 159200 378654 160000
rect 379610 159200 379666 160000
rect 380622 159200 380678 160000
rect 381542 159200 381598 160000
rect 382554 159200 382610 160000
rect 383474 159200 383530 160000
rect 384486 159200 384542 160000
rect 385498 159200 385554 160000
rect 386418 159200 386474 160000
rect 387430 159200 387486 160000
rect 388350 159200 388406 160000
rect 389362 159200 389418 160000
rect 390282 159200 390338 160000
rect 391294 159200 391350 160000
rect 392306 159200 392362 160000
rect 393226 159200 393282 160000
rect 394238 159200 394294 160000
rect 395158 159200 395214 160000
rect 396170 159200 396226 160000
rect 397182 159200 397238 160000
rect 398102 159200 398158 160000
rect 399114 159200 399170 160000
rect 400034 159200 400090 160000
rect 401046 159200 401102 160000
rect 402058 159200 402114 160000
rect 402978 159200 403034 160000
rect 403990 159200 404046 160000
rect 404910 159200 404966 160000
rect 405922 159200 405978 160000
rect 406934 159200 406990 160000
rect 407854 159200 407910 160000
rect 408866 159200 408922 160000
rect 409786 159200 409842 160000
rect 410798 159200 410854 160000
rect 411810 159200 411866 160000
rect 412730 159200 412786 160000
rect 413742 159200 413798 160000
rect 414662 159200 414718 160000
rect 415674 159200 415730 160000
rect 416686 159200 416742 160000
rect 417606 159200 417662 160000
rect 418618 159200 418674 160000
rect 419538 159200 419594 160000
rect 420550 159200 420606 160000
rect 421562 159200 421618 160000
rect 422482 159200 422538 160000
rect 423494 159200 423550 160000
rect 424414 159200 424470 160000
rect 425426 159200 425482 160000
rect 426346 159200 426402 160000
rect 427358 159200 427414 160000
rect 428370 159200 428426 160000
rect 429290 159200 429346 160000
rect 430302 159200 430358 160000
rect 431222 159200 431278 160000
rect 432234 159200 432290 160000
rect 433246 159200 433302 160000
rect 434166 159200 434222 160000
rect 435178 159200 435234 160000
rect 436098 159200 436154 160000
rect 437110 159200 437166 160000
rect 438122 159200 438178 160000
rect 439042 159200 439098 160000
rect 440054 159200 440110 160000
rect 440974 159200 441030 160000
rect 441986 159200 442042 160000
rect 442998 159200 443054 160000
rect 443918 159200 443974 160000
rect 444930 159200 444986 160000
rect 445850 159200 445906 160000
rect 446862 159200 446918 160000
rect 447874 159200 447930 160000
rect 448794 159200 448850 160000
rect 449806 159200 449862 160000
rect 450726 159200 450782 160000
rect 451738 159200 451794 160000
rect 452750 159200 452806 160000
rect 453670 159200 453726 160000
rect 454682 159200 454738 160000
rect 455602 159200 455658 160000
rect 456614 159200 456670 160000
rect 457626 159200 457682 160000
rect 458546 159200 458602 160000
rect 459558 159200 459614 160000
rect 460478 159200 460534 160000
rect 461490 159200 461546 160000
rect 462502 159200 462558 160000
rect 463422 159200 463478 160000
rect 464434 159200 464490 160000
rect 465354 159200 465410 160000
rect 466366 159200 466422 160000
rect 467286 159200 467342 160000
rect 468298 159200 468354 160000
rect 469310 159200 469366 160000
rect 470230 159200 470286 160000
rect 471242 159200 471298 160000
rect 472162 159200 472218 160000
rect 473174 159200 473230 160000
rect 474186 159200 474242 160000
rect 475106 159200 475162 160000
rect 476118 159200 476174 160000
rect 477038 159200 477094 160000
rect 478050 159200 478106 160000
rect 479062 159200 479118 160000
rect 479982 159200 480038 160000
rect 480994 159200 481050 160000
rect 481914 159200 481970 160000
rect 482926 159200 482982 160000
rect 483938 159200 483994 160000
rect 484858 159200 484914 160000
rect 485870 159200 485926 160000
rect 486790 159200 486846 160000
rect 487802 159200 487858 160000
rect 488814 159200 488870 160000
rect 489734 159200 489790 160000
rect 490746 159200 490802 160000
rect 491666 159200 491722 160000
rect 492678 159200 492734 160000
rect 493690 159200 493746 160000
rect 494610 159200 494666 160000
rect 495622 159200 495678 160000
rect 496542 159200 496598 160000
rect 497554 159200 497610 160000
rect 498566 159200 498622 160000
rect 499486 159200 499542 160000
rect 500498 159200 500554 160000
rect 501418 159200 501474 160000
rect 502430 159200 502486 160000
rect 503350 159200 503406 160000
rect 504362 159200 504418 160000
rect 505374 159200 505430 160000
rect 506294 159200 506350 160000
rect 507306 159200 507362 160000
rect 508226 159200 508282 160000
rect 509238 159200 509294 160000
rect 510250 159200 510306 160000
rect 511170 159200 511226 160000
rect 512182 159200 512238 160000
rect 513102 159200 513158 160000
rect 514114 159200 514170 160000
rect 515126 159200 515182 160000
rect 516046 159200 516102 160000
rect 517058 159200 517114 160000
rect 517978 159200 518034 160000
rect 518990 159200 519046 160000
rect 520002 159200 520058 160000
rect 520922 159200 520978 160000
rect 521934 159200 521990 160000
rect 522854 159200 522910 160000
rect 523866 159200 523922 160000
rect 524878 159200 524934 160000
rect 525798 159200 525854 160000
rect 526810 159200 526866 160000
rect 527730 159200 527786 160000
rect 528742 159200 528798 160000
rect 529754 159200 529810 160000
rect 530674 159200 530730 160000
rect 531686 159200 531742 160000
rect 532606 159200 532662 160000
rect 533618 159200 533674 160000
rect 534630 159200 534686 160000
rect 535550 159200 535606 160000
rect 536562 159200 536618 160000
rect 537482 159200 537538 160000
rect 538494 159200 538550 160000
rect 539506 159200 539562 160000
rect 540426 159200 540482 160000
rect 541438 159200 541494 160000
rect 542358 159200 542414 160000
rect 543370 159200 543426 160000
rect 544290 159200 544346 160000
rect 545302 159200 545358 160000
rect 546314 159200 546370 160000
rect 547234 159200 547290 160000
rect 548246 159200 548302 160000
rect 549166 159200 549222 160000
rect 550178 159200 550234 160000
rect 551190 159200 551246 160000
rect 552110 159200 552166 160000
rect 553122 159200 553178 160000
rect 554042 159200 554098 160000
rect 555054 159200 555110 160000
rect 556066 159200 556122 160000
rect 556986 159200 557042 160000
rect 557998 159200 558054 160000
rect 558918 159200 558974 160000
rect 559930 159200 559986 160000
rect 560942 159200 560998 160000
rect 561862 159200 561918 160000
rect 562874 159200 562930 160000
rect 563794 159200 563850 160000
rect 564806 159200 564862 160000
rect 565818 159200 565874 160000
rect 566738 159200 566794 160000
rect 567750 159200 567806 160000
rect 568670 159200 568726 160000
rect 569682 159200 569738 160000
rect 570694 159200 570750 160000
rect 571614 159200 571670 160000
rect 572626 159200 572682 160000
rect 573546 159200 573602 160000
rect 574558 159200 574614 160000
rect 575570 159200 575626 160000
rect 576490 159200 576546 160000
rect 577502 159200 577558 160000
rect 578422 159200 578478 160000
rect 579434 159200 579490 160000
rect 2594 0 2650 800
rect 7838 0 7894 800
rect 13174 0 13230 800
rect 18510 0 18566 800
rect 23846 0 23902 800
rect 29182 0 29238 800
rect 34518 0 34574 800
rect 39762 0 39818 800
rect 45098 0 45154 800
rect 50434 0 50490 800
rect 55770 0 55826 800
rect 61106 0 61162 800
rect 66442 0 66498 800
rect 71686 0 71742 800
rect 77022 0 77078 800
rect 82358 0 82414 800
rect 87694 0 87750 800
rect 93030 0 93086 800
rect 98366 0 98422 800
rect 103610 0 103666 800
rect 108946 0 109002 800
rect 114282 0 114338 800
rect 119618 0 119674 800
rect 124954 0 125010 800
rect 130290 0 130346 800
rect 135534 0 135590 800
rect 140870 0 140926 800
rect 146206 0 146262 800
rect 151542 0 151598 800
rect 156878 0 156934 800
rect 162214 0 162270 800
rect 167458 0 167514 800
rect 172794 0 172850 800
rect 178130 0 178186 800
rect 183466 0 183522 800
rect 188802 0 188858 800
rect 194138 0 194194 800
rect 199382 0 199438 800
rect 204718 0 204774 800
rect 210054 0 210110 800
rect 215390 0 215446 800
rect 220726 0 220782 800
rect 226062 0 226118 800
rect 231306 0 231362 800
rect 236642 0 236698 800
rect 241978 0 242034 800
rect 247314 0 247370 800
rect 252650 0 252706 800
rect 257986 0 258042 800
rect 263230 0 263286 800
rect 268566 0 268622 800
rect 273902 0 273958 800
rect 279238 0 279294 800
rect 284574 0 284630 800
rect 289910 0 289966 800
rect 295154 0 295210 800
rect 300490 0 300546 800
rect 305826 0 305882 800
rect 311162 0 311218 800
rect 316498 0 316554 800
rect 321834 0 321890 800
rect 327078 0 327134 800
rect 332414 0 332470 800
rect 337750 0 337806 800
rect 343086 0 343142 800
rect 348422 0 348478 800
rect 353758 0 353814 800
rect 359002 0 359058 800
rect 364338 0 364394 800
rect 369674 0 369730 800
rect 375010 0 375066 800
rect 380346 0 380402 800
rect 385682 0 385738 800
rect 390926 0 390982 800
rect 396262 0 396318 800
rect 401598 0 401654 800
rect 406934 0 406990 800
rect 412270 0 412326 800
rect 417606 0 417662 800
rect 422850 0 422906 800
rect 428186 0 428242 800
rect 433522 0 433578 800
rect 438858 0 438914 800
rect 444194 0 444250 800
rect 449530 0 449586 800
rect 454774 0 454830 800
rect 460110 0 460166 800
rect 465446 0 465502 800
rect 470782 0 470838 800
rect 476118 0 476174 800
rect 481454 0 481510 800
rect 486698 0 486754 800
rect 492034 0 492090 800
rect 497370 0 497426 800
rect 502706 0 502762 800
rect 508042 0 508098 800
rect 513378 0 513434 800
rect 518622 0 518678 800
rect 523958 0 524014 800
rect 529294 0 529350 800
rect 534630 0 534686 800
rect 539966 0 540022 800
rect 545302 0 545358 800
rect 550546 0 550602 800
rect 555882 0 555938 800
rect 561218 0 561274 800
rect 566554 0 566610 800
rect 571890 0 571946 800
rect 577226 0 577282 800
<< obsm2 >>
rect 590 159144 1342 159338
rect 1510 159144 2354 159338
rect 2522 159144 3274 159338
rect 3442 159144 4286 159338
rect 4454 159144 5206 159338
rect 5374 159144 6218 159338
rect 6386 159144 7230 159338
rect 7398 159144 8150 159338
rect 8318 159144 9162 159338
rect 9330 159144 10082 159338
rect 10250 159144 11094 159338
rect 11262 159144 12106 159338
rect 12274 159144 13026 159338
rect 13194 159144 14038 159338
rect 14206 159144 14958 159338
rect 15126 159144 15970 159338
rect 16138 159144 16982 159338
rect 17150 159144 17902 159338
rect 18070 159144 18914 159338
rect 19082 159144 19834 159338
rect 20002 159144 20846 159338
rect 21014 159144 21858 159338
rect 22026 159144 22778 159338
rect 22946 159144 23790 159338
rect 23958 159144 24710 159338
rect 24878 159144 25722 159338
rect 25890 159144 26734 159338
rect 26902 159144 27654 159338
rect 27822 159144 28666 159338
rect 28834 159144 29586 159338
rect 29754 159144 30598 159338
rect 30766 159144 31610 159338
rect 31778 159144 32530 159338
rect 32698 159144 33542 159338
rect 33710 159144 34462 159338
rect 34630 159144 35474 159338
rect 35642 159144 36486 159338
rect 36654 159144 37406 159338
rect 37574 159144 38418 159338
rect 38586 159144 39338 159338
rect 39506 159144 40350 159338
rect 40518 159144 41270 159338
rect 41438 159144 42282 159338
rect 42450 159144 43294 159338
rect 43462 159144 44214 159338
rect 44382 159144 45226 159338
rect 45394 159144 46146 159338
rect 46314 159144 47158 159338
rect 47326 159144 48170 159338
rect 48338 159144 49090 159338
rect 49258 159144 50102 159338
rect 50270 159144 51022 159338
rect 51190 159144 52034 159338
rect 52202 159144 53046 159338
rect 53214 159144 53966 159338
rect 54134 159144 54978 159338
rect 55146 159144 55898 159338
rect 56066 159144 56910 159338
rect 57078 159144 57922 159338
rect 58090 159144 58842 159338
rect 59010 159144 59854 159338
rect 60022 159144 60774 159338
rect 60942 159144 61786 159338
rect 61954 159144 62798 159338
rect 62966 159144 63718 159338
rect 63886 159144 64730 159338
rect 64898 159144 65650 159338
rect 65818 159144 66662 159338
rect 66830 159144 67674 159338
rect 67842 159144 68594 159338
rect 68762 159144 69606 159338
rect 69774 159144 70526 159338
rect 70694 159144 71538 159338
rect 71706 159144 72550 159338
rect 72718 159144 73470 159338
rect 73638 159144 74482 159338
rect 74650 159144 75402 159338
rect 75570 159144 76414 159338
rect 76582 159144 77426 159338
rect 77594 159144 78346 159338
rect 78514 159144 79358 159338
rect 79526 159144 80278 159338
rect 80446 159144 81290 159338
rect 81458 159144 82210 159338
rect 82378 159144 83222 159338
rect 83390 159144 84234 159338
rect 84402 159144 85154 159338
rect 85322 159144 86166 159338
rect 86334 159144 87086 159338
rect 87254 159144 88098 159338
rect 88266 159144 89110 159338
rect 89278 159144 90030 159338
rect 90198 159144 91042 159338
rect 91210 159144 91962 159338
rect 92130 159144 92974 159338
rect 93142 159144 93986 159338
rect 94154 159144 94906 159338
rect 95074 159144 95918 159338
rect 96086 159144 96838 159338
rect 97006 159144 97850 159338
rect 98018 159144 98862 159338
rect 99030 159144 99782 159338
rect 99950 159144 100794 159338
rect 100962 159144 101714 159338
rect 101882 159144 102726 159338
rect 102894 159144 103738 159338
rect 103906 159144 104658 159338
rect 104826 159144 105670 159338
rect 105838 159144 106590 159338
rect 106758 159144 107602 159338
rect 107770 159144 108614 159338
rect 108782 159144 109534 159338
rect 109702 159144 110546 159338
rect 110714 159144 111466 159338
rect 111634 159144 112478 159338
rect 112646 159144 113490 159338
rect 113658 159144 114410 159338
rect 114578 159144 115422 159338
rect 115590 159144 116342 159338
rect 116510 159144 117354 159338
rect 117522 159144 118274 159338
rect 118442 159144 119286 159338
rect 119454 159144 120298 159338
rect 120466 159144 121218 159338
rect 121386 159144 122230 159338
rect 122398 159144 123150 159338
rect 123318 159144 124162 159338
rect 124330 159144 125174 159338
rect 125342 159144 126094 159338
rect 126262 159144 127106 159338
rect 127274 159144 128026 159338
rect 128194 159144 129038 159338
rect 129206 159144 130050 159338
rect 130218 159144 130970 159338
rect 131138 159144 131982 159338
rect 132150 159144 132902 159338
rect 133070 159144 133914 159338
rect 134082 159144 134926 159338
rect 135094 159144 135846 159338
rect 136014 159144 136858 159338
rect 137026 159144 137778 159338
rect 137946 159144 138790 159338
rect 138958 159144 139802 159338
rect 139970 159144 140722 159338
rect 140890 159144 141734 159338
rect 141902 159144 142654 159338
rect 142822 159144 143666 159338
rect 143834 159144 144678 159338
rect 144846 159144 145598 159338
rect 145766 159144 146610 159338
rect 146778 159144 147530 159338
rect 147698 159144 148542 159338
rect 148710 159144 149554 159338
rect 149722 159144 150474 159338
rect 150642 159144 151486 159338
rect 151654 159144 152406 159338
rect 152574 159144 153418 159338
rect 153586 159144 154430 159338
rect 154598 159144 155350 159338
rect 155518 159144 156362 159338
rect 156530 159144 157282 159338
rect 157450 159144 158294 159338
rect 158462 159144 159214 159338
rect 159382 159144 160226 159338
rect 160394 159144 161238 159338
rect 161406 159144 162158 159338
rect 162326 159144 163170 159338
rect 163338 159144 164090 159338
rect 164258 159144 165102 159338
rect 165270 159144 166114 159338
rect 166282 159144 167034 159338
rect 167202 159144 168046 159338
rect 168214 159144 168966 159338
rect 169134 159144 169978 159338
rect 170146 159144 170990 159338
rect 171158 159144 171910 159338
rect 172078 159144 172922 159338
rect 173090 159144 173842 159338
rect 174010 159144 174854 159338
rect 175022 159144 175866 159338
rect 176034 159144 176786 159338
rect 176954 159144 177798 159338
rect 177966 159144 178718 159338
rect 178886 159144 179730 159338
rect 179898 159144 180742 159338
rect 180910 159144 181662 159338
rect 181830 159144 182674 159338
rect 182842 159144 183594 159338
rect 183762 159144 184606 159338
rect 184774 159144 185618 159338
rect 185786 159144 186538 159338
rect 186706 159144 187550 159338
rect 187718 159144 188470 159338
rect 188638 159144 189482 159338
rect 189650 159144 190494 159338
rect 190662 159144 191414 159338
rect 191582 159144 192426 159338
rect 192594 159144 193346 159338
rect 193514 159144 194358 159338
rect 194526 159144 195278 159338
rect 195446 159144 196290 159338
rect 196458 159144 197302 159338
rect 197470 159144 198222 159338
rect 198390 159144 199234 159338
rect 199402 159144 200154 159338
rect 200322 159144 201166 159338
rect 201334 159144 202178 159338
rect 202346 159144 203098 159338
rect 203266 159144 204110 159338
rect 204278 159144 205030 159338
rect 205198 159144 206042 159338
rect 206210 159144 207054 159338
rect 207222 159144 207974 159338
rect 208142 159144 208986 159338
rect 209154 159144 209906 159338
rect 210074 159144 210918 159338
rect 211086 159144 211930 159338
rect 212098 159144 212850 159338
rect 213018 159144 213862 159338
rect 214030 159144 214782 159338
rect 214950 159144 215794 159338
rect 215962 159144 216806 159338
rect 216974 159144 217726 159338
rect 217894 159144 218738 159338
rect 218906 159144 219658 159338
rect 219826 159144 220670 159338
rect 220838 159144 221682 159338
rect 221850 159144 222602 159338
rect 222770 159144 223614 159338
rect 223782 159144 224534 159338
rect 224702 159144 225546 159338
rect 225714 159144 226558 159338
rect 226726 159144 227478 159338
rect 227646 159144 228490 159338
rect 228658 159144 229410 159338
rect 229578 159144 230422 159338
rect 230590 159144 231434 159338
rect 231602 159144 232354 159338
rect 232522 159144 233366 159338
rect 233534 159144 234286 159338
rect 234454 159144 235298 159338
rect 235466 159144 236218 159338
rect 236386 159144 237230 159338
rect 237398 159144 238242 159338
rect 238410 159144 239162 159338
rect 239330 159144 240174 159338
rect 240342 159144 241094 159338
rect 241262 159144 242106 159338
rect 242274 159144 243118 159338
rect 243286 159144 244038 159338
rect 244206 159144 245050 159338
rect 245218 159144 245970 159338
rect 246138 159144 246982 159338
rect 247150 159144 247994 159338
rect 248162 159144 248914 159338
rect 249082 159144 249926 159338
rect 250094 159144 250846 159338
rect 251014 159144 251858 159338
rect 252026 159144 252870 159338
rect 253038 159144 253790 159338
rect 253958 159144 254802 159338
rect 254970 159144 255722 159338
rect 255890 159144 256734 159338
rect 256902 159144 257746 159338
rect 257914 159144 258666 159338
rect 258834 159144 259678 159338
rect 259846 159144 260598 159338
rect 260766 159144 261610 159338
rect 261778 159144 262622 159338
rect 262790 159144 263542 159338
rect 263710 159144 264554 159338
rect 264722 159144 265474 159338
rect 265642 159144 266486 159338
rect 266654 159144 267498 159338
rect 267666 159144 268418 159338
rect 268586 159144 269430 159338
rect 269598 159144 270350 159338
rect 270518 159144 271362 159338
rect 271530 159144 272282 159338
rect 272450 159144 273294 159338
rect 273462 159144 274306 159338
rect 274474 159144 275226 159338
rect 275394 159144 276238 159338
rect 276406 159144 277158 159338
rect 277326 159144 278170 159338
rect 278338 159144 279182 159338
rect 279350 159144 280102 159338
rect 280270 159144 281114 159338
rect 281282 159144 282034 159338
rect 282202 159144 283046 159338
rect 283214 159144 284058 159338
rect 284226 159144 284978 159338
rect 285146 159144 285990 159338
rect 286158 159144 286910 159338
rect 287078 159144 287922 159338
rect 288090 159144 288934 159338
rect 289102 159144 289854 159338
rect 290022 159144 290866 159338
rect 291034 159144 291786 159338
rect 291954 159144 292798 159338
rect 292966 159144 293810 159338
rect 293978 159144 294730 159338
rect 294898 159144 295742 159338
rect 295910 159144 296662 159338
rect 296830 159144 297674 159338
rect 297842 159144 298686 159338
rect 298854 159144 299606 159338
rect 299774 159144 300618 159338
rect 300786 159144 301538 159338
rect 301706 159144 302550 159338
rect 302718 159144 303562 159338
rect 303730 159144 304482 159338
rect 304650 159144 305494 159338
rect 305662 159144 306414 159338
rect 306582 159144 307426 159338
rect 307594 159144 308438 159338
rect 308606 159144 309358 159338
rect 309526 159144 310370 159338
rect 310538 159144 311290 159338
rect 311458 159144 312302 159338
rect 312470 159144 313222 159338
rect 313390 159144 314234 159338
rect 314402 159144 315246 159338
rect 315414 159144 316166 159338
rect 316334 159144 317178 159338
rect 317346 159144 318098 159338
rect 318266 159144 319110 159338
rect 319278 159144 320122 159338
rect 320290 159144 321042 159338
rect 321210 159144 322054 159338
rect 322222 159144 322974 159338
rect 323142 159144 323986 159338
rect 324154 159144 324998 159338
rect 325166 159144 325918 159338
rect 326086 159144 326930 159338
rect 327098 159144 327850 159338
rect 328018 159144 328862 159338
rect 329030 159144 329874 159338
rect 330042 159144 330794 159338
rect 330962 159144 331806 159338
rect 331974 159144 332726 159338
rect 332894 159144 333738 159338
rect 333906 159144 334750 159338
rect 334918 159144 335670 159338
rect 335838 159144 336682 159338
rect 336850 159144 337602 159338
rect 337770 159144 338614 159338
rect 338782 159144 339626 159338
rect 339794 159144 340546 159338
rect 340714 159144 341558 159338
rect 341726 159144 342478 159338
rect 342646 159144 343490 159338
rect 343658 159144 344502 159338
rect 344670 159144 345422 159338
rect 345590 159144 346434 159338
rect 346602 159144 347354 159338
rect 347522 159144 348366 159338
rect 348534 159144 349286 159338
rect 349454 159144 350298 159338
rect 350466 159144 351310 159338
rect 351478 159144 352230 159338
rect 352398 159144 353242 159338
rect 353410 159144 354162 159338
rect 354330 159144 355174 159338
rect 355342 159144 356186 159338
rect 356354 159144 357106 159338
rect 357274 159144 358118 159338
rect 358286 159144 359038 159338
rect 359206 159144 360050 159338
rect 360218 159144 361062 159338
rect 361230 159144 361982 159338
rect 362150 159144 362994 159338
rect 363162 159144 363914 159338
rect 364082 159144 364926 159338
rect 365094 159144 365938 159338
rect 366106 159144 366858 159338
rect 367026 159144 367870 159338
rect 368038 159144 368790 159338
rect 368958 159144 369802 159338
rect 369970 159144 370814 159338
rect 370982 159144 371734 159338
rect 371902 159144 372746 159338
rect 372914 159144 373666 159338
rect 373834 159144 374678 159338
rect 374846 159144 375690 159338
rect 375858 159144 376610 159338
rect 376778 159144 377622 159338
rect 377790 159144 378542 159338
rect 378710 159144 379554 159338
rect 379722 159144 380566 159338
rect 380734 159144 381486 159338
rect 381654 159144 382498 159338
rect 382666 159144 383418 159338
rect 383586 159144 384430 159338
rect 384598 159144 385442 159338
rect 385610 159144 386362 159338
rect 386530 159144 387374 159338
rect 387542 159144 388294 159338
rect 388462 159144 389306 159338
rect 389474 159144 390226 159338
rect 390394 159144 391238 159338
rect 391406 159144 392250 159338
rect 392418 159144 393170 159338
rect 393338 159144 394182 159338
rect 394350 159144 395102 159338
rect 395270 159144 396114 159338
rect 396282 159144 397126 159338
rect 397294 159144 398046 159338
rect 398214 159144 399058 159338
rect 399226 159144 399978 159338
rect 400146 159144 400990 159338
rect 401158 159144 402002 159338
rect 402170 159144 402922 159338
rect 403090 159144 403934 159338
rect 404102 159144 404854 159338
rect 405022 159144 405866 159338
rect 406034 159144 406878 159338
rect 407046 159144 407798 159338
rect 407966 159144 408810 159338
rect 408978 159144 409730 159338
rect 409898 159144 410742 159338
rect 410910 159144 411754 159338
rect 411922 159144 412674 159338
rect 412842 159144 413686 159338
rect 413854 159144 414606 159338
rect 414774 159144 415618 159338
rect 415786 159144 416630 159338
rect 416798 159144 417550 159338
rect 417718 159144 418562 159338
rect 418730 159144 419482 159338
rect 419650 159144 420494 159338
rect 420662 159144 421506 159338
rect 421674 159144 422426 159338
rect 422594 159144 423438 159338
rect 423606 159144 424358 159338
rect 424526 159144 425370 159338
rect 425538 159144 426290 159338
rect 426458 159144 427302 159338
rect 427470 159144 428314 159338
rect 428482 159144 429234 159338
rect 429402 159144 430246 159338
rect 430414 159144 431166 159338
rect 431334 159144 432178 159338
rect 432346 159144 433190 159338
rect 433358 159144 434110 159338
rect 434278 159144 435122 159338
rect 435290 159144 436042 159338
rect 436210 159144 437054 159338
rect 437222 159144 438066 159338
rect 438234 159144 438986 159338
rect 439154 159144 439998 159338
rect 440166 159144 440918 159338
rect 441086 159144 441930 159338
rect 442098 159144 442942 159338
rect 443110 159144 443862 159338
rect 444030 159144 444874 159338
rect 445042 159144 445794 159338
rect 445962 159144 446806 159338
rect 446974 159144 447818 159338
rect 447986 159144 448738 159338
rect 448906 159144 449750 159338
rect 449918 159144 450670 159338
rect 450838 159144 451682 159338
rect 451850 159144 452694 159338
rect 452862 159144 453614 159338
rect 453782 159144 454626 159338
rect 454794 159144 455546 159338
rect 455714 159144 456558 159338
rect 456726 159144 457570 159338
rect 457738 159144 458490 159338
rect 458658 159144 459502 159338
rect 459670 159144 460422 159338
rect 460590 159144 461434 159338
rect 461602 159144 462446 159338
rect 462614 159144 463366 159338
rect 463534 159144 464378 159338
rect 464546 159144 465298 159338
rect 465466 159144 466310 159338
rect 466478 159144 467230 159338
rect 467398 159144 468242 159338
rect 468410 159144 469254 159338
rect 469422 159144 470174 159338
rect 470342 159144 471186 159338
rect 471354 159144 472106 159338
rect 472274 159144 473118 159338
rect 473286 159144 474130 159338
rect 474298 159144 475050 159338
rect 475218 159144 476062 159338
rect 476230 159144 476982 159338
rect 477150 159144 477994 159338
rect 478162 159144 479006 159338
rect 479174 159144 479926 159338
rect 480094 159144 480938 159338
rect 481106 159144 481858 159338
rect 482026 159144 482870 159338
rect 483038 159144 483882 159338
rect 484050 159144 484802 159338
rect 484970 159144 485814 159338
rect 485982 159144 486734 159338
rect 486902 159144 487746 159338
rect 487914 159144 488758 159338
rect 488926 159144 489678 159338
rect 489846 159144 490690 159338
rect 490858 159144 491610 159338
rect 491778 159144 492622 159338
rect 492790 159144 493634 159338
rect 493802 159144 494554 159338
rect 494722 159144 495566 159338
rect 495734 159144 496486 159338
rect 496654 159144 497498 159338
rect 497666 159144 498510 159338
rect 498678 159144 499430 159338
rect 499598 159144 500442 159338
rect 500610 159144 501362 159338
rect 501530 159144 502374 159338
rect 502542 159144 503294 159338
rect 503462 159144 504306 159338
rect 504474 159144 505318 159338
rect 505486 159144 506238 159338
rect 506406 159144 507250 159338
rect 507418 159144 508170 159338
rect 508338 159144 509182 159338
rect 509350 159144 510194 159338
rect 510362 159144 511114 159338
rect 511282 159144 512126 159338
rect 512294 159144 513046 159338
rect 513214 159144 514058 159338
rect 514226 159144 515070 159338
rect 515238 159144 515990 159338
rect 516158 159144 517002 159338
rect 517170 159144 517922 159338
rect 518090 159144 518934 159338
rect 519102 159144 519946 159338
rect 520114 159144 520866 159338
rect 521034 159144 521878 159338
rect 522046 159144 522798 159338
rect 522966 159144 523810 159338
rect 523978 159144 524822 159338
rect 524990 159144 525742 159338
rect 525910 159144 526754 159338
rect 526922 159144 527674 159338
rect 527842 159144 528686 159338
rect 528854 159144 529698 159338
rect 529866 159144 530618 159338
rect 530786 159144 531630 159338
rect 531798 159144 532550 159338
rect 532718 159144 533562 159338
rect 533730 159144 534574 159338
rect 534742 159144 535494 159338
rect 535662 159144 536506 159338
rect 536674 159144 537426 159338
rect 537594 159144 538438 159338
rect 538606 159144 539450 159338
rect 539618 159144 540370 159338
rect 540538 159144 541382 159338
rect 541550 159144 542302 159338
rect 542470 159144 543314 159338
rect 543482 159144 544234 159338
rect 544402 159144 545246 159338
rect 545414 159144 546258 159338
rect 546426 159144 547178 159338
rect 547346 159144 548190 159338
rect 548358 159144 549110 159338
rect 549278 159144 550122 159338
rect 550290 159144 551134 159338
rect 551302 159144 552054 159338
rect 552222 159144 553066 159338
rect 553234 159144 553986 159338
rect 554154 159144 554998 159338
rect 555166 159144 556010 159338
rect 556178 159144 556930 159338
rect 557098 159144 557942 159338
rect 558110 159144 558862 159338
rect 559030 159144 559874 159338
rect 560042 159144 560886 159338
rect 561054 159144 561806 159338
rect 561974 159144 562818 159338
rect 562986 159144 563738 159338
rect 563906 159144 564750 159338
rect 564918 159144 565762 159338
rect 565930 159144 566682 159338
rect 566850 159144 567694 159338
rect 567862 159144 568614 159338
rect 568782 159144 569626 159338
rect 569794 159144 570638 159338
rect 570806 159144 571558 159338
rect 571726 159144 572570 159338
rect 572738 159144 573490 159338
rect 573658 159144 574502 159338
rect 574670 159144 575514 159338
rect 575682 159144 576434 159338
rect 576602 159144 577446 159338
rect 577614 159144 578366 159338
rect 578534 159144 579378 159338
rect 480 856 579490 159144
rect 480 734 2538 856
rect 2706 734 7782 856
rect 7950 734 13118 856
rect 13286 734 18454 856
rect 18622 734 23790 856
rect 23958 734 29126 856
rect 29294 734 34462 856
rect 34630 734 39706 856
rect 39874 734 45042 856
rect 45210 734 50378 856
rect 50546 734 55714 856
rect 55882 734 61050 856
rect 61218 734 66386 856
rect 66554 734 71630 856
rect 71798 734 76966 856
rect 77134 734 82302 856
rect 82470 734 87638 856
rect 87806 734 92974 856
rect 93142 734 98310 856
rect 98478 734 103554 856
rect 103722 734 108890 856
rect 109058 734 114226 856
rect 114394 734 119562 856
rect 119730 734 124898 856
rect 125066 734 130234 856
rect 130402 734 135478 856
rect 135646 734 140814 856
rect 140982 734 146150 856
rect 146318 734 151486 856
rect 151654 734 156822 856
rect 156990 734 162158 856
rect 162326 734 167402 856
rect 167570 734 172738 856
rect 172906 734 178074 856
rect 178242 734 183410 856
rect 183578 734 188746 856
rect 188914 734 194082 856
rect 194250 734 199326 856
rect 199494 734 204662 856
rect 204830 734 209998 856
rect 210166 734 215334 856
rect 215502 734 220670 856
rect 220838 734 226006 856
rect 226174 734 231250 856
rect 231418 734 236586 856
rect 236754 734 241922 856
rect 242090 734 247258 856
rect 247426 734 252594 856
rect 252762 734 257930 856
rect 258098 734 263174 856
rect 263342 734 268510 856
rect 268678 734 273846 856
rect 274014 734 279182 856
rect 279350 734 284518 856
rect 284686 734 289854 856
rect 290022 734 295098 856
rect 295266 734 300434 856
rect 300602 734 305770 856
rect 305938 734 311106 856
rect 311274 734 316442 856
rect 316610 734 321778 856
rect 321946 734 327022 856
rect 327190 734 332358 856
rect 332526 734 337694 856
rect 337862 734 343030 856
rect 343198 734 348366 856
rect 348534 734 353702 856
rect 353870 734 358946 856
rect 359114 734 364282 856
rect 364450 734 369618 856
rect 369786 734 374954 856
rect 375122 734 380290 856
rect 380458 734 385626 856
rect 385794 734 390870 856
rect 391038 734 396206 856
rect 396374 734 401542 856
rect 401710 734 406878 856
rect 407046 734 412214 856
rect 412382 734 417550 856
rect 417718 734 422794 856
rect 422962 734 428130 856
rect 428298 734 433466 856
rect 433634 734 438802 856
rect 438970 734 444138 856
rect 444306 734 449474 856
rect 449642 734 454718 856
rect 454886 734 460054 856
rect 460222 734 465390 856
rect 465558 734 470726 856
rect 470894 734 476062 856
rect 476230 734 481398 856
rect 481566 734 486642 856
rect 486810 734 491978 856
rect 492146 734 497314 856
rect 497482 734 502650 856
rect 502818 734 507986 856
rect 508154 734 513322 856
rect 513490 734 518566 856
rect 518734 734 523902 856
rect 524070 734 529238 856
rect 529406 734 534574 856
rect 534742 734 539910 856
rect 540078 734 545246 856
rect 545414 734 550490 856
rect 550658 734 555826 856
rect 555994 734 561162 856
rect 561330 734 566498 856
rect 566666 734 571834 856
rect 572002 734 577170 856
rect 577338 734 579490 856
<< metal3 >>
rect 0 157496 800 157616
rect 0 152872 800 152992
rect 0 148384 800 148504
rect 0 143760 800 143880
rect 0 139272 800 139392
rect 0 134648 800 134768
rect 0 130024 800 130144
rect 0 125536 800 125656
rect 0 120912 800 121032
rect 0 116424 800 116544
rect 0 111800 800 111920
rect 0 107176 800 107296
rect 0 102688 800 102808
rect 0 98064 800 98184
rect 0 93576 800 93696
rect 0 88952 800 89072
rect 0 84328 800 84448
rect 0 79840 800 79960
rect 0 75216 800 75336
rect 0 70728 800 70848
rect 0 66104 800 66224
rect 0 61480 800 61600
rect 0 56992 800 57112
rect 0 52368 800 52488
rect 0 47880 800 48000
rect 0 43256 800 43376
rect 0 38632 800 38752
rect 0 34144 800 34264
rect 0 29520 800 29640
rect 0 25032 800 25152
rect 0 20408 800 20528
rect 0 15784 800 15904
rect 0 11296 800 11416
rect 0 6672 800 6792
rect 0 2184 800 2304
<< obsm3 >>
rect 880 157416 579495 157589
rect 800 153072 579495 157416
rect 880 152792 579495 153072
rect 800 148584 579495 152792
rect 880 148304 579495 148584
rect 800 143960 579495 148304
rect 880 143680 579495 143960
rect 800 139472 579495 143680
rect 880 139192 579495 139472
rect 800 134848 579495 139192
rect 880 134568 579495 134848
rect 800 130224 579495 134568
rect 880 129944 579495 130224
rect 800 125736 579495 129944
rect 880 125456 579495 125736
rect 800 121112 579495 125456
rect 880 120832 579495 121112
rect 800 116624 579495 120832
rect 880 116344 579495 116624
rect 800 112000 579495 116344
rect 880 111720 579495 112000
rect 800 107376 579495 111720
rect 880 107096 579495 107376
rect 800 102888 579495 107096
rect 880 102608 579495 102888
rect 800 98264 579495 102608
rect 880 97984 579495 98264
rect 800 93776 579495 97984
rect 880 93496 579495 93776
rect 800 89152 579495 93496
rect 880 88872 579495 89152
rect 800 84528 579495 88872
rect 880 84248 579495 84528
rect 800 80040 579495 84248
rect 880 79760 579495 80040
rect 800 75416 579495 79760
rect 880 75136 579495 75416
rect 800 70928 579495 75136
rect 880 70648 579495 70928
rect 800 66304 579495 70648
rect 880 66024 579495 66304
rect 800 61680 579495 66024
rect 880 61400 579495 61680
rect 800 57192 579495 61400
rect 880 56912 579495 57192
rect 800 52568 579495 56912
rect 880 52288 579495 52568
rect 800 48080 579495 52288
rect 880 47800 579495 48080
rect 800 43456 579495 47800
rect 880 43176 579495 43456
rect 800 38832 579495 43176
rect 880 38552 579495 38832
rect 800 34344 579495 38552
rect 880 34064 579495 34344
rect 800 29720 579495 34064
rect 880 29440 579495 29720
rect 800 25232 579495 29440
rect 880 24952 579495 25232
rect 800 20608 579495 24952
rect 880 20328 579495 20608
rect 800 15984 579495 20328
rect 880 15704 579495 15984
rect 800 11496 579495 15704
rect 880 11216 579495 11496
rect 800 6872 579495 11216
rect 880 6592 579495 6872
rect 800 2384 579495 6592
rect 880 2104 579495 2384
rect 800 1803 579495 2104
<< metal4 >>
rect 4208 154000 4528 157760
rect 9208 154000 9528 157760
rect 14208 154000 14528 157760
rect 19208 154000 19528 157760
rect 24208 154000 24528 157760
rect 29208 154000 29528 157760
rect 34208 154000 34528 157760
rect 39208 154000 39528 157760
rect 44208 154000 44528 157760
rect 49208 154000 49528 157760
rect 54208 154000 54528 157760
rect 59208 154000 59528 157760
rect 64208 154000 64528 157760
rect 69208 154000 69528 157760
rect 74208 154000 74528 157760
rect 79208 154000 79528 157760
rect 84208 154000 84528 157760
rect 89208 154000 89528 157760
rect 94208 154000 94528 157760
rect 99208 154000 99528 157760
rect 104208 154000 104528 157760
rect 109208 154000 109528 157760
rect 114208 154000 114528 157760
rect 119208 154000 119528 157760
rect 124208 154000 124528 157760
rect 129208 154000 129528 157760
rect 134208 154000 134528 157760
rect 139208 154000 139528 157760
rect 144208 154000 144528 157760
rect 149208 154000 149528 157760
rect 154208 154000 154528 157760
rect 159208 154000 159528 157760
rect 164208 154000 164528 157760
rect 169208 154000 169528 157760
rect 174208 154000 174528 157760
rect 179208 154000 179528 157760
rect 184208 154000 184528 157760
rect 189208 154000 189528 157760
rect 194208 154000 194528 157760
rect 199208 154000 199528 157760
rect 204208 154000 204528 157760
rect 209208 154000 209528 157760
rect 214208 154000 214528 157760
rect 219208 154000 219528 157760
rect 224208 154000 224528 157760
rect 229208 154000 229528 157760
rect 234208 154000 234528 157760
rect 239208 154000 239528 157760
rect 244208 154000 244528 157760
rect 249208 154000 249528 157760
rect 254208 154000 254528 157760
rect 259208 154000 259528 157760
rect 264208 154000 264528 157760
rect 269208 154000 269528 157760
rect 274208 154000 274528 157760
rect 279208 154000 279528 157760
rect 284208 154000 284528 157760
rect 289208 154000 289528 157760
rect 294208 154000 294528 157760
rect 299208 154000 299528 157760
rect 304208 154000 304528 157760
rect 309208 154000 309528 157760
rect 314208 154000 314528 157760
rect 319208 154000 319528 157760
rect 324208 154000 324528 157760
rect 329208 154000 329528 157760
rect 334208 154000 334528 157760
rect 339208 154000 339528 157760
rect 344208 154000 344528 157760
rect 349208 154000 349528 157760
rect 354208 154000 354528 157760
rect 359208 154000 359528 157760
rect 364208 154000 364528 157760
rect 369208 154000 369528 157760
rect 374208 154000 374528 157760
rect 379208 154000 379528 157760
rect 384208 154000 384528 157760
rect 389208 154000 389528 157760
rect 394208 154000 394528 157760
rect 399208 154000 399528 157760
rect 404208 154000 404528 157760
rect 409208 154000 409528 157760
rect 414208 154000 414528 157760
rect 419208 154000 419528 157760
rect 424208 154000 424528 157760
rect 429208 154000 429528 157760
rect 434208 154000 434528 157760
rect 439208 154000 439528 157760
rect 444208 154000 444528 157760
rect 449208 154000 449528 157760
rect 454208 154000 454528 157760
rect 459208 154000 459528 157760
rect 464208 154000 464528 157760
rect 469208 154000 469528 157760
rect 474208 154000 474528 157760
rect 479208 154000 479528 157760
rect 484208 154000 484528 157760
rect 489208 154000 489528 157760
rect 494208 154000 494528 157760
rect 499208 154000 499528 157760
rect 504208 154000 504528 157760
rect 509208 154000 509528 157760
rect 514208 154000 514528 157760
rect 519208 154000 519528 157760
rect 524208 2176 524528 157760
rect 529208 2176 529528 157760
rect 534208 2176 534528 157760
rect 539208 2176 539528 157760
rect 544208 2176 544528 157760
rect 549208 2176 549528 157760
rect 554208 2176 554528 157760
rect 559208 2176 559528 157760
rect 564208 2176 564528 157760
rect 569208 2176 569528 157760
rect 574208 2176 574528 157760
<< obsm4 >>
rect 4004 4156 522218 151812
<< metal5 >>
rect 1104 148346 2000 148666
rect 116000 148346 118000 148666
rect 522000 148346 578864 148666
rect 1104 135346 2000 135666
rect 116000 135346 118000 135666
rect 522000 135346 578864 135666
rect 1104 122346 2000 122666
rect 116000 122346 118000 122666
rect 522000 122346 578864 122666
rect 1104 109346 2000 109666
rect 116000 109346 118000 109666
rect 522000 109346 578864 109666
rect 1104 96346 2000 96666
rect 116000 96346 118000 96666
rect 522000 96346 578864 96666
rect 1104 83346 2000 83666
rect 116000 83346 118000 83666
rect 522000 83346 578864 83666
rect 1104 70346 2000 70666
rect 116000 70346 118000 70666
rect 522000 70346 578864 70666
rect 1104 57346 2000 57666
rect 116000 57346 118000 57666
rect 522000 57346 578864 57666
rect 1104 44346 2000 44666
rect 116000 44346 118000 44666
rect 522000 44346 578864 44666
rect 1104 31346 2000 31666
rect 116000 31346 118000 31666
rect 522000 31346 578864 31666
rect 1104 18346 2000 18666
rect 116000 18346 118000 18666
rect 522000 18346 578864 18666
rect 1104 5346 2000 5666
rect 116000 5346 118000 5666
rect 522000 5346 578864 5666
<< obsm5 >>
rect 4004 148986 522260 151812
rect 4004 148026 115680 148986
rect 118320 148026 521680 148986
rect 4004 135986 522260 148026
rect 4004 135026 115680 135986
rect 118320 135026 521680 135986
rect 4004 122986 522260 135026
rect 4004 122026 115680 122986
rect 118320 122026 521680 122986
rect 4004 109986 522260 122026
rect 4004 109026 115680 109986
rect 118320 109026 521680 109986
rect 4004 96986 522260 109026
rect 4004 96026 115680 96986
rect 118320 96026 521680 96986
rect 4004 83986 522260 96026
rect 4004 83026 115680 83986
rect 118320 83026 521680 83986
rect 4004 70986 522260 83026
rect 4004 70026 115680 70986
rect 118320 70026 521680 70986
rect 4004 57986 522260 70026
rect 4004 57026 115680 57986
rect 118320 57026 521680 57986
rect 4004 44986 522260 57026
rect 4004 44026 115680 44986
rect 118320 44026 521680 44986
rect 4004 31986 522260 44026
rect 4004 31026 115680 31986
rect 118320 31026 521680 31986
rect 4004 18986 522260 31026
rect 4004 18026 115680 18986
rect 118320 18026 521680 18986
rect 4004 5986 522260 18026
rect 4004 5026 115680 5986
rect 118320 5026 521680 5986
rect 4004 4156 522260 5026
<< labels >>
rlabel metal5 s 1104 18346 2000 18666 6 VGND
port 1 nsew ground input
rlabel metal5 s 116000 18346 118000 18666 6 VGND
port 1 nsew ground input
rlabel metal5 s 522000 18346 578864 18666 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 44346 2000 44666 6 VGND
port 1 nsew ground input
rlabel metal5 s 116000 44346 118000 44666 6 VGND
port 1 nsew ground input
rlabel metal5 s 522000 44346 578864 44666 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 70346 2000 70666 6 VGND
port 1 nsew ground input
rlabel metal5 s 116000 70346 118000 70666 6 VGND
port 1 nsew ground input
rlabel metal5 s 522000 70346 578864 70666 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 96346 2000 96666 6 VGND
port 1 nsew ground input
rlabel metal5 s 116000 96346 118000 96666 6 VGND
port 1 nsew ground input
rlabel metal5 s 522000 96346 578864 96666 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 122346 2000 122666 6 VGND
port 1 nsew ground input
rlabel metal5 s 116000 122346 118000 122666 6 VGND
port 1 nsew ground input
rlabel metal5 s 522000 122346 578864 122666 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 148346 2000 148666 6 VGND
port 1 nsew ground input
rlabel metal5 s 116000 148346 118000 148666 6 VGND
port 1 nsew ground input
rlabel metal5 s 522000 148346 578864 148666 6 VGND
port 1 nsew ground input
rlabel metal4 s 9208 154000 9528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 19208 154000 19528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 29208 154000 29528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 39208 154000 39528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 49208 154000 49528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 59208 154000 59528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 69208 154000 69528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 79208 154000 79528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 89208 154000 89528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 99208 154000 99528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 109208 154000 109528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 119208 154000 119528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 129208 154000 129528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 139208 154000 139528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 149208 154000 149528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 159208 154000 159528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 169208 154000 169528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 179208 154000 179528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 189208 154000 189528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 199208 154000 199528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 209208 154000 209528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 219208 154000 219528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 229208 154000 229528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 239208 154000 239528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 249208 154000 249528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 259208 154000 259528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 269208 154000 269528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 279208 154000 279528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 289208 154000 289528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 299208 154000 299528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 309208 154000 309528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 319208 154000 319528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 329208 154000 329528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 339208 154000 339528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 349208 154000 349528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 359208 154000 359528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 369208 154000 369528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 379208 154000 379528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 389208 154000 389528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 399208 154000 399528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 409208 154000 409528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 419208 154000 419528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 429208 154000 429528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 439208 154000 439528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 449208 154000 449528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 459208 154000 459528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 469208 154000 469528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 479208 154000 479528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 489208 154000 489528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 499208 154000 499528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 509208 154000 509528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 519208 154000 519528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 529208 2176 529528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 539208 2176 539528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 549208 2176 549528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 559208 2176 559528 157760 6 VGND
port 1 nsew ground input
rlabel metal4 s 569208 2176 569528 157760 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 5346 2000 5666 6 VPWR
port 2 nsew power input
rlabel metal5 s 116000 5346 118000 5666 6 VPWR
port 2 nsew power input
rlabel metal5 s 522000 5346 578864 5666 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 31346 2000 31666 6 VPWR
port 2 nsew power input
rlabel metal5 s 116000 31346 118000 31666 6 VPWR
port 2 nsew power input
rlabel metal5 s 522000 31346 578864 31666 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 57346 2000 57666 6 VPWR
port 2 nsew power input
rlabel metal5 s 116000 57346 118000 57666 6 VPWR
port 2 nsew power input
rlabel metal5 s 522000 57346 578864 57666 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 83346 2000 83666 6 VPWR
port 2 nsew power input
rlabel metal5 s 116000 83346 118000 83666 6 VPWR
port 2 nsew power input
rlabel metal5 s 522000 83346 578864 83666 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 109346 2000 109666 6 VPWR
port 2 nsew power input
rlabel metal5 s 116000 109346 118000 109666 6 VPWR
port 2 nsew power input
rlabel metal5 s 522000 109346 578864 109666 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 135346 2000 135666 6 VPWR
port 2 nsew power input
rlabel metal5 s 116000 135346 118000 135666 6 VPWR
port 2 nsew power input
rlabel metal5 s 522000 135346 578864 135666 6 VPWR
port 2 nsew power input
rlabel metal4 s 4208 154000 4528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 14208 154000 14528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 24208 154000 24528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 34208 154000 34528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 44208 154000 44528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 54208 154000 54528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 64208 154000 64528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 74208 154000 74528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 84208 154000 84528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 94208 154000 94528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 104208 154000 104528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 114208 154000 114528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 124208 154000 124528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 134208 154000 134528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 144208 154000 144528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 154208 154000 154528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 164208 154000 164528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 174208 154000 174528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 184208 154000 184528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 194208 154000 194528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 204208 154000 204528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 214208 154000 214528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 224208 154000 224528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 234208 154000 234528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 244208 154000 244528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 254208 154000 254528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 264208 154000 264528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 274208 154000 274528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 284208 154000 284528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 294208 154000 294528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 304208 154000 304528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 314208 154000 314528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 324208 154000 324528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 334208 154000 334528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 344208 154000 344528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 354208 154000 354528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 364208 154000 364528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 374208 154000 374528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 384208 154000 384528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 394208 154000 394528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 404208 154000 404528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 414208 154000 414528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 424208 154000 424528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 434208 154000 434528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 444208 154000 444528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 454208 154000 454528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 464208 154000 464528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 474208 154000 474528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 484208 154000 484528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 494208 154000 494528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 504208 154000 504528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 514208 154000 514528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 524208 2176 524528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 534208 2176 534528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 544208 2176 544528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 554208 2176 554528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 564208 2176 564528 157760 6 VPWR
port 2 nsew power input
rlabel metal4 s 574208 2176 574528 157760 6 VPWR
port 2 nsew power input
rlabel metal2 s 478 159200 534 160000 6 core_clk
port 3 nsew signal input
rlabel metal2 s 1398 159200 1454 160000 6 core_rstn
port 4 nsew signal input
rlabel metal2 s 508042 0 508098 800 6 debug_in
port 5 nsew signal input
rlabel metal2 s 513378 0 513434 800 6 debug_mode
port 6 nsew signal output
rlabel metal2 s 523958 0 524014 800 6 debug_oeb
port 7 nsew signal output
rlabel metal2 s 518622 0 518678 800 6 debug_out
port 8 nsew signal output
rlabel metal2 s 39762 0 39818 800 6 flash_clk
port 9 nsew signal output
rlabel metal2 s 34518 0 34574 800 6 flash_csb
port 10 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 flash_io0_di
port 11 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 flash_io0_do
port 12 nsew signal output
rlabel metal2 s 55770 0 55826 800 6 flash_io0_oeb
port 13 nsew signal output
rlabel metal2 s 61106 0 61162 800 6 flash_io1_di
port 14 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 flash_io1_do
port 15 nsew signal output
rlabel metal2 s 71686 0 71742 800 6 flash_io1_oeb
port 16 nsew signal output
rlabel metal2 s 77022 0 77078 800 6 flash_io2_di
port 17 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 flash_io2_do
port 18 nsew signal output
rlabel metal3 s 0 6672 800 6792 6 flash_io2_oeb
port 19 nsew signal output
rlabel metal2 s 87694 0 87750 800 6 flash_io3_di
port 20 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 flash_io3_do
port 21 nsew signal output
rlabel metal3 s 0 2184 800 2304 6 flash_io3_oeb
port 22 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 gpio_in_pad
port 23 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 gpio_inenb_pad
port 24 nsew signal output
rlabel metal2 s 13174 0 13230 800 6 gpio_mode0_pad
port 25 nsew signal output
rlabel metal2 s 18510 0 18566 800 6 gpio_mode1_pad
port 26 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 gpio_out_pad
port 27 nsew signal output
rlabel metal2 s 29182 0 29238 800 6 gpio_outenb_pad
port 28 nsew signal output
rlabel metal2 s 103610 0 103666 800 6 hk_ack_i
port 29 nsew signal input
rlabel metal2 s 114282 0 114338 800 6 hk_dat_i[0]
port 30 nsew signal input
rlabel metal2 s 167458 0 167514 800 6 hk_dat_i[10]
port 31 nsew signal input
rlabel metal2 s 172794 0 172850 800 6 hk_dat_i[11]
port 32 nsew signal input
rlabel metal2 s 178130 0 178186 800 6 hk_dat_i[12]
port 33 nsew signal input
rlabel metal2 s 183466 0 183522 800 6 hk_dat_i[13]
port 34 nsew signal input
rlabel metal2 s 188802 0 188858 800 6 hk_dat_i[14]
port 35 nsew signal input
rlabel metal2 s 194138 0 194194 800 6 hk_dat_i[15]
port 36 nsew signal input
rlabel metal2 s 199382 0 199438 800 6 hk_dat_i[16]
port 37 nsew signal input
rlabel metal2 s 204718 0 204774 800 6 hk_dat_i[17]
port 38 nsew signal input
rlabel metal2 s 210054 0 210110 800 6 hk_dat_i[18]
port 39 nsew signal input
rlabel metal2 s 215390 0 215446 800 6 hk_dat_i[19]
port 40 nsew signal input
rlabel metal2 s 119618 0 119674 800 6 hk_dat_i[1]
port 41 nsew signal input
rlabel metal2 s 220726 0 220782 800 6 hk_dat_i[20]
port 42 nsew signal input
rlabel metal2 s 226062 0 226118 800 6 hk_dat_i[21]
port 43 nsew signal input
rlabel metal2 s 231306 0 231362 800 6 hk_dat_i[22]
port 44 nsew signal input
rlabel metal2 s 236642 0 236698 800 6 hk_dat_i[23]
port 45 nsew signal input
rlabel metal2 s 241978 0 242034 800 6 hk_dat_i[24]
port 46 nsew signal input
rlabel metal2 s 247314 0 247370 800 6 hk_dat_i[25]
port 47 nsew signal input
rlabel metal2 s 252650 0 252706 800 6 hk_dat_i[26]
port 48 nsew signal input
rlabel metal2 s 257986 0 258042 800 6 hk_dat_i[27]
port 49 nsew signal input
rlabel metal2 s 263230 0 263286 800 6 hk_dat_i[28]
port 50 nsew signal input
rlabel metal2 s 268566 0 268622 800 6 hk_dat_i[29]
port 51 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 hk_dat_i[2]
port 52 nsew signal input
rlabel metal2 s 273902 0 273958 800 6 hk_dat_i[30]
port 53 nsew signal input
rlabel metal2 s 279238 0 279294 800 6 hk_dat_i[31]
port 54 nsew signal input
rlabel metal2 s 130290 0 130346 800 6 hk_dat_i[3]
port 55 nsew signal input
rlabel metal2 s 135534 0 135590 800 6 hk_dat_i[4]
port 56 nsew signal input
rlabel metal2 s 140870 0 140926 800 6 hk_dat_i[5]
port 57 nsew signal input
rlabel metal2 s 146206 0 146262 800 6 hk_dat_i[6]
port 58 nsew signal input
rlabel metal2 s 151542 0 151598 800 6 hk_dat_i[7]
port 59 nsew signal input
rlabel metal2 s 156878 0 156934 800 6 hk_dat_i[8]
port 60 nsew signal input
rlabel metal2 s 162214 0 162270 800 6 hk_dat_i[9]
port 61 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 hk_stb_o
port 62 nsew signal output
rlabel metal2 s 574558 159200 574614 160000 6 irq[0]
port 63 nsew signal input
rlabel metal2 s 575570 159200 575626 160000 6 irq[1]
port 64 nsew signal input
rlabel metal2 s 576490 159200 576546 160000 6 irq[2]
port 65 nsew signal input
rlabel metal2 s 577502 159200 577558 160000 6 irq[3]
port 66 nsew signal input
rlabel metal2 s 578422 159200 578478 160000 6 irq[4]
port 67 nsew signal input
rlabel metal2 s 579434 159200 579490 160000 6 irq[5]
port 68 nsew signal input
rlabel metal2 s 2410 159200 2466 160000 6 la_iena[0]
port 69 nsew signal output
rlabel metal2 s 392306 159200 392362 160000 6 la_iena[100]
port 70 nsew signal output
rlabel metal2 s 396170 159200 396226 160000 6 la_iena[101]
port 71 nsew signal output
rlabel metal2 s 400034 159200 400090 160000 6 la_iena[102]
port 72 nsew signal output
rlabel metal2 s 403990 159200 404046 160000 6 la_iena[103]
port 73 nsew signal output
rlabel metal2 s 407854 159200 407910 160000 6 la_iena[104]
port 74 nsew signal output
rlabel metal2 s 411810 159200 411866 160000 6 la_iena[105]
port 75 nsew signal output
rlabel metal2 s 415674 159200 415730 160000 6 la_iena[106]
port 76 nsew signal output
rlabel metal2 s 419538 159200 419594 160000 6 la_iena[107]
port 77 nsew signal output
rlabel metal2 s 423494 159200 423550 160000 6 la_iena[108]
port 78 nsew signal output
rlabel metal2 s 427358 159200 427414 160000 6 la_iena[109]
port 79 nsew signal output
rlabel metal2 s 41326 159200 41382 160000 6 la_iena[10]
port 80 nsew signal output
rlabel metal2 s 431222 159200 431278 160000 6 la_iena[110]
port 81 nsew signal output
rlabel metal2 s 435178 159200 435234 160000 6 la_iena[111]
port 82 nsew signal output
rlabel metal2 s 439042 159200 439098 160000 6 la_iena[112]
port 83 nsew signal output
rlabel metal2 s 442998 159200 443054 160000 6 la_iena[113]
port 84 nsew signal output
rlabel metal2 s 446862 159200 446918 160000 6 la_iena[114]
port 85 nsew signal output
rlabel metal2 s 450726 159200 450782 160000 6 la_iena[115]
port 86 nsew signal output
rlabel metal2 s 454682 159200 454738 160000 6 la_iena[116]
port 87 nsew signal output
rlabel metal2 s 458546 159200 458602 160000 6 la_iena[117]
port 88 nsew signal output
rlabel metal2 s 462502 159200 462558 160000 6 la_iena[118]
port 89 nsew signal output
rlabel metal2 s 466366 159200 466422 160000 6 la_iena[119]
port 90 nsew signal output
rlabel metal2 s 45282 159200 45338 160000 6 la_iena[11]
port 91 nsew signal output
rlabel metal2 s 470230 159200 470286 160000 6 la_iena[120]
port 92 nsew signal output
rlabel metal2 s 474186 159200 474242 160000 6 la_iena[121]
port 93 nsew signal output
rlabel metal2 s 478050 159200 478106 160000 6 la_iena[122]
port 94 nsew signal output
rlabel metal2 s 481914 159200 481970 160000 6 la_iena[123]
port 95 nsew signal output
rlabel metal2 s 485870 159200 485926 160000 6 la_iena[124]
port 96 nsew signal output
rlabel metal2 s 489734 159200 489790 160000 6 la_iena[125]
port 97 nsew signal output
rlabel metal2 s 493690 159200 493746 160000 6 la_iena[126]
port 98 nsew signal output
rlabel metal2 s 497554 159200 497610 160000 6 la_iena[127]
port 99 nsew signal output
rlabel metal2 s 49146 159200 49202 160000 6 la_iena[12]
port 100 nsew signal output
rlabel metal2 s 53102 159200 53158 160000 6 la_iena[13]
port 101 nsew signal output
rlabel metal2 s 56966 159200 57022 160000 6 la_iena[14]
port 102 nsew signal output
rlabel metal2 s 60830 159200 60886 160000 6 la_iena[15]
port 103 nsew signal output
rlabel metal2 s 64786 159200 64842 160000 6 la_iena[16]
port 104 nsew signal output
rlabel metal2 s 68650 159200 68706 160000 6 la_iena[17]
port 105 nsew signal output
rlabel metal2 s 72606 159200 72662 160000 6 la_iena[18]
port 106 nsew signal output
rlabel metal2 s 76470 159200 76526 160000 6 la_iena[19]
port 107 nsew signal output
rlabel metal2 s 6274 159200 6330 160000 6 la_iena[1]
port 108 nsew signal output
rlabel metal2 s 80334 159200 80390 160000 6 la_iena[20]
port 109 nsew signal output
rlabel metal2 s 84290 159200 84346 160000 6 la_iena[21]
port 110 nsew signal output
rlabel metal2 s 88154 159200 88210 160000 6 la_iena[22]
port 111 nsew signal output
rlabel metal2 s 92018 159200 92074 160000 6 la_iena[23]
port 112 nsew signal output
rlabel metal2 s 95974 159200 96030 160000 6 la_iena[24]
port 113 nsew signal output
rlabel metal2 s 99838 159200 99894 160000 6 la_iena[25]
port 114 nsew signal output
rlabel metal2 s 103794 159200 103850 160000 6 la_iena[26]
port 115 nsew signal output
rlabel metal2 s 107658 159200 107714 160000 6 la_iena[27]
port 116 nsew signal output
rlabel metal2 s 111522 159200 111578 160000 6 la_iena[28]
port 117 nsew signal output
rlabel metal2 s 115478 159200 115534 160000 6 la_iena[29]
port 118 nsew signal output
rlabel metal2 s 10138 159200 10194 160000 6 la_iena[2]
port 119 nsew signal output
rlabel metal2 s 119342 159200 119398 160000 6 la_iena[30]
port 120 nsew signal output
rlabel metal2 s 123206 159200 123262 160000 6 la_iena[31]
port 121 nsew signal output
rlabel metal2 s 127162 159200 127218 160000 6 la_iena[32]
port 122 nsew signal output
rlabel metal2 s 131026 159200 131082 160000 6 la_iena[33]
port 123 nsew signal output
rlabel metal2 s 134982 159200 135038 160000 6 la_iena[34]
port 124 nsew signal output
rlabel metal2 s 138846 159200 138902 160000 6 la_iena[35]
port 125 nsew signal output
rlabel metal2 s 142710 159200 142766 160000 6 la_iena[36]
port 126 nsew signal output
rlabel metal2 s 146666 159200 146722 160000 6 la_iena[37]
port 127 nsew signal output
rlabel metal2 s 150530 159200 150586 160000 6 la_iena[38]
port 128 nsew signal output
rlabel metal2 s 154486 159200 154542 160000 6 la_iena[39]
port 129 nsew signal output
rlabel metal2 s 14094 159200 14150 160000 6 la_iena[3]
port 130 nsew signal output
rlabel metal2 s 158350 159200 158406 160000 6 la_iena[40]
port 131 nsew signal output
rlabel metal2 s 162214 159200 162270 160000 6 la_iena[41]
port 132 nsew signal output
rlabel metal2 s 166170 159200 166226 160000 6 la_iena[42]
port 133 nsew signal output
rlabel metal2 s 170034 159200 170090 160000 6 la_iena[43]
port 134 nsew signal output
rlabel metal2 s 173898 159200 173954 160000 6 la_iena[44]
port 135 nsew signal output
rlabel metal2 s 177854 159200 177910 160000 6 la_iena[45]
port 136 nsew signal output
rlabel metal2 s 181718 159200 181774 160000 6 la_iena[46]
port 137 nsew signal output
rlabel metal2 s 185674 159200 185730 160000 6 la_iena[47]
port 138 nsew signal output
rlabel metal2 s 189538 159200 189594 160000 6 la_iena[48]
port 139 nsew signal output
rlabel metal2 s 193402 159200 193458 160000 6 la_iena[49]
port 140 nsew signal output
rlabel metal2 s 17958 159200 18014 160000 6 la_iena[4]
port 141 nsew signal output
rlabel metal2 s 197358 159200 197414 160000 6 la_iena[50]
port 142 nsew signal output
rlabel metal2 s 201222 159200 201278 160000 6 la_iena[51]
port 143 nsew signal output
rlabel metal2 s 205086 159200 205142 160000 6 la_iena[52]
port 144 nsew signal output
rlabel metal2 s 209042 159200 209098 160000 6 la_iena[53]
port 145 nsew signal output
rlabel metal2 s 212906 159200 212962 160000 6 la_iena[54]
port 146 nsew signal output
rlabel metal2 s 216862 159200 216918 160000 6 la_iena[55]
port 147 nsew signal output
rlabel metal2 s 220726 159200 220782 160000 6 la_iena[56]
port 148 nsew signal output
rlabel metal2 s 224590 159200 224646 160000 6 la_iena[57]
port 149 nsew signal output
rlabel metal2 s 228546 159200 228602 160000 6 la_iena[58]
port 150 nsew signal output
rlabel metal2 s 232410 159200 232466 160000 6 la_iena[59]
port 151 nsew signal output
rlabel metal2 s 21914 159200 21970 160000 6 la_iena[5]
port 152 nsew signal output
rlabel metal2 s 236274 159200 236330 160000 6 la_iena[60]
port 153 nsew signal output
rlabel metal2 s 240230 159200 240286 160000 6 la_iena[61]
port 154 nsew signal output
rlabel metal2 s 244094 159200 244150 160000 6 la_iena[62]
port 155 nsew signal output
rlabel metal2 s 248050 159200 248106 160000 6 la_iena[63]
port 156 nsew signal output
rlabel metal2 s 251914 159200 251970 160000 6 la_iena[64]
port 157 nsew signal output
rlabel metal2 s 255778 159200 255834 160000 6 la_iena[65]
port 158 nsew signal output
rlabel metal2 s 259734 159200 259790 160000 6 la_iena[66]
port 159 nsew signal output
rlabel metal2 s 263598 159200 263654 160000 6 la_iena[67]
port 160 nsew signal output
rlabel metal2 s 267554 159200 267610 160000 6 la_iena[68]
port 161 nsew signal output
rlabel metal2 s 271418 159200 271474 160000 6 la_iena[69]
port 162 nsew signal output
rlabel metal2 s 25778 159200 25834 160000 6 la_iena[6]
port 163 nsew signal output
rlabel metal2 s 275282 159200 275338 160000 6 la_iena[70]
port 164 nsew signal output
rlabel metal2 s 279238 159200 279294 160000 6 la_iena[71]
port 165 nsew signal output
rlabel metal2 s 283102 159200 283158 160000 6 la_iena[72]
port 166 nsew signal output
rlabel metal2 s 286966 159200 287022 160000 6 la_iena[73]
port 167 nsew signal output
rlabel metal2 s 290922 159200 290978 160000 6 la_iena[74]
port 168 nsew signal output
rlabel metal2 s 294786 159200 294842 160000 6 la_iena[75]
port 169 nsew signal output
rlabel metal2 s 298742 159200 298798 160000 6 la_iena[76]
port 170 nsew signal output
rlabel metal2 s 302606 159200 302662 160000 6 la_iena[77]
port 171 nsew signal output
rlabel metal2 s 306470 159200 306526 160000 6 la_iena[78]
port 172 nsew signal output
rlabel metal2 s 310426 159200 310482 160000 6 la_iena[79]
port 173 nsew signal output
rlabel metal2 s 29642 159200 29698 160000 6 la_iena[7]
port 174 nsew signal output
rlabel metal2 s 314290 159200 314346 160000 6 la_iena[80]
port 175 nsew signal output
rlabel metal2 s 318154 159200 318210 160000 6 la_iena[81]
port 176 nsew signal output
rlabel metal2 s 322110 159200 322166 160000 6 la_iena[82]
port 177 nsew signal output
rlabel metal2 s 325974 159200 326030 160000 6 la_iena[83]
port 178 nsew signal output
rlabel metal2 s 329930 159200 329986 160000 6 la_iena[84]
port 179 nsew signal output
rlabel metal2 s 333794 159200 333850 160000 6 la_iena[85]
port 180 nsew signal output
rlabel metal2 s 337658 159200 337714 160000 6 la_iena[86]
port 181 nsew signal output
rlabel metal2 s 341614 159200 341670 160000 6 la_iena[87]
port 182 nsew signal output
rlabel metal2 s 345478 159200 345534 160000 6 la_iena[88]
port 183 nsew signal output
rlabel metal2 s 349342 159200 349398 160000 6 la_iena[89]
port 184 nsew signal output
rlabel metal2 s 33598 159200 33654 160000 6 la_iena[8]
port 185 nsew signal output
rlabel metal2 s 353298 159200 353354 160000 6 la_iena[90]
port 186 nsew signal output
rlabel metal2 s 357162 159200 357218 160000 6 la_iena[91]
port 187 nsew signal output
rlabel metal2 s 361118 159200 361174 160000 6 la_iena[92]
port 188 nsew signal output
rlabel metal2 s 364982 159200 365038 160000 6 la_iena[93]
port 189 nsew signal output
rlabel metal2 s 368846 159200 368902 160000 6 la_iena[94]
port 190 nsew signal output
rlabel metal2 s 372802 159200 372858 160000 6 la_iena[95]
port 191 nsew signal output
rlabel metal2 s 376666 159200 376722 160000 6 la_iena[96]
port 192 nsew signal output
rlabel metal2 s 380622 159200 380678 160000 6 la_iena[97]
port 193 nsew signal output
rlabel metal2 s 384486 159200 384542 160000 6 la_iena[98]
port 194 nsew signal output
rlabel metal2 s 388350 159200 388406 160000 6 la_iena[99]
port 195 nsew signal output
rlabel metal2 s 37462 159200 37518 160000 6 la_iena[9]
port 196 nsew signal output
rlabel metal2 s 3330 159200 3386 160000 6 la_input[0]
port 197 nsew signal input
rlabel metal2 s 393226 159200 393282 160000 6 la_input[100]
port 198 nsew signal input
rlabel metal2 s 397182 159200 397238 160000 6 la_input[101]
port 199 nsew signal input
rlabel metal2 s 401046 159200 401102 160000 6 la_input[102]
port 200 nsew signal input
rlabel metal2 s 404910 159200 404966 160000 6 la_input[103]
port 201 nsew signal input
rlabel metal2 s 408866 159200 408922 160000 6 la_input[104]
port 202 nsew signal input
rlabel metal2 s 412730 159200 412786 160000 6 la_input[105]
port 203 nsew signal input
rlabel metal2 s 416686 159200 416742 160000 6 la_input[106]
port 204 nsew signal input
rlabel metal2 s 420550 159200 420606 160000 6 la_input[107]
port 205 nsew signal input
rlabel metal2 s 424414 159200 424470 160000 6 la_input[108]
port 206 nsew signal input
rlabel metal2 s 428370 159200 428426 160000 6 la_input[109]
port 207 nsew signal input
rlabel metal2 s 42338 159200 42394 160000 6 la_input[10]
port 208 nsew signal input
rlabel metal2 s 432234 159200 432290 160000 6 la_input[110]
port 209 nsew signal input
rlabel metal2 s 436098 159200 436154 160000 6 la_input[111]
port 210 nsew signal input
rlabel metal2 s 440054 159200 440110 160000 6 la_input[112]
port 211 nsew signal input
rlabel metal2 s 443918 159200 443974 160000 6 la_input[113]
port 212 nsew signal input
rlabel metal2 s 447874 159200 447930 160000 6 la_input[114]
port 213 nsew signal input
rlabel metal2 s 451738 159200 451794 160000 6 la_input[115]
port 214 nsew signal input
rlabel metal2 s 455602 159200 455658 160000 6 la_input[116]
port 215 nsew signal input
rlabel metal2 s 459558 159200 459614 160000 6 la_input[117]
port 216 nsew signal input
rlabel metal2 s 463422 159200 463478 160000 6 la_input[118]
port 217 nsew signal input
rlabel metal2 s 467286 159200 467342 160000 6 la_input[119]
port 218 nsew signal input
rlabel metal2 s 46202 159200 46258 160000 6 la_input[11]
port 219 nsew signal input
rlabel metal2 s 471242 159200 471298 160000 6 la_input[120]
port 220 nsew signal input
rlabel metal2 s 475106 159200 475162 160000 6 la_input[121]
port 221 nsew signal input
rlabel metal2 s 479062 159200 479118 160000 6 la_input[122]
port 222 nsew signal input
rlabel metal2 s 482926 159200 482982 160000 6 la_input[123]
port 223 nsew signal input
rlabel metal2 s 486790 159200 486846 160000 6 la_input[124]
port 224 nsew signal input
rlabel metal2 s 490746 159200 490802 160000 6 la_input[125]
port 225 nsew signal input
rlabel metal2 s 494610 159200 494666 160000 6 la_input[126]
port 226 nsew signal input
rlabel metal2 s 498566 159200 498622 160000 6 la_input[127]
port 227 nsew signal input
rlabel metal2 s 50158 159200 50214 160000 6 la_input[12]
port 228 nsew signal input
rlabel metal2 s 54022 159200 54078 160000 6 la_input[13]
port 229 nsew signal input
rlabel metal2 s 57978 159200 58034 160000 6 la_input[14]
port 230 nsew signal input
rlabel metal2 s 61842 159200 61898 160000 6 la_input[15]
port 231 nsew signal input
rlabel metal2 s 65706 159200 65762 160000 6 la_input[16]
port 232 nsew signal input
rlabel metal2 s 69662 159200 69718 160000 6 la_input[17]
port 233 nsew signal input
rlabel metal2 s 73526 159200 73582 160000 6 la_input[18]
port 234 nsew signal input
rlabel metal2 s 77482 159200 77538 160000 6 la_input[19]
port 235 nsew signal input
rlabel metal2 s 7286 159200 7342 160000 6 la_input[1]
port 236 nsew signal input
rlabel metal2 s 81346 159200 81402 160000 6 la_input[20]
port 237 nsew signal input
rlabel metal2 s 85210 159200 85266 160000 6 la_input[21]
port 238 nsew signal input
rlabel metal2 s 89166 159200 89222 160000 6 la_input[22]
port 239 nsew signal input
rlabel metal2 s 93030 159200 93086 160000 6 la_input[23]
port 240 nsew signal input
rlabel metal2 s 96894 159200 96950 160000 6 la_input[24]
port 241 nsew signal input
rlabel metal2 s 100850 159200 100906 160000 6 la_input[25]
port 242 nsew signal input
rlabel metal2 s 104714 159200 104770 160000 6 la_input[26]
port 243 nsew signal input
rlabel metal2 s 108670 159200 108726 160000 6 la_input[27]
port 244 nsew signal input
rlabel metal2 s 112534 159200 112590 160000 6 la_input[28]
port 245 nsew signal input
rlabel metal2 s 116398 159200 116454 160000 6 la_input[29]
port 246 nsew signal input
rlabel metal2 s 11150 159200 11206 160000 6 la_input[2]
port 247 nsew signal input
rlabel metal2 s 120354 159200 120410 160000 6 la_input[30]
port 248 nsew signal input
rlabel metal2 s 124218 159200 124274 160000 6 la_input[31]
port 249 nsew signal input
rlabel metal2 s 128082 159200 128138 160000 6 la_input[32]
port 250 nsew signal input
rlabel metal2 s 132038 159200 132094 160000 6 la_input[33]
port 251 nsew signal input
rlabel metal2 s 135902 159200 135958 160000 6 la_input[34]
port 252 nsew signal input
rlabel metal2 s 139858 159200 139914 160000 6 la_input[35]
port 253 nsew signal input
rlabel metal2 s 143722 159200 143778 160000 6 la_input[36]
port 254 nsew signal input
rlabel metal2 s 147586 159200 147642 160000 6 la_input[37]
port 255 nsew signal input
rlabel metal2 s 151542 159200 151598 160000 6 la_input[38]
port 256 nsew signal input
rlabel metal2 s 155406 159200 155462 160000 6 la_input[39]
port 257 nsew signal input
rlabel metal2 s 15014 159200 15070 160000 6 la_input[3]
port 258 nsew signal input
rlabel metal2 s 159270 159200 159326 160000 6 la_input[40]
port 259 nsew signal input
rlabel metal2 s 163226 159200 163282 160000 6 la_input[41]
port 260 nsew signal input
rlabel metal2 s 167090 159200 167146 160000 6 la_input[42]
port 261 nsew signal input
rlabel metal2 s 171046 159200 171102 160000 6 la_input[43]
port 262 nsew signal input
rlabel metal2 s 174910 159200 174966 160000 6 la_input[44]
port 263 nsew signal input
rlabel metal2 s 178774 159200 178830 160000 6 la_input[45]
port 264 nsew signal input
rlabel metal2 s 182730 159200 182786 160000 6 la_input[46]
port 265 nsew signal input
rlabel metal2 s 186594 159200 186650 160000 6 la_input[47]
port 266 nsew signal input
rlabel metal2 s 190550 159200 190606 160000 6 la_input[48]
port 267 nsew signal input
rlabel metal2 s 194414 159200 194470 160000 6 la_input[49]
port 268 nsew signal input
rlabel metal2 s 18970 159200 19026 160000 6 la_input[4]
port 269 nsew signal input
rlabel metal2 s 198278 159200 198334 160000 6 la_input[50]
port 270 nsew signal input
rlabel metal2 s 202234 159200 202290 160000 6 la_input[51]
port 271 nsew signal input
rlabel metal2 s 206098 159200 206154 160000 6 la_input[52]
port 272 nsew signal input
rlabel metal2 s 209962 159200 210018 160000 6 la_input[53]
port 273 nsew signal input
rlabel metal2 s 213918 159200 213974 160000 6 la_input[54]
port 274 nsew signal input
rlabel metal2 s 217782 159200 217838 160000 6 la_input[55]
port 275 nsew signal input
rlabel metal2 s 221738 159200 221794 160000 6 la_input[56]
port 276 nsew signal input
rlabel metal2 s 225602 159200 225658 160000 6 la_input[57]
port 277 nsew signal input
rlabel metal2 s 229466 159200 229522 160000 6 la_input[58]
port 278 nsew signal input
rlabel metal2 s 233422 159200 233478 160000 6 la_input[59]
port 279 nsew signal input
rlabel metal2 s 22834 159200 22890 160000 6 la_input[5]
port 280 nsew signal input
rlabel metal2 s 237286 159200 237342 160000 6 la_input[60]
port 281 nsew signal input
rlabel metal2 s 241150 159200 241206 160000 6 la_input[61]
port 282 nsew signal input
rlabel metal2 s 245106 159200 245162 160000 6 la_input[62]
port 283 nsew signal input
rlabel metal2 s 248970 159200 249026 160000 6 la_input[63]
port 284 nsew signal input
rlabel metal2 s 252926 159200 252982 160000 6 la_input[64]
port 285 nsew signal input
rlabel metal2 s 256790 159200 256846 160000 6 la_input[65]
port 286 nsew signal input
rlabel metal2 s 260654 159200 260710 160000 6 la_input[66]
port 287 nsew signal input
rlabel metal2 s 264610 159200 264666 160000 6 la_input[67]
port 288 nsew signal input
rlabel metal2 s 268474 159200 268530 160000 6 la_input[68]
port 289 nsew signal input
rlabel metal2 s 272338 159200 272394 160000 6 la_input[69]
port 290 nsew signal input
rlabel metal2 s 26790 159200 26846 160000 6 la_input[6]
port 291 nsew signal input
rlabel metal2 s 276294 159200 276350 160000 6 la_input[70]
port 292 nsew signal input
rlabel metal2 s 280158 159200 280214 160000 6 la_input[71]
port 293 nsew signal input
rlabel metal2 s 284114 159200 284170 160000 6 la_input[72]
port 294 nsew signal input
rlabel metal2 s 287978 159200 288034 160000 6 la_input[73]
port 295 nsew signal input
rlabel metal2 s 291842 159200 291898 160000 6 la_input[74]
port 296 nsew signal input
rlabel metal2 s 295798 159200 295854 160000 6 la_input[75]
port 297 nsew signal input
rlabel metal2 s 299662 159200 299718 160000 6 la_input[76]
port 298 nsew signal input
rlabel metal2 s 303618 159200 303674 160000 6 la_input[77]
port 299 nsew signal input
rlabel metal2 s 307482 159200 307538 160000 6 la_input[78]
port 300 nsew signal input
rlabel metal2 s 311346 159200 311402 160000 6 la_input[79]
port 301 nsew signal input
rlabel metal2 s 30654 159200 30710 160000 6 la_input[7]
port 302 nsew signal input
rlabel metal2 s 315302 159200 315358 160000 6 la_input[80]
port 303 nsew signal input
rlabel metal2 s 319166 159200 319222 160000 6 la_input[81]
port 304 nsew signal input
rlabel metal2 s 323030 159200 323086 160000 6 la_input[82]
port 305 nsew signal input
rlabel metal2 s 326986 159200 327042 160000 6 la_input[83]
port 306 nsew signal input
rlabel metal2 s 330850 159200 330906 160000 6 la_input[84]
port 307 nsew signal input
rlabel metal2 s 334806 159200 334862 160000 6 la_input[85]
port 308 nsew signal input
rlabel metal2 s 338670 159200 338726 160000 6 la_input[86]
port 309 nsew signal input
rlabel metal2 s 342534 159200 342590 160000 6 la_input[87]
port 310 nsew signal input
rlabel metal2 s 346490 159200 346546 160000 6 la_input[88]
port 311 nsew signal input
rlabel metal2 s 350354 159200 350410 160000 6 la_input[89]
port 312 nsew signal input
rlabel metal2 s 34518 159200 34574 160000 6 la_input[8]
port 313 nsew signal input
rlabel metal2 s 354218 159200 354274 160000 6 la_input[90]
port 314 nsew signal input
rlabel metal2 s 358174 159200 358230 160000 6 la_input[91]
port 315 nsew signal input
rlabel metal2 s 362038 159200 362094 160000 6 la_input[92]
port 316 nsew signal input
rlabel metal2 s 365994 159200 366050 160000 6 la_input[93]
port 317 nsew signal input
rlabel metal2 s 369858 159200 369914 160000 6 la_input[94]
port 318 nsew signal input
rlabel metal2 s 373722 159200 373778 160000 6 la_input[95]
port 319 nsew signal input
rlabel metal2 s 377678 159200 377734 160000 6 la_input[96]
port 320 nsew signal input
rlabel metal2 s 381542 159200 381598 160000 6 la_input[97]
port 321 nsew signal input
rlabel metal2 s 385498 159200 385554 160000 6 la_input[98]
port 322 nsew signal input
rlabel metal2 s 389362 159200 389418 160000 6 la_input[99]
port 323 nsew signal input
rlabel metal2 s 38474 159200 38530 160000 6 la_input[9]
port 324 nsew signal input
rlabel metal2 s 4342 159200 4398 160000 6 la_oenb[0]
port 325 nsew signal output
rlabel metal2 s 394238 159200 394294 160000 6 la_oenb[100]
port 326 nsew signal output
rlabel metal2 s 398102 159200 398158 160000 6 la_oenb[101]
port 327 nsew signal output
rlabel metal2 s 402058 159200 402114 160000 6 la_oenb[102]
port 328 nsew signal output
rlabel metal2 s 405922 159200 405978 160000 6 la_oenb[103]
port 329 nsew signal output
rlabel metal2 s 409786 159200 409842 160000 6 la_oenb[104]
port 330 nsew signal output
rlabel metal2 s 413742 159200 413798 160000 6 la_oenb[105]
port 331 nsew signal output
rlabel metal2 s 417606 159200 417662 160000 6 la_oenb[106]
port 332 nsew signal output
rlabel metal2 s 421562 159200 421618 160000 6 la_oenb[107]
port 333 nsew signal output
rlabel metal2 s 425426 159200 425482 160000 6 la_oenb[108]
port 334 nsew signal output
rlabel metal2 s 429290 159200 429346 160000 6 la_oenb[109]
port 335 nsew signal output
rlabel metal2 s 43350 159200 43406 160000 6 la_oenb[10]
port 336 nsew signal output
rlabel metal2 s 433246 159200 433302 160000 6 la_oenb[110]
port 337 nsew signal output
rlabel metal2 s 437110 159200 437166 160000 6 la_oenb[111]
port 338 nsew signal output
rlabel metal2 s 440974 159200 441030 160000 6 la_oenb[112]
port 339 nsew signal output
rlabel metal2 s 444930 159200 444986 160000 6 la_oenb[113]
port 340 nsew signal output
rlabel metal2 s 448794 159200 448850 160000 6 la_oenb[114]
port 341 nsew signal output
rlabel metal2 s 452750 159200 452806 160000 6 la_oenb[115]
port 342 nsew signal output
rlabel metal2 s 456614 159200 456670 160000 6 la_oenb[116]
port 343 nsew signal output
rlabel metal2 s 460478 159200 460534 160000 6 la_oenb[117]
port 344 nsew signal output
rlabel metal2 s 464434 159200 464490 160000 6 la_oenb[118]
port 345 nsew signal output
rlabel metal2 s 468298 159200 468354 160000 6 la_oenb[119]
port 346 nsew signal output
rlabel metal2 s 47214 159200 47270 160000 6 la_oenb[11]
port 347 nsew signal output
rlabel metal2 s 472162 159200 472218 160000 6 la_oenb[120]
port 348 nsew signal output
rlabel metal2 s 476118 159200 476174 160000 6 la_oenb[121]
port 349 nsew signal output
rlabel metal2 s 479982 159200 480038 160000 6 la_oenb[122]
port 350 nsew signal output
rlabel metal2 s 483938 159200 483994 160000 6 la_oenb[123]
port 351 nsew signal output
rlabel metal2 s 487802 159200 487858 160000 6 la_oenb[124]
port 352 nsew signal output
rlabel metal2 s 491666 159200 491722 160000 6 la_oenb[125]
port 353 nsew signal output
rlabel metal2 s 495622 159200 495678 160000 6 la_oenb[126]
port 354 nsew signal output
rlabel metal2 s 499486 159200 499542 160000 6 la_oenb[127]
port 355 nsew signal output
rlabel metal2 s 51078 159200 51134 160000 6 la_oenb[12]
port 356 nsew signal output
rlabel metal2 s 55034 159200 55090 160000 6 la_oenb[13]
port 357 nsew signal output
rlabel metal2 s 58898 159200 58954 160000 6 la_oenb[14]
port 358 nsew signal output
rlabel metal2 s 62854 159200 62910 160000 6 la_oenb[15]
port 359 nsew signal output
rlabel metal2 s 66718 159200 66774 160000 6 la_oenb[16]
port 360 nsew signal output
rlabel metal2 s 70582 159200 70638 160000 6 la_oenb[17]
port 361 nsew signal output
rlabel metal2 s 74538 159200 74594 160000 6 la_oenb[18]
port 362 nsew signal output
rlabel metal2 s 78402 159200 78458 160000 6 la_oenb[19]
port 363 nsew signal output
rlabel metal2 s 8206 159200 8262 160000 6 la_oenb[1]
port 364 nsew signal output
rlabel metal2 s 82266 159200 82322 160000 6 la_oenb[20]
port 365 nsew signal output
rlabel metal2 s 86222 159200 86278 160000 6 la_oenb[21]
port 366 nsew signal output
rlabel metal2 s 90086 159200 90142 160000 6 la_oenb[22]
port 367 nsew signal output
rlabel metal2 s 94042 159200 94098 160000 6 la_oenb[23]
port 368 nsew signal output
rlabel metal2 s 97906 159200 97962 160000 6 la_oenb[24]
port 369 nsew signal output
rlabel metal2 s 101770 159200 101826 160000 6 la_oenb[25]
port 370 nsew signal output
rlabel metal2 s 105726 159200 105782 160000 6 la_oenb[26]
port 371 nsew signal output
rlabel metal2 s 109590 159200 109646 160000 6 la_oenb[27]
port 372 nsew signal output
rlabel metal2 s 113546 159200 113602 160000 6 la_oenb[28]
port 373 nsew signal output
rlabel metal2 s 117410 159200 117466 160000 6 la_oenb[29]
port 374 nsew signal output
rlabel metal2 s 12162 159200 12218 160000 6 la_oenb[2]
port 375 nsew signal output
rlabel metal2 s 121274 159200 121330 160000 6 la_oenb[30]
port 376 nsew signal output
rlabel metal2 s 125230 159200 125286 160000 6 la_oenb[31]
port 377 nsew signal output
rlabel metal2 s 129094 159200 129150 160000 6 la_oenb[32]
port 378 nsew signal output
rlabel metal2 s 132958 159200 133014 160000 6 la_oenb[33]
port 379 nsew signal output
rlabel metal2 s 136914 159200 136970 160000 6 la_oenb[34]
port 380 nsew signal output
rlabel metal2 s 140778 159200 140834 160000 6 la_oenb[35]
port 381 nsew signal output
rlabel metal2 s 144734 159200 144790 160000 6 la_oenb[36]
port 382 nsew signal output
rlabel metal2 s 148598 159200 148654 160000 6 la_oenb[37]
port 383 nsew signal output
rlabel metal2 s 152462 159200 152518 160000 6 la_oenb[38]
port 384 nsew signal output
rlabel metal2 s 156418 159200 156474 160000 6 la_oenb[39]
port 385 nsew signal output
rlabel metal2 s 16026 159200 16082 160000 6 la_oenb[3]
port 386 nsew signal output
rlabel metal2 s 160282 159200 160338 160000 6 la_oenb[40]
port 387 nsew signal output
rlabel metal2 s 164146 159200 164202 160000 6 la_oenb[41]
port 388 nsew signal output
rlabel metal2 s 168102 159200 168158 160000 6 la_oenb[42]
port 389 nsew signal output
rlabel metal2 s 171966 159200 172022 160000 6 la_oenb[43]
port 390 nsew signal output
rlabel metal2 s 175922 159200 175978 160000 6 la_oenb[44]
port 391 nsew signal output
rlabel metal2 s 179786 159200 179842 160000 6 la_oenb[45]
port 392 nsew signal output
rlabel metal2 s 183650 159200 183706 160000 6 la_oenb[46]
port 393 nsew signal output
rlabel metal2 s 187606 159200 187662 160000 6 la_oenb[47]
port 394 nsew signal output
rlabel metal2 s 191470 159200 191526 160000 6 la_oenb[48]
port 395 nsew signal output
rlabel metal2 s 195334 159200 195390 160000 6 la_oenb[49]
port 396 nsew signal output
rlabel metal2 s 19890 159200 19946 160000 6 la_oenb[4]
port 397 nsew signal output
rlabel metal2 s 199290 159200 199346 160000 6 la_oenb[50]
port 398 nsew signal output
rlabel metal2 s 203154 159200 203210 160000 6 la_oenb[51]
port 399 nsew signal output
rlabel metal2 s 207110 159200 207166 160000 6 la_oenb[52]
port 400 nsew signal output
rlabel metal2 s 210974 159200 211030 160000 6 la_oenb[53]
port 401 nsew signal output
rlabel metal2 s 214838 159200 214894 160000 6 la_oenb[54]
port 402 nsew signal output
rlabel metal2 s 218794 159200 218850 160000 6 la_oenb[55]
port 403 nsew signal output
rlabel metal2 s 222658 159200 222714 160000 6 la_oenb[56]
port 404 nsew signal output
rlabel metal2 s 226614 159200 226670 160000 6 la_oenb[57]
port 405 nsew signal output
rlabel metal2 s 230478 159200 230534 160000 6 la_oenb[58]
port 406 nsew signal output
rlabel metal2 s 234342 159200 234398 160000 6 la_oenb[59]
port 407 nsew signal output
rlabel metal2 s 23846 159200 23902 160000 6 la_oenb[5]
port 408 nsew signal output
rlabel metal2 s 238298 159200 238354 160000 6 la_oenb[60]
port 409 nsew signal output
rlabel metal2 s 242162 159200 242218 160000 6 la_oenb[61]
port 410 nsew signal output
rlabel metal2 s 246026 159200 246082 160000 6 la_oenb[62]
port 411 nsew signal output
rlabel metal2 s 249982 159200 250038 160000 6 la_oenb[63]
port 412 nsew signal output
rlabel metal2 s 253846 159200 253902 160000 6 la_oenb[64]
port 413 nsew signal output
rlabel metal2 s 257802 159200 257858 160000 6 la_oenb[65]
port 414 nsew signal output
rlabel metal2 s 261666 159200 261722 160000 6 la_oenb[66]
port 415 nsew signal output
rlabel metal2 s 265530 159200 265586 160000 6 la_oenb[67]
port 416 nsew signal output
rlabel metal2 s 269486 159200 269542 160000 6 la_oenb[68]
port 417 nsew signal output
rlabel metal2 s 273350 159200 273406 160000 6 la_oenb[69]
port 418 nsew signal output
rlabel metal2 s 27710 159200 27766 160000 6 la_oenb[6]
port 419 nsew signal output
rlabel metal2 s 277214 159200 277270 160000 6 la_oenb[70]
port 420 nsew signal output
rlabel metal2 s 281170 159200 281226 160000 6 la_oenb[71]
port 421 nsew signal output
rlabel metal2 s 285034 159200 285090 160000 6 la_oenb[72]
port 422 nsew signal output
rlabel metal2 s 288990 159200 289046 160000 6 la_oenb[73]
port 423 nsew signal output
rlabel metal2 s 292854 159200 292910 160000 6 la_oenb[74]
port 424 nsew signal output
rlabel metal2 s 296718 159200 296774 160000 6 la_oenb[75]
port 425 nsew signal output
rlabel metal2 s 300674 159200 300730 160000 6 la_oenb[76]
port 426 nsew signal output
rlabel metal2 s 304538 159200 304594 160000 6 la_oenb[77]
port 427 nsew signal output
rlabel metal2 s 308494 159200 308550 160000 6 la_oenb[78]
port 428 nsew signal output
rlabel metal2 s 312358 159200 312414 160000 6 la_oenb[79]
port 429 nsew signal output
rlabel metal2 s 31666 159200 31722 160000 6 la_oenb[7]
port 430 nsew signal output
rlabel metal2 s 316222 159200 316278 160000 6 la_oenb[80]
port 431 nsew signal output
rlabel metal2 s 320178 159200 320234 160000 6 la_oenb[81]
port 432 nsew signal output
rlabel metal2 s 324042 159200 324098 160000 6 la_oenb[82]
port 433 nsew signal output
rlabel metal2 s 327906 159200 327962 160000 6 la_oenb[83]
port 434 nsew signal output
rlabel metal2 s 331862 159200 331918 160000 6 la_oenb[84]
port 435 nsew signal output
rlabel metal2 s 335726 159200 335782 160000 6 la_oenb[85]
port 436 nsew signal output
rlabel metal2 s 339682 159200 339738 160000 6 la_oenb[86]
port 437 nsew signal output
rlabel metal2 s 343546 159200 343602 160000 6 la_oenb[87]
port 438 nsew signal output
rlabel metal2 s 347410 159200 347466 160000 6 la_oenb[88]
port 439 nsew signal output
rlabel metal2 s 351366 159200 351422 160000 6 la_oenb[89]
port 440 nsew signal output
rlabel metal2 s 35530 159200 35586 160000 6 la_oenb[8]
port 441 nsew signal output
rlabel metal2 s 355230 159200 355286 160000 6 la_oenb[90]
port 442 nsew signal output
rlabel metal2 s 359094 159200 359150 160000 6 la_oenb[91]
port 443 nsew signal output
rlabel metal2 s 363050 159200 363106 160000 6 la_oenb[92]
port 444 nsew signal output
rlabel metal2 s 366914 159200 366970 160000 6 la_oenb[93]
port 445 nsew signal output
rlabel metal2 s 370870 159200 370926 160000 6 la_oenb[94]
port 446 nsew signal output
rlabel metal2 s 374734 159200 374790 160000 6 la_oenb[95]
port 447 nsew signal output
rlabel metal2 s 378598 159200 378654 160000 6 la_oenb[96]
port 448 nsew signal output
rlabel metal2 s 382554 159200 382610 160000 6 la_oenb[97]
port 449 nsew signal output
rlabel metal2 s 386418 159200 386474 160000 6 la_oenb[98]
port 450 nsew signal output
rlabel metal2 s 390282 159200 390338 160000 6 la_oenb[99]
port 451 nsew signal output
rlabel metal2 s 39394 159200 39450 160000 6 la_oenb[9]
port 452 nsew signal output
rlabel metal2 s 5262 159200 5318 160000 6 la_output[0]
port 453 nsew signal output
rlabel metal2 s 395158 159200 395214 160000 6 la_output[100]
port 454 nsew signal output
rlabel metal2 s 399114 159200 399170 160000 6 la_output[101]
port 455 nsew signal output
rlabel metal2 s 402978 159200 403034 160000 6 la_output[102]
port 456 nsew signal output
rlabel metal2 s 406934 159200 406990 160000 6 la_output[103]
port 457 nsew signal output
rlabel metal2 s 410798 159200 410854 160000 6 la_output[104]
port 458 nsew signal output
rlabel metal2 s 414662 159200 414718 160000 6 la_output[105]
port 459 nsew signal output
rlabel metal2 s 418618 159200 418674 160000 6 la_output[106]
port 460 nsew signal output
rlabel metal2 s 422482 159200 422538 160000 6 la_output[107]
port 461 nsew signal output
rlabel metal2 s 426346 159200 426402 160000 6 la_output[108]
port 462 nsew signal output
rlabel metal2 s 430302 159200 430358 160000 6 la_output[109]
port 463 nsew signal output
rlabel metal2 s 44270 159200 44326 160000 6 la_output[10]
port 464 nsew signal output
rlabel metal2 s 434166 159200 434222 160000 6 la_output[110]
port 465 nsew signal output
rlabel metal2 s 438122 159200 438178 160000 6 la_output[111]
port 466 nsew signal output
rlabel metal2 s 441986 159200 442042 160000 6 la_output[112]
port 467 nsew signal output
rlabel metal2 s 445850 159200 445906 160000 6 la_output[113]
port 468 nsew signal output
rlabel metal2 s 449806 159200 449862 160000 6 la_output[114]
port 469 nsew signal output
rlabel metal2 s 453670 159200 453726 160000 6 la_output[115]
port 470 nsew signal output
rlabel metal2 s 457626 159200 457682 160000 6 la_output[116]
port 471 nsew signal output
rlabel metal2 s 461490 159200 461546 160000 6 la_output[117]
port 472 nsew signal output
rlabel metal2 s 465354 159200 465410 160000 6 la_output[118]
port 473 nsew signal output
rlabel metal2 s 469310 159200 469366 160000 6 la_output[119]
port 474 nsew signal output
rlabel metal2 s 48226 159200 48282 160000 6 la_output[11]
port 475 nsew signal output
rlabel metal2 s 473174 159200 473230 160000 6 la_output[120]
port 476 nsew signal output
rlabel metal2 s 477038 159200 477094 160000 6 la_output[121]
port 477 nsew signal output
rlabel metal2 s 480994 159200 481050 160000 6 la_output[122]
port 478 nsew signal output
rlabel metal2 s 484858 159200 484914 160000 6 la_output[123]
port 479 nsew signal output
rlabel metal2 s 488814 159200 488870 160000 6 la_output[124]
port 480 nsew signal output
rlabel metal2 s 492678 159200 492734 160000 6 la_output[125]
port 481 nsew signal output
rlabel metal2 s 496542 159200 496598 160000 6 la_output[126]
port 482 nsew signal output
rlabel metal2 s 500498 159200 500554 160000 6 la_output[127]
port 483 nsew signal output
rlabel metal2 s 52090 159200 52146 160000 6 la_output[12]
port 484 nsew signal output
rlabel metal2 s 55954 159200 56010 160000 6 la_output[13]
port 485 nsew signal output
rlabel metal2 s 59910 159200 59966 160000 6 la_output[14]
port 486 nsew signal output
rlabel metal2 s 63774 159200 63830 160000 6 la_output[15]
port 487 nsew signal output
rlabel metal2 s 67730 159200 67786 160000 6 la_output[16]
port 488 nsew signal output
rlabel metal2 s 71594 159200 71650 160000 6 la_output[17]
port 489 nsew signal output
rlabel metal2 s 75458 159200 75514 160000 6 la_output[18]
port 490 nsew signal output
rlabel metal2 s 79414 159200 79470 160000 6 la_output[19]
port 491 nsew signal output
rlabel metal2 s 9218 159200 9274 160000 6 la_output[1]
port 492 nsew signal output
rlabel metal2 s 83278 159200 83334 160000 6 la_output[20]
port 493 nsew signal output
rlabel metal2 s 87142 159200 87198 160000 6 la_output[21]
port 494 nsew signal output
rlabel metal2 s 91098 159200 91154 160000 6 la_output[22]
port 495 nsew signal output
rlabel metal2 s 94962 159200 95018 160000 6 la_output[23]
port 496 nsew signal output
rlabel metal2 s 98918 159200 98974 160000 6 la_output[24]
port 497 nsew signal output
rlabel metal2 s 102782 159200 102838 160000 6 la_output[25]
port 498 nsew signal output
rlabel metal2 s 106646 159200 106702 160000 6 la_output[26]
port 499 nsew signal output
rlabel metal2 s 110602 159200 110658 160000 6 la_output[27]
port 500 nsew signal output
rlabel metal2 s 114466 159200 114522 160000 6 la_output[28]
port 501 nsew signal output
rlabel metal2 s 118330 159200 118386 160000 6 la_output[29]
port 502 nsew signal output
rlabel metal2 s 13082 159200 13138 160000 6 la_output[2]
port 503 nsew signal output
rlabel metal2 s 122286 159200 122342 160000 6 la_output[30]
port 504 nsew signal output
rlabel metal2 s 126150 159200 126206 160000 6 la_output[31]
port 505 nsew signal output
rlabel metal2 s 130106 159200 130162 160000 6 la_output[32]
port 506 nsew signal output
rlabel metal2 s 133970 159200 134026 160000 6 la_output[33]
port 507 nsew signal output
rlabel metal2 s 137834 159200 137890 160000 6 la_output[34]
port 508 nsew signal output
rlabel metal2 s 141790 159200 141846 160000 6 la_output[35]
port 509 nsew signal output
rlabel metal2 s 145654 159200 145710 160000 6 la_output[36]
port 510 nsew signal output
rlabel metal2 s 149610 159200 149666 160000 6 la_output[37]
port 511 nsew signal output
rlabel metal2 s 153474 159200 153530 160000 6 la_output[38]
port 512 nsew signal output
rlabel metal2 s 157338 159200 157394 160000 6 la_output[39]
port 513 nsew signal output
rlabel metal2 s 17038 159200 17094 160000 6 la_output[3]
port 514 nsew signal output
rlabel metal2 s 161294 159200 161350 160000 6 la_output[40]
port 515 nsew signal output
rlabel metal2 s 165158 159200 165214 160000 6 la_output[41]
port 516 nsew signal output
rlabel metal2 s 169022 159200 169078 160000 6 la_output[42]
port 517 nsew signal output
rlabel metal2 s 172978 159200 173034 160000 6 la_output[43]
port 518 nsew signal output
rlabel metal2 s 176842 159200 176898 160000 6 la_output[44]
port 519 nsew signal output
rlabel metal2 s 180798 159200 180854 160000 6 la_output[45]
port 520 nsew signal output
rlabel metal2 s 184662 159200 184718 160000 6 la_output[46]
port 521 nsew signal output
rlabel metal2 s 188526 159200 188582 160000 6 la_output[47]
port 522 nsew signal output
rlabel metal2 s 192482 159200 192538 160000 6 la_output[48]
port 523 nsew signal output
rlabel metal2 s 196346 159200 196402 160000 6 la_output[49]
port 524 nsew signal output
rlabel metal2 s 20902 159200 20958 160000 6 la_output[4]
port 525 nsew signal output
rlabel metal2 s 200210 159200 200266 160000 6 la_output[50]
port 526 nsew signal output
rlabel metal2 s 204166 159200 204222 160000 6 la_output[51]
port 527 nsew signal output
rlabel metal2 s 208030 159200 208086 160000 6 la_output[52]
port 528 nsew signal output
rlabel metal2 s 211986 159200 212042 160000 6 la_output[53]
port 529 nsew signal output
rlabel metal2 s 215850 159200 215906 160000 6 la_output[54]
port 530 nsew signal output
rlabel metal2 s 219714 159200 219770 160000 6 la_output[55]
port 531 nsew signal output
rlabel metal2 s 223670 159200 223726 160000 6 la_output[56]
port 532 nsew signal output
rlabel metal2 s 227534 159200 227590 160000 6 la_output[57]
port 533 nsew signal output
rlabel metal2 s 231490 159200 231546 160000 6 la_output[58]
port 534 nsew signal output
rlabel metal2 s 235354 159200 235410 160000 6 la_output[59]
port 535 nsew signal output
rlabel metal2 s 24766 159200 24822 160000 6 la_output[5]
port 536 nsew signal output
rlabel metal2 s 239218 159200 239274 160000 6 la_output[60]
port 537 nsew signal output
rlabel metal2 s 243174 159200 243230 160000 6 la_output[61]
port 538 nsew signal output
rlabel metal2 s 247038 159200 247094 160000 6 la_output[62]
port 539 nsew signal output
rlabel metal2 s 250902 159200 250958 160000 6 la_output[63]
port 540 nsew signal output
rlabel metal2 s 254858 159200 254914 160000 6 la_output[64]
port 541 nsew signal output
rlabel metal2 s 258722 159200 258778 160000 6 la_output[65]
port 542 nsew signal output
rlabel metal2 s 262678 159200 262734 160000 6 la_output[66]
port 543 nsew signal output
rlabel metal2 s 266542 159200 266598 160000 6 la_output[67]
port 544 nsew signal output
rlabel metal2 s 270406 159200 270462 160000 6 la_output[68]
port 545 nsew signal output
rlabel metal2 s 274362 159200 274418 160000 6 la_output[69]
port 546 nsew signal output
rlabel metal2 s 28722 159200 28778 160000 6 la_output[6]
port 547 nsew signal output
rlabel metal2 s 278226 159200 278282 160000 6 la_output[70]
port 548 nsew signal output
rlabel metal2 s 282090 159200 282146 160000 6 la_output[71]
port 549 nsew signal output
rlabel metal2 s 286046 159200 286102 160000 6 la_output[72]
port 550 nsew signal output
rlabel metal2 s 289910 159200 289966 160000 6 la_output[73]
port 551 nsew signal output
rlabel metal2 s 293866 159200 293922 160000 6 la_output[74]
port 552 nsew signal output
rlabel metal2 s 297730 159200 297786 160000 6 la_output[75]
port 553 nsew signal output
rlabel metal2 s 301594 159200 301650 160000 6 la_output[76]
port 554 nsew signal output
rlabel metal2 s 305550 159200 305606 160000 6 la_output[77]
port 555 nsew signal output
rlabel metal2 s 309414 159200 309470 160000 6 la_output[78]
port 556 nsew signal output
rlabel metal2 s 313278 159200 313334 160000 6 la_output[79]
port 557 nsew signal output
rlabel metal2 s 32586 159200 32642 160000 6 la_output[7]
port 558 nsew signal output
rlabel metal2 s 317234 159200 317290 160000 6 la_output[80]
port 559 nsew signal output
rlabel metal2 s 321098 159200 321154 160000 6 la_output[81]
port 560 nsew signal output
rlabel metal2 s 325054 159200 325110 160000 6 la_output[82]
port 561 nsew signal output
rlabel metal2 s 328918 159200 328974 160000 6 la_output[83]
port 562 nsew signal output
rlabel metal2 s 332782 159200 332838 160000 6 la_output[84]
port 563 nsew signal output
rlabel metal2 s 336738 159200 336794 160000 6 la_output[85]
port 564 nsew signal output
rlabel metal2 s 340602 159200 340658 160000 6 la_output[86]
port 565 nsew signal output
rlabel metal2 s 344558 159200 344614 160000 6 la_output[87]
port 566 nsew signal output
rlabel metal2 s 348422 159200 348478 160000 6 la_output[88]
port 567 nsew signal output
rlabel metal2 s 352286 159200 352342 160000 6 la_output[89]
port 568 nsew signal output
rlabel metal2 s 36542 159200 36598 160000 6 la_output[8]
port 569 nsew signal output
rlabel metal2 s 356242 159200 356298 160000 6 la_output[90]
port 570 nsew signal output
rlabel metal2 s 360106 159200 360162 160000 6 la_output[91]
port 571 nsew signal output
rlabel metal2 s 363970 159200 364026 160000 6 la_output[92]
port 572 nsew signal output
rlabel metal2 s 367926 159200 367982 160000 6 la_output[93]
port 573 nsew signal output
rlabel metal2 s 371790 159200 371846 160000 6 la_output[94]
port 574 nsew signal output
rlabel metal2 s 375746 159200 375802 160000 6 la_output[95]
port 575 nsew signal output
rlabel metal2 s 379610 159200 379666 160000 6 la_output[96]
port 576 nsew signal output
rlabel metal2 s 383474 159200 383530 160000 6 la_output[97]
port 577 nsew signal output
rlabel metal2 s 387430 159200 387486 160000 6 la_output[98]
port 578 nsew signal output
rlabel metal2 s 391294 159200 391350 160000 6 la_output[99]
port 579 nsew signal output
rlabel metal2 s 40406 159200 40462 160000 6 la_output[9]
port 580 nsew signal output
rlabel metal3 s 0 157496 800 157616 6 mprj_ack_i
port 581 nsew signal input
rlabel metal2 s 504362 159200 504418 160000 6 mprj_adr_o[0]
port 582 nsew signal output
rlabel metal2 s 527730 159200 527786 160000 6 mprj_adr_o[10]
port 583 nsew signal output
rlabel metal2 s 529754 159200 529810 160000 6 mprj_adr_o[11]
port 584 nsew signal output
rlabel metal2 s 531686 159200 531742 160000 6 mprj_adr_o[12]
port 585 nsew signal output
rlabel metal2 s 533618 159200 533674 160000 6 mprj_adr_o[13]
port 586 nsew signal output
rlabel metal2 s 535550 159200 535606 160000 6 mprj_adr_o[14]
port 587 nsew signal output
rlabel metal2 s 537482 159200 537538 160000 6 mprj_adr_o[15]
port 588 nsew signal output
rlabel metal2 s 539506 159200 539562 160000 6 mprj_adr_o[16]
port 589 nsew signal output
rlabel metal2 s 541438 159200 541494 160000 6 mprj_adr_o[17]
port 590 nsew signal output
rlabel metal2 s 543370 159200 543426 160000 6 mprj_adr_o[18]
port 591 nsew signal output
rlabel metal2 s 545302 159200 545358 160000 6 mprj_adr_o[19]
port 592 nsew signal output
rlabel metal2 s 507306 159200 507362 160000 6 mprj_adr_o[1]
port 593 nsew signal output
rlabel metal2 s 547234 159200 547290 160000 6 mprj_adr_o[20]
port 594 nsew signal output
rlabel metal2 s 549166 159200 549222 160000 6 mprj_adr_o[21]
port 595 nsew signal output
rlabel metal2 s 551190 159200 551246 160000 6 mprj_adr_o[22]
port 596 nsew signal output
rlabel metal2 s 553122 159200 553178 160000 6 mprj_adr_o[23]
port 597 nsew signal output
rlabel metal2 s 555054 159200 555110 160000 6 mprj_adr_o[24]
port 598 nsew signal output
rlabel metal2 s 556986 159200 557042 160000 6 mprj_adr_o[25]
port 599 nsew signal output
rlabel metal2 s 558918 159200 558974 160000 6 mprj_adr_o[26]
port 600 nsew signal output
rlabel metal2 s 560942 159200 560998 160000 6 mprj_adr_o[27]
port 601 nsew signal output
rlabel metal2 s 562874 159200 562930 160000 6 mprj_adr_o[28]
port 602 nsew signal output
rlabel metal2 s 564806 159200 564862 160000 6 mprj_adr_o[29]
port 603 nsew signal output
rlabel metal2 s 510250 159200 510306 160000 6 mprj_adr_o[2]
port 604 nsew signal output
rlabel metal2 s 566738 159200 566794 160000 6 mprj_adr_o[30]
port 605 nsew signal output
rlabel metal2 s 568670 159200 568726 160000 6 mprj_adr_o[31]
port 606 nsew signal output
rlabel metal2 s 513102 159200 513158 160000 6 mprj_adr_o[3]
port 607 nsew signal output
rlabel metal2 s 516046 159200 516102 160000 6 mprj_adr_o[4]
port 608 nsew signal output
rlabel metal2 s 517978 159200 518034 160000 6 mprj_adr_o[5]
port 609 nsew signal output
rlabel metal2 s 520002 159200 520058 160000 6 mprj_adr_o[6]
port 610 nsew signal output
rlabel metal2 s 521934 159200 521990 160000 6 mprj_adr_o[7]
port 611 nsew signal output
rlabel metal2 s 523866 159200 523922 160000 6 mprj_adr_o[8]
port 612 nsew signal output
rlabel metal2 s 525798 159200 525854 160000 6 mprj_adr_o[9]
port 613 nsew signal output
rlabel metal2 s 501418 159200 501474 160000 6 mprj_cyc_o
port 614 nsew signal output
rlabel metal3 s 0 11296 800 11416 6 mprj_dat_i[0]
port 615 nsew signal input
rlabel metal3 s 0 56992 800 57112 6 mprj_dat_i[10]
port 616 nsew signal input
rlabel metal3 s 0 61480 800 61600 6 mprj_dat_i[11]
port 617 nsew signal input
rlabel metal3 s 0 66104 800 66224 6 mprj_dat_i[12]
port 618 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 mprj_dat_i[13]
port 619 nsew signal input
rlabel metal3 s 0 75216 800 75336 6 mprj_dat_i[14]
port 620 nsew signal input
rlabel metal3 s 0 79840 800 79960 6 mprj_dat_i[15]
port 621 nsew signal input
rlabel metal3 s 0 84328 800 84448 6 mprj_dat_i[16]
port 622 nsew signal input
rlabel metal3 s 0 88952 800 89072 6 mprj_dat_i[17]
port 623 nsew signal input
rlabel metal3 s 0 93576 800 93696 6 mprj_dat_i[18]
port 624 nsew signal input
rlabel metal3 s 0 98064 800 98184 6 mprj_dat_i[19]
port 625 nsew signal input
rlabel metal3 s 0 15784 800 15904 6 mprj_dat_i[1]
port 626 nsew signal input
rlabel metal3 s 0 102688 800 102808 6 mprj_dat_i[20]
port 627 nsew signal input
rlabel metal3 s 0 107176 800 107296 6 mprj_dat_i[21]
port 628 nsew signal input
rlabel metal3 s 0 111800 800 111920 6 mprj_dat_i[22]
port 629 nsew signal input
rlabel metal3 s 0 116424 800 116544 6 mprj_dat_i[23]
port 630 nsew signal input
rlabel metal3 s 0 120912 800 121032 6 mprj_dat_i[24]
port 631 nsew signal input
rlabel metal3 s 0 125536 800 125656 6 mprj_dat_i[25]
port 632 nsew signal input
rlabel metal3 s 0 130024 800 130144 6 mprj_dat_i[26]
port 633 nsew signal input
rlabel metal3 s 0 134648 800 134768 6 mprj_dat_i[27]
port 634 nsew signal input
rlabel metal3 s 0 139272 800 139392 6 mprj_dat_i[28]
port 635 nsew signal input
rlabel metal3 s 0 143760 800 143880 6 mprj_dat_i[29]
port 636 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 mprj_dat_i[2]
port 637 nsew signal input
rlabel metal3 s 0 148384 800 148504 6 mprj_dat_i[30]
port 638 nsew signal input
rlabel metal3 s 0 152872 800 152992 6 mprj_dat_i[31]
port 639 nsew signal input
rlabel metal3 s 0 25032 800 25152 6 mprj_dat_i[3]
port 640 nsew signal input
rlabel metal3 s 0 29520 800 29640 6 mprj_dat_i[4]
port 641 nsew signal input
rlabel metal3 s 0 34144 800 34264 6 mprj_dat_i[5]
port 642 nsew signal input
rlabel metal3 s 0 38632 800 38752 6 mprj_dat_i[6]
port 643 nsew signal input
rlabel metal3 s 0 43256 800 43376 6 mprj_dat_i[7]
port 644 nsew signal input
rlabel metal3 s 0 47880 800 48000 6 mprj_dat_i[8]
port 645 nsew signal input
rlabel metal3 s 0 52368 800 52488 6 mprj_dat_i[9]
port 646 nsew signal input
rlabel metal2 s 505374 159200 505430 160000 6 mprj_dat_o[0]
port 647 nsew signal output
rlabel metal2 s 528742 159200 528798 160000 6 mprj_dat_o[10]
port 648 nsew signal output
rlabel metal2 s 530674 159200 530730 160000 6 mprj_dat_o[11]
port 649 nsew signal output
rlabel metal2 s 532606 159200 532662 160000 6 mprj_dat_o[12]
port 650 nsew signal output
rlabel metal2 s 534630 159200 534686 160000 6 mprj_dat_o[13]
port 651 nsew signal output
rlabel metal2 s 536562 159200 536618 160000 6 mprj_dat_o[14]
port 652 nsew signal output
rlabel metal2 s 538494 159200 538550 160000 6 mprj_dat_o[15]
port 653 nsew signal output
rlabel metal2 s 540426 159200 540482 160000 6 mprj_dat_o[16]
port 654 nsew signal output
rlabel metal2 s 542358 159200 542414 160000 6 mprj_dat_o[17]
port 655 nsew signal output
rlabel metal2 s 544290 159200 544346 160000 6 mprj_dat_o[18]
port 656 nsew signal output
rlabel metal2 s 546314 159200 546370 160000 6 mprj_dat_o[19]
port 657 nsew signal output
rlabel metal2 s 508226 159200 508282 160000 6 mprj_dat_o[1]
port 658 nsew signal output
rlabel metal2 s 548246 159200 548302 160000 6 mprj_dat_o[20]
port 659 nsew signal output
rlabel metal2 s 550178 159200 550234 160000 6 mprj_dat_o[21]
port 660 nsew signal output
rlabel metal2 s 552110 159200 552166 160000 6 mprj_dat_o[22]
port 661 nsew signal output
rlabel metal2 s 554042 159200 554098 160000 6 mprj_dat_o[23]
port 662 nsew signal output
rlabel metal2 s 556066 159200 556122 160000 6 mprj_dat_o[24]
port 663 nsew signal output
rlabel metal2 s 557998 159200 558054 160000 6 mprj_dat_o[25]
port 664 nsew signal output
rlabel metal2 s 559930 159200 559986 160000 6 mprj_dat_o[26]
port 665 nsew signal output
rlabel metal2 s 561862 159200 561918 160000 6 mprj_dat_o[27]
port 666 nsew signal output
rlabel metal2 s 563794 159200 563850 160000 6 mprj_dat_o[28]
port 667 nsew signal output
rlabel metal2 s 565818 159200 565874 160000 6 mprj_dat_o[29]
port 668 nsew signal output
rlabel metal2 s 511170 159200 511226 160000 6 mprj_dat_o[2]
port 669 nsew signal output
rlabel metal2 s 567750 159200 567806 160000 6 mprj_dat_o[30]
port 670 nsew signal output
rlabel metal2 s 569682 159200 569738 160000 6 mprj_dat_o[31]
port 671 nsew signal output
rlabel metal2 s 514114 159200 514170 160000 6 mprj_dat_o[3]
port 672 nsew signal output
rlabel metal2 s 517058 159200 517114 160000 6 mprj_dat_o[4]
port 673 nsew signal output
rlabel metal2 s 518990 159200 519046 160000 6 mprj_dat_o[5]
port 674 nsew signal output
rlabel metal2 s 520922 159200 520978 160000 6 mprj_dat_o[6]
port 675 nsew signal output
rlabel metal2 s 522854 159200 522910 160000 6 mprj_dat_o[7]
port 676 nsew signal output
rlabel metal2 s 524878 159200 524934 160000 6 mprj_dat_o[8]
port 677 nsew signal output
rlabel metal2 s 526810 159200 526866 160000 6 mprj_dat_o[9]
port 678 nsew signal output
rlabel metal2 s 506294 159200 506350 160000 6 mprj_sel_o[0]
port 679 nsew signal output
rlabel metal2 s 509238 159200 509294 160000 6 mprj_sel_o[1]
port 680 nsew signal output
rlabel metal2 s 512182 159200 512238 160000 6 mprj_sel_o[2]
port 681 nsew signal output
rlabel metal2 s 515126 159200 515182 160000 6 mprj_sel_o[3]
port 682 nsew signal output
rlabel metal2 s 502430 159200 502486 160000 6 mprj_stb_o
port 683 nsew signal output
rlabel metal2 s 570694 159200 570750 160000 6 mprj_wb_iena
port 684 nsew signal output
rlabel metal2 s 503350 159200 503406 160000 6 mprj_we_o
port 685 nsew signal output
rlabel metal2 s 98366 0 98422 800 6 qspi_enabled
port 686 nsew signal output
rlabel metal2 s 577226 0 577282 800 6 ser_rx
port 687 nsew signal input
rlabel metal2 s 566554 0 566610 800 6 ser_tx
port 688 nsew signal output
rlabel metal2 s 529294 0 529350 800 6 spi_csb
port 689 nsew signal output
rlabel metal2 s 534630 0 534686 800 6 spi_enabled
port 690 nsew signal output
rlabel metal2 s 539966 0 540022 800 6 spi_sck
port 691 nsew signal output
rlabel metal2 s 545302 0 545358 800 6 spi_sdi
port 692 nsew signal input
rlabel metal2 s 550546 0 550602 800 6 spi_sdo
port 693 nsew signal output
rlabel metal2 s 555882 0 555938 800 6 spi_sdoenb
port 694 nsew signal output
rlabel metal2 s 295154 0 295210 800 6 sram_ro_addr[0]
port 695 nsew signal input
rlabel metal2 s 300490 0 300546 800 6 sram_ro_addr[1]
port 696 nsew signal input
rlabel metal2 s 305826 0 305882 800 6 sram_ro_addr[2]
port 697 nsew signal input
rlabel metal2 s 311162 0 311218 800 6 sram_ro_addr[3]
port 698 nsew signal input
rlabel metal2 s 316498 0 316554 800 6 sram_ro_addr[4]
port 699 nsew signal input
rlabel metal2 s 321834 0 321890 800 6 sram_ro_addr[5]
port 700 nsew signal input
rlabel metal2 s 327078 0 327134 800 6 sram_ro_addr[6]
port 701 nsew signal input
rlabel metal2 s 332414 0 332470 800 6 sram_ro_addr[7]
port 702 nsew signal input
rlabel metal2 s 284574 0 284630 800 6 sram_ro_clk
port 703 nsew signal input
rlabel metal2 s 289910 0 289966 800 6 sram_ro_csb
port 704 nsew signal input
rlabel metal2 s 337750 0 337806 800 6 sram_ro_data[0]
port 705 nsew signal output
rlabel metal2 s 390926 0 390982 800 6 sram_ro_data[10]
port 706 nsew signal output
rlabel metal2 s 396262 0 396318 800 6 sram_ro_data[11]
port 707 nsew signal output
rlabel metal2 s 401598 0 401654 800 6 sram_ro_data[12]
port 708 nsew signal output
rlabel metal2 s 406934 0 406990 800 6 sram_ro_data[13]
port 709 nsew signal output
rlabel metal2 s 412270 0 412326 800 6 sram_ro_data[14]
port 710 nsew signal output
rlabel metal2 s 417606 0 417662 800 6 sram_ro_data[15]
port 711 nsew signal output
rlabel metal2 s 422850 0 422906 800 6 sram_ro_data[16]
port 712 nsew signal output
rlabel metal2 s 428186 0 428242 800 6 sram_ro_data[17]
port 713 nsew signal output
rlabel metal2 s 433522 0 433578 800 6 sram_ro_data[18]
port 714 nsew signal output
rlabel metal2 s 438858 0 438914 800 6 sram_ro_data[19]
port 715 nsew signal output
rlabel metal2 s 343086 0 343142 800 6 sram_ro_data[1]
port 716 nsew signal output
rlabel metal2 s 444194 0 444250 800 6 sram_ro_data[20]
port 717 nsew signal output
rlabel metal2 s 449530 0 449586 800 6 sram_ro_data[21]
port 718 nsew signal output
rlabel metal2 s 454774 0 454830 800 6 sram_ro_data[22]
port 719 nsew signal output
rlabel metal2 s 460110 0 460166 800 6 sram_ro_data[23]
port 720 nsew signal output
rlabel metal2 s 465446 0 465502 800 6 sram_ro_data[24]
port 721 nsew signal output
rlabel metal2 s 470782 0 470838 800 6 sram_ro_data[25]
port 722 nsew signal output
rlabel metal2 s 476118 0 476174 800 6 sram_ro_data[26]
port 723 nsew signal output
rlabel metal2 s 481454 0 481510 800 6 sram_ro_data[27]
port 724 nsew signal output
rlabel metal2 s 486698 0 486754 800 6 sram_ro_data[28]
port 725 nsew signal output
rlabel metal2 s 492034 0 492090 800 6 sram_ro_data[29]
port 726 nsew signal output
rlabel metal2 s 348422 0 348478 800 6 sram_ro_data[2]
port 727 nsew signal output
rlabel metal2 s 497370 0 497426 800 6 sram_ro_data[30]
port 728 nsew signal output
rlabel metal2 s 502706 0 502762 800 6 sram_ro_data[31]
port 729 nsew signal output
rlabel metal2 s 353758 0 353814 800 6 sram_ro_data[3]
port 730 nsew signal output
rlabel metal2 s 359002 0 359058 800 6 sram_ro_data[4]
port 731 nsew signal output
rlabel metal2 s 364338 0 364394 800 6 sram_ro_data[5]
port 732 nsew signal output
rlabel metal2 s 369674 0 369730 800 6 sram_ro_data[6]
port 733 nsew signal output
rlabel metal2 s 375010 0 375066 800 6 sram_ro_data[7]
port 734 nsew signal output
rlabel metal2 s 380346 0 380402 800 6 sram_ro_data[8]
port 735 nsew signal output
rlabel metal2 s 385682 0 385738 800 6 sram_ro_data[9]
port 736 nsew signal output
rlabel metal2 s 561218 0 561274 800 6 trap
port 737 nsew signal output
rlabel metal2 s 571890 0 571946 800 6 uart_enabled
port 738 nsew signal output
rlabel metal2 s 571614 159200 571670 160000 6 user_irq_ena[0]
port 739 nsew signal output
rlabel metal2 s 572626 159200 572682 160000 6 user_irq_ena[1]
port 740 nsew signal output
rlabel metal2 s 573546 159200 573602 160000 6 user_irq_ena[2]
port 741 nsew signal output
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 580000 160000
string LEFview TRUE
string GDS_FILE /project/openlane/mgmt_core_wrapper/runs/xyzs/results/magic/mgmt_core_wrapper.gds
string GDS_END 179210478
string GDS_START 178062148
<< end >>

