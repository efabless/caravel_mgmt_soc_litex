* NGSPICE file created from RAM128.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dlclkp_1 abstract view
.subckt sky130_fd_sc_hd__dlclkp_1 CLK GATE VGND VNB VPB VPWR GCLK
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_2 abstract view
.subckt sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtp_1 abstract view
.subckt sky130_fd_sc_hd__dlxtp_1 D GATE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

.subckt RAM128 A0[0] A0[1] A0[2] A0[3] A0[4] A0[5] A0[6] CLK Di0[0] Di0[10] Di0[11]
+ Di0[12] Di0[13] Di0[14] Di0[15] Di0[16] Di0[17] Di0[18] Di0[19] Di0[1] Di0[20] Di0[21]
+ Di0[22] Di0[23] Di0[24] Di0[25] Di0[26] Di0[27] Di0[28] Di0[29] Di0[2] Di0[30] Di0[31]
+ Di0[3] Di0[4] Di0[5] Di0[6] Di0[7] Di0[8] Di0[9] Do0[0] Do0[10] Do0[11] Do0[12]
+ Do0[13] Do0[14] Do0[15] Do0[16] Do0[17] Do0[18] Do0[19] Do0[1] Do0[20] Do0[21] Do0[22]
+ Do0[23] Do0[24] Do0[25] Do0[26] Do0[27] Do0[28] Do0[29] Do0[2] Do0[30] Do0[31] Do0[3]
+ Do0[4] Do0[5] Do0[6] Do0[7] Do0[8] Do0[9] EN0 VGND VPWR WE0[0] WE0[1] WE0[2] WE0[3]
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_111_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_91_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_3_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.Do0_REG.Root_CLKBUF BLOCK\[0\].RAM32.CLKBUF.cell/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.Do0_REG.Root_CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xtap_111_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[12\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[30\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_24_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_93_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_138_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_86_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[24\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_40_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_79_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[13\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND4 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND4/X
+ sky130_fd_sc_hd__and4bb_2
Xtap_40_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_40_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_136_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[3\].Do_FF\[1\] BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X
+ BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[3\].MUX\[1\]/A2
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[25\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_136_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_136_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_49_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_49_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[14\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_49_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[23\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[8\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[2\].Do_FF\[6\] BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X
+ BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[2\].MUX\[6\]/A0
+ sky130_fd_sc_hd__dfxtp_1
Xtap_22_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_65_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_65_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.TIE0\[1\].cell VGND VGND VPWR VPWR BLOCK\[0\].RAM32.TIE0\[1\].cell/HI
+ BLOCK\[0\].RAM32.TIE0\[1\].cell/LO sky130_fd_sc_hd__conb_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[9\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_81_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[18\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_141_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_0_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[6\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[15\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell BLOCK\[3\].RAM32.WEBUF\[3\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.A0BUF\[0\].cell A0BUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.A0BUF\[0\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[31\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[27\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_50_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[14\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[5\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_36_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[1\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF BLOCK\[2\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[10\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[28\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_29_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell BLOCK\[1\].RAM32.CLKBUF.cell/X VGND
+ VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[15\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[27\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[11\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_58_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_86_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[10\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_106_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_106_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_19_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[24\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_19_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_122_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_122_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_35_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_35_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[0\].DIODE\[4\] BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_91_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_51_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_51_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_136_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[7\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_84_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_51_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_142_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_129_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_77_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND4/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xfill_128_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[19\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.DIBUF\[20\].cell DIBUF\[20\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DIBUF\[20\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[2\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[20\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[29\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_76_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.ENBUF BLOCK\[3\].RAM32.DEC0.AND2/X VGND VGND
+ VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[3\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[30\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[4\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[2\].DIODE\[1\] BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell BLOCK\[1\].RAM32.TIE0\[1\].cell/LO
+ BLOCK\[1\].RAM32.FBUFENBUF0\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[13\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[31\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[16\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[25\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[14\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[26\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_2_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[9\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[0\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_41_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND4 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND4/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[23\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_122_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF BLOCK\[3\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xtap_21_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_70_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_115_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_63_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_117_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_108_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_97_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_97_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell BLOCK\[1\].RAM32.TIE0\[2\].cell/LO
+ BLOCK\[1\].RAM32.FBUFENBUF0\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_56_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[22\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[6\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_117_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_49_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_69_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_69_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[18\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_133_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_133_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_133_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[23\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[5\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_46_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_46_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_46_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[1\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_106_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[19\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDIBUF\[1\].cell Di0[1] VGND VGND VPWR VPWR DIBUF\[1\].cell/X sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[6\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_62_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_62_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_141_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_62_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[2\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[18\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.FBUFENBUF0\[1\].cell DEC0.AND0/Y VGND VGND VPWR VPWR BLOCK\[0\].RAM32.FBUFENBUF0\[1\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
Xfill_34_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_34_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_134_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_34_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_140_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_133_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[1\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_126_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_119_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[24\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[15\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[1\].DIODE_A3MUX\[13\] Do0MUX.M\[1\].MUX\[5\]/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[1\].Do_FF\[2\] BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X
+ BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[1\].MUX\[2\]/A1
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[27\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[10\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_96_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[11\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[20\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND2/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xfill_89_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell BLOCK\[0\].RAM32.WEBUF\[0\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[21\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_103_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_103_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF BLOCK\[0\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xtap_16_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[4\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[22\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_32_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_71_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_32_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[16\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_120_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[5\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[2\].DIODE_A3MUX\[17\] Do0MUX.M\[2\].MUX\[1\]/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_128_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_128_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_113_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_61_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_106_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[17\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_54_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_47_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_105_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_57_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_57_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_57_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[0\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[31\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_73_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_73_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[14\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[30\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[26\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[13\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[9\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell BLOCK\[2\].RAM32.TIE0\[1\].cell/LO
+ BLOCK\[2\].RAM32.FBUFENBUF0\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[23\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[14\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.DIBUF\[24\].cell DIBUF\[24\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DIBUF\[24\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xfill_68_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[10\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[19\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[9\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[18\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_11_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xtap_8_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_40_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[2\] BLOCK\[1\].RAM32.Do0_REG.Root_CLKBUF/X VGND
+ VGND VPWR VPWR BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X sky130_fd_sc_hd__clkbuf_4
Xtap_33_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[6\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_26_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[0\].DIODE\[2\] BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[15\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_114_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_114_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_94_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[27\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND1 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND1/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_130_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_130_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_43_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_43_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[1\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[10\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_43_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.Do0_REG.Root_CLKBUF BLOCK\[3\].RAM32.CLKBUF.cell/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.Do0_REG.Root_CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[28\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_111_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[11\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[29\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_104_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_52_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_68_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_68_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[12\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_84_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[24\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[13\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[22\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[3\].DIODE\[7\] BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[25\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND5/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.WEBUF\[2\].cell WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.WEBUF\[2\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[8\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell BLOCK\[1\].RAM32.TIE0\[0\].cell/LO
+ BLOCK\[1\].RAM32.FBUFENBUF0\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_66_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[31\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_59_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[5\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[14\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[30\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.ABUF\[2\] BLOCK\[0\].RAM32.A0BUF\[2\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[17\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[26\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_100_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_100_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_7_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_13_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_88_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[31\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_13_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[13\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[4\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[0\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_109_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_109_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_89_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[27\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[14\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_125_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_125_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[1\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[26\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_31_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_38_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[10\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_24_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_38_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_38_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_17_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_141_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_141_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[0\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_54_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_54_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_54_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[9\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XDo0MUX.M\[0\].DIODE_A2MUX\[3\] Do0MUX.M\[0\].MUX\[3\]/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_70_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_70_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[23\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_79_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_139_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_139_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[6\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_139_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_139_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_139_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_101_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[18\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[7\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF BLOCK\[2\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[1\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[19\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_0_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_104_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_104_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[2\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[20\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[29\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_5_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[3\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_5_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[30\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_71_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell BLOCK\[1\].RAM32.WEBUF\[2\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[24\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[13\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[4\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell BLOCK\[0\].RAM32.CLKBUF.cell/X VGND
+ VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.DIBUF\[28\].cell DIBUF\[28\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DIBUF\[28\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xtap_111_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[25\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_111_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_24_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_93_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_138_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[8\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_86_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND3/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_79_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND5 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND5/X
+ sky130_fd_sc_hd__and4b_2
Xtap_40_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_40_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_40_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_136_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_136_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_49_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_49_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[22\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_49_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_22_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_65_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_65_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_65_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[21\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[5\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[17\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_81_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_81_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[22\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[4\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_0_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[0\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[18\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[5\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[1\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[17\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.ABUF\[0\] BLOCK\[2\].RAM32.A0BUF\[0\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[0\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_50_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfill_43_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[31\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell BLOCK\[0\].RAM32.WEBUF\[3\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X sky130_fd_sc_hd__clkbuf_2
Xfill_36_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XA0BUF\[1\].cell A0[1] VGND VGND VPWR VPWR A0BUF\[1\].cell/X sky130_fd_sc_hd__clkbuf_2
Xfill_29_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell BLOCK\[3\].RAM32.TIE0\[3\].cell/LO
+ BLOCK\[3\].RAM32.FBUFENBUF0\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[14\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[3\].MUX\[2\] Do0MUX.M\[3\].MUX\[2\]/A0 Do0MUX.M\[3\].MUX\[2\]/A1 Do0MUX.M\[3\].MUX\[2\]/A2
+ Do0MUX.M\[3\].MUX\[2\]/A3 Do0MUX.SEL0BUF\[3\]/X Do0MUX.SEL1BUF\[3\]/X VGND VGND
+ VPWR VPWR Do0[26] sky130_fd_sc_hd__mux4_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[26\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[15\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_10_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[9\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_106_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_106_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_19_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_122_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_122_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[10\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[19\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF BLOCK\[3\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_35_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_35_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_91_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[20\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_51_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_136_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_84_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_51_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_51_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_142_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_129_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_77_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[3\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[21\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_128_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[3\].DIODE\[5\] BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[4\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[2\].MUX\[4\] Do0MUX.M\[2\].MUX\[4\]/A0 Do0MUX.M\[2\].MUX\[4\]/A1 Do0MUX.M\[2\].MUX\[4\]/A2
+ Do0MUX.M\[2\].MUX\[4\]/A3 Do0MUX.SEL0BUF\[2\]/X Do0MUX.SEL1BUF\[2\]/X VGND VGND
+ VPWR VPWR Do0[20] sky130_fd_sc_hd__mux4_1
Xtap_76_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_76_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[16\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_92_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.DIBUF\[11\].cell DIBUF\[11\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DIBUF\[11\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.DIBUF\[3\].cell DIBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DIBUF\[3\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[30\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND1/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[13\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[29\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[3\].DIODE_A0MUX\[31\] Do0MUX.M\[3\].MUX\[7\]/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[25\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_2_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[12\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF BLOCK\[0\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND6/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[8\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[26\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_41_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[22\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[13\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_34_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[9\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[25\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[1\].MUX\[6\] Do0MUX.M\[1\].MUX\[6\]/A0 Do0MUX.M\[1\].MUX\[6\]/A1 Do0MUX.M\[1\].MUX\[6\]/A2
+ Do0MUX.M\[1\].MUX\[6\]/A3 Do0MUX.SEL0BUF\[1\]/X Do0MUX.SEL1BUF\[1\]/X VGND VGND
+ VPWR VPWR Do0[14] sky130_fd_sc_hd__mux4_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND5 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND5/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_70_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[8\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_21_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_115_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_63_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_117_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_108_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_97_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_56_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_117_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_49_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_69_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell BLOCK\[2\].RAM32.TIE0\[0\].cell/LO
+ BLOCK\[2\].RAM32.FBUFENBUF0\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_133_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_133_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[31\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_46_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_46_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_46_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xfill_106_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[5\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_62_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_62_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_141_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[14\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_62_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[3\].Do_FF\[1\] BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X
+ BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[3\].MUX\[1\]/A3
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[17\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_34_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_34_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_134_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[26\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_82_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_34_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_140_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_127_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[15\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_34_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[2\].Do_FF\[6\] BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X
+ BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[2\].MUX\[6\]/A1
+ sky130_fd_sc_hd__dfxtp_1
Xfill_126_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[0\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[27\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_119_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_87_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[1\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[10\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[28\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[11\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[29\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[12\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[24\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_96_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_89_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XDIBUF\[15\].cell Di0[15] VGND VGND VPWR VPWR DIBUF\[15\].cell/X sky130_fd_sc_hd__clkbuf_16
Xtap_103_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[7\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_103_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_16_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[21\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[30\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_32_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell BLOCK\[0\].RAM32.TIE0\[3\].cell/LO
+ BLOCK\[0\].RAM32.FBUFENBUF0\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_120_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[20\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[4\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_128_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_113_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[29\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_128_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_61_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[16\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[25\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_106_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_54_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[30\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[3\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_47_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.FBUFENBUF0\[0\].cell DEC0.AND1/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.FBUFENBUF0\[0\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_105_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_57_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_57_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_57_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[0\].DIODE\[4\] BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[26\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[4\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF BLOCK\[1\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[13\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_73_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_73_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_73_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[3\].DIODE_A1MUX\[29\] Do0MUX.M\[3\].MUX\[5\]/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[0\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND4/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[25\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[9\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[8\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_131_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[22\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_68_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[5\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[2\].DIODE\[1\] BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[23\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[17\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.DIBUF\[15\].cell DIBUF\[15\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DIBUF\[15\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[1\].DIODE\[6\] BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[6\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_11_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.ABUF\[1\] BLOCK\[1\].RAM32.A0BUF\[1\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[0\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[18\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[7\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[1\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[19\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[28\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_33_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_114_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_114_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[2\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_19_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND2 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND2/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[29\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_130_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_130_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_43_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_43_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[12\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[3\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_43_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[24\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_111_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.DIBUF\[30\].cell DIBUF\[30\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DIBUF\[30\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xtap_104_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[15\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_52_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_68_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_68_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_68_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_45_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_103_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xtap_84_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_84_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[21\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[20\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[4\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[16\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[21\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[3\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[1\].Do_FF\[2\] BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X
+ BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[1\].MUX\[2\]/A2
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[17\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[4\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_66_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_59_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[0\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[16\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[0\].Do_FF\[7\] BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X
+ BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[0\].MUX\[7\]/A0
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_100_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_7_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xtap_13_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_13_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND2/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[30\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_109_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_109_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[13\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_125_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_125_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_38_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[25\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_24_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_38_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_38_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[14\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_17_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_141_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[23\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_141_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[8\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[26\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_54_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_54_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_54_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_70_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[9\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.DIBUF\[6\].cell DIBUF\[6\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DIBUF\[6\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xtap_70_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[7\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_79_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[10\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_79_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[19\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_139_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_139_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_139_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_139_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_139_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_101_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_95_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[20\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[3\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell BLOCK\[3\].RAM32.TIE0\[0\].cell/LO
+ BLOCK\[3\].RAM32.FBUFENBUF0\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_0_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_104_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_104_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_104_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[15\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_5_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[29\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_71_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF BLOCK\[3\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_64_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[12\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[28\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[24\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_111_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_111_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[29\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_24_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[11\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.A0BUF\[3\].cell A0BUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DEC0.AND3/B
+ sky130_fd_sc_hd__clkbuf_2
Xtap_24_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_93_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_138_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[25\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_86_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_79_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND6 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND6/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[12\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_40_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_40_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[0\].DIODE\[2\] BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[8\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[24\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_136_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_136_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_49_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_49_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_49_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_22_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_65_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_65_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_65_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_81_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_81_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.ENBUF BLOCK\[0\].RAM32.DEC0.AND0/Y VGND VGND
+ VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[21\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_81_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[30\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xfill_0_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[4\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND0/Y
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[31\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[16\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[25\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[5\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[14\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[0\] BLOCK\[0\].RAM32.Do0_REG.Root_CLKBUF/X VGND
+ VGND VPWR VPWR BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND5/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[26\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[15\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[0\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_36_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[9\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[27\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_29_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[10\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[28\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_10_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF BLOCK\[0\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[11\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_106_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_106_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_19_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_122_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_122_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_35_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_35_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[23\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_1_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_91_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_51_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XDo0MUX.M\[2\].DIODE_A0MUX\[20\] Do0MUX.M\[2\].MUX\[4\]/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_136_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_84_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[6\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_51_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_51_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_142_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_129_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_77_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[20\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[29\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_128_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[7\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[3\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_76_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[19\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_76_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_76_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[28\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_92_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[29\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[2\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_92_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[16\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[25\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[3\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[12\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[1\].Do_FF\[0\] BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X
+ BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[1\].MUX\[0\]/A0
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[24\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XDo0MUX.M\[3\].DIODE_A0MUX\[24\] Do0MUX.M\[3\].MUX\[0\]/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_41_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_34_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[21\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_27_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND6 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND6/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_142_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[4\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[22\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_21_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[16\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_63_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_108_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_56_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_117_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_117_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[5\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[23\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_49_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[17\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF BLOCK\[1\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xtap_133_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_133_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell BLOCK\[2\].RAM32.TIE0\[2\].cell/LO
+ BLOCK\[2\].RAM32.FBUFENBUF0\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[6\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_46_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_46_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_46_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_106_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND3/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[0\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[18\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_62_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_62_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_62_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_141_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[1\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_34_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[19\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_34_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDo0MUX.M\[1\].DIODE_A1MUX\[14\] Do0MUX.M\[1\].MUX\[6\]/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_134_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_82_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[28\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_34_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_34_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_140_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_127_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.CLKBUF.cell CLKBUF.cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.CLKBUF.cell/X
+ sky130_fd_sc_hd__clkbuf_4
Xtap_75_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBLOCK\[3\].RAM32.WEBUF\[1\].cell WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.WEBUF\[1\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[2\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_119_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[2\] BLOCK\[2\].RAM32.Do0_REG.Root_CLKBUF/X VGND
+ VGND VPWR VPWR BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X sky130_fd_sc_hd__clkbuf_4
Xtap_87_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_87_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[14\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[23\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[11\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[20\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[7\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[19\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[10\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[2\].DIODE_A1MUX\[18\] Do0MUX.M\[2\].MUX\[2\]/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[20\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_103_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_16_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[16\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[3\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_32_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_120_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_128_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_128_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_113_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_61_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_106_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_54_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_47_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[29\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_105_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_3_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_57_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_57_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_57_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[12\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[30\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_73_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_73_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_73_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[24\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[13\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[25\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[3\].DIODE\[5\] BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDIBUF\[21\].cell Di0[21] VGND VGND VPWR VPWR DIBUF\[21\].cell/X sky130_fd_sc_hd__clkbuf_16
Xfill_131_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[14\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[23\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_124_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_98_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[8\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[9\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[18\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell BLOCK\[3\].RAM32.TIE0\[1\].cell/LO
+ BLOCK\[3\].RAM32.FBUFENBUF0\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[19\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND1/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_8_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[2\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_94_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[31\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[5\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_114_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_114_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[14\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_26_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[28\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND3 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND3/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[15\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_130_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_130_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_43_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[27\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_43_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_43_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[11\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XDo0MUX.M\[2\].DIODE_A3MUX\[22\] Do0MUX.M\[2\].MUX\[6\]/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_111_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[28\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[10\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_104_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_52_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_68_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[24\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_68_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_68_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_45_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_103_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[11\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_38_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.DIBUF\[21\].cell DIBUF\[21\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DIBUF\[21\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_84_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_84_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_84_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[2\].Do_FF\[6\] BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X
+ BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[2\].MUX\[6\]/A2
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[3\].RAM32.DIBUF\[26\].cell DIBUF\[26\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DIBUF\[26\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[20\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[29\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XDo0MUX.M\[3\].DIODE_A3MUX\[26\] Do0MUX.M\[3\].MUX\[2\]/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[3\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_66_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[30\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[4\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[13\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[31\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[16\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[25\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_7_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_13_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[14\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_109_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_109_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[26\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.ABUF\[2\] BLOCK\[1\].RAM32.A0BUF\[2\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_125_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_125_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[0\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_31_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[9\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_24_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[27\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_38_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_38_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_141_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_141_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_54_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_54_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[10\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_54_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.DIBUF\[2\].cell DIBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DIBUF\[2\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_70_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_70_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[22\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[0\].DIODE_A0MUX\[2\] Do0MUX.M\[0\].MUX\[2\]/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_79_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_79_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_102_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_79_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_139_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[5\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[23\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDIBUF\[7\].cell Di0[7] VGND VGND VPWR VPWR DIBUF\[7\].cell/X sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_139_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_139_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_139_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_101_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_95_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_95_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[19\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND4/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[6\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[2\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[18\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[7\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_0_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_104_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_104_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_104_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_104_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[28\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[19\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[1\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[24\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[2\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[2\].DIODE\[1\] BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_71_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_64_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[1\].DIODE\[6\] BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_57_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_111_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell BLOCK\[0\].RAM32.TIE0\[1\].cell/LO
+ BLOCK\[0\].RAM32.FBUFENBUF0\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_24_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_93_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_138_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_86_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[11\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_79_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/X
+ sky130_fd_sc_hd__and4_2
Xtap_40_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_40_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[20\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_136_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_136_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_49_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[21\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_49_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_49_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_22_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_65_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_65_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_65_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_15_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[4\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[22\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[3\].DIODE\[3\] BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[16\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_81_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_101_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_81_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_81_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[5\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_0_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[17\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[0\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[18\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[27\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[1\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[30\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.ABUF\[0\] BLOCK\[3\].RAM32.A0BUF\[0\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_36_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[13\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[1\].Do_FF\[2\] BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X
+ BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[1\].MUX\[2\]/A3
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[14\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_10_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF BLOCK\[1\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[23\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[0\].Do_FF\[7\] BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X
+ BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[0\].MUX\[7\]/A1
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[10\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[19\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_106_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_19_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_122_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[18\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[9\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_122_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND2/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_35_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_35_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_1_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[7\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_91_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[19\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_136_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_84_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_51_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_51_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_51_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_142_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_129_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_77_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[2\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_6_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_76_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_76_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_76_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[2\].Do_FF\[4\] BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X
+ BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[2\].MUX\[4\]/A0
+ sky130_fd_sc_hd__dfxtp_1
Xtap_20_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_92_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_92_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[28\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_92_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[11\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[29\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[12\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[24\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[13\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[22\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[25\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_34_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[8\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_27_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/X
+ sky130_fd_sc_hd__and4_2
Xfill_142_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_142_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_21_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[9\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND0/Y
+ sky130_fd_sc_hd__nor4b_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_56_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[18\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_117_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_117_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_49_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_133_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_133_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[30\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_46_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_46_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[4\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_62_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[0\].DIODE\[2\] BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[13\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_62_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_62_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[31\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_141_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[27\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_134_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_82_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_34_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_34_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_140_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_127_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_75_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[14\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_68_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[1\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_126_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.DIBUF\[13\].cell DIBUF\[13\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DIBUF\[13\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[26\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[10\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF BLOCK\[2\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xtap_87_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_87_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_87_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[15\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[0\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[27\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[9\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[10\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND0/Y
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[7\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[19\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_16_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[2\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[20\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[29\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[7\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_32_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[3\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_120_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[30\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_128_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_128_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_113_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_61_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_106_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[24\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_54_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell BLOCK\[1\].RAM32.TIE0\[3\].cell/LO
+ BLOCK\[1\].RAM32.FBUFENBUF0\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[4\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_47_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_105_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[13\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_3_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_57_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_57_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_57_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[25\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_73_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_73_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_73_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[8\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[26\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_132_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[9\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_131_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xtap_98_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_124_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_98_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_117_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[21\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF BLOCK\[3\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[4\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[22\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[1\].DIODE_A3MUX\[11\] Do0MUX.M\[1\].MUX\[3\]/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[1\].Do_FF\[0\] BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X
+ BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[1\].MUX\[0\]/A1
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[18\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[23\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[5\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.A0BUF\[2\].cell A0BUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.A0BUF\[2\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[1\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[17\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[6\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_94_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.ABUF\[1\] BLOCK\[2\].RAM32.A0BUF\[1\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B sky130_fd_sc_hd__clkbuf_2
Xfill_87_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[27\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[18\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[0\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_114_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[1\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_19_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND4 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND4/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_130_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_130_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_43_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_43_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[15\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_111_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_104_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_68_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_52_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_68_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_68_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_45_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[10\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND3/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_38_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[19\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[0\].DIODE_A1MUX\[7\] Do0MUX.M\[0\].MUX\[7\]/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_84_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_84_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_84_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[20\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[7\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[3\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[21\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[4\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF BLOCK\[0\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.DIBUF\[17\].cell DIBUF\[17\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DIBUF\[17\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[16\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.DIBUF\[9\].cell DIBUF\[9\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DIBUF\[9\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xfill_66_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xfill_59_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[17\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[0\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_13_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[29\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_109_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[12\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_125_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_125_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[0\] BLOCK\[1\].RAM32.Do0_REG.Root_CLKBUF/X VGND
+ VGND VPWR VPWR BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X sky130_fd_sc_hd__clkbuf_4
Xtap_31_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[26\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[0\].DIODE\[0\] BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_38_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_38_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[13\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_24_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_0_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[22\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_141_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_141_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_54_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[25\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[9\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_54_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[23\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_70_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_70_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[8\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[6\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_79_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[9\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_102_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_79_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_79_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_50_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[18\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xfill_139_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_139_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_139_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_95_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_95_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_95_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[3\].DIODE\[5\] BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[15\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_104_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_104_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_104_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_104_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_104_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[27\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[1\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[10\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[28\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[15\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_71_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_64_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[11\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND1/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[29\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_57_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[12\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_24_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF BLOCK\[1\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xfill_5_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.ABUF\[0\] BLOCK\[0\].RAM32.A0BUF\[0\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A sky130_fd_sc_hd__clkbuf_2
Xtap_86_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[24\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND6/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_79_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_40_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_40_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_136_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_136_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_49_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_49_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_49_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[7\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_22_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[8\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_65_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_65_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[17\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_65_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_81_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_101_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_101_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_81_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_81_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[20\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[0\].DIODE_A2MUX\[1\] Do0MUX.M\[0\].MUX\[1\]/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_98_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[29\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xfill_0_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[3\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell BLOCK\[0\].RAM32.TIE0\[0\].cell/LO
+ BLOCK\[0\].RAM32.FBUFENBUF0\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[30\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[26\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[4\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[31\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[13\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[2\].Do_FF\[6\] BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X
+ BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[2\].MUX\[6\]/A3
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[0\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[25\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[9\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[14\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_36_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[26\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[8\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[9\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_10_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[2\] BLOCK\[3\].RAM32.Do0_REG.Root_CLKBUF/X VGND
+ VGND VPWR VPWR BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_19_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[23\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_122_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_35_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[6\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_1_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_35_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[18\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_91_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_136_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_51_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_51_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[23\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[7\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_84_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_129_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.DEC0.AND0 BLOCK\[2\].RAM32.DEC0.AND3/B BLOCK\[2\].RAM32.DEC0.AND3/A
+ BLOCK\[2\].RAM32.DEC0.AND3/C VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DEC0.AND0/Y sky130_fd_sc_hd__nor3b_2
Xtap_77_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[1\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[19\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF BLOCK\[2\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xtap_6_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[28\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[6\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[2\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_76_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_76_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_76_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[29\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_20_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_92_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[3\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_112_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_92_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_92_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[12\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[24\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[15\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[25\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[8\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell BLOCK\[1\].RAM32.WEBUF\[0\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[20\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_34_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_142_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfill_142_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_142_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDo0MUX.M\[3\].MUX\[0\] Do0MUX.M\[3\].MUX\[0\]/A0 Do0MUX.M\[3\].MUX\[0\]/A1 Do0MUX.M\[3\].MUX\[0\]/A2
+ Do0MUX.M\[3\].MUX\[0\]/A3 Do0MUX.SEL0BUF\[3\]/X Do0MUX.SEL1BUF\[3\]/X VGND VGND
+ VPWR VPWR Do0[24] sky130_fd_sc_hd__mux4_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[3\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[21\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_21_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[17\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_117_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND1 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND1/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[1\].DIODE\[6\] BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[22\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[4\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_49_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[31\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[0\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[16\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_133_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[5\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_133_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_46_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_46_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[17\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell BLOCK\[3\].RAM32.TIE0\[2\].cell/LO
+ BLOCK\[3\].RAM32.FBUFENBUF0\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_62_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_62_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_141_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[0\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_34_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_134_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_82_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_34_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_140_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_127_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_75_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_68_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[14\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_107_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_87_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_87_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_87_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[23\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[3\].DIODE\[3\] BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XDo0MUX.M\[2\].MUX\[2\] Do0MUX.M\[2\].MUX\[2\]/A0 Do0MUX.M\[2\].MUX\[2\]/A1 Do0MUX.M\[2\].MUX\[2\]/A2
+ Do0MUX.M\[2\].MUX\[2\]/A3 Do0MUX.SEL0BUF\[2\]/X Do0MUX.SEL1BUF\[2\]/X VGND VGND
+ VPWR VPWR Do0[18] sky130_fd_sc_hd__mux4_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[26\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.SEL0BUF\[2\] DEC0.AND3/B VGND VGND VPWR VPWR Do0MUX.SEL0BUF\[2\]/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[9\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[7\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[23\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[10\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[19\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[6\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF BLOCK\[3\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[20\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[3\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_16_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_16_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_32_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[1\].MUX\[4\] Do0MUX.M\[1\].MUX\[4\]/A0 Do0MUX.M\[1\].MUX\[4\]/A1 Do0MUX.M\[1\].MUX\[4\]/A2
+ Do0MUX.M\[1\].MUX\[4\]/A3 Do0MUX.SEL0BUF\[1\]/X Do0MUX.SEL1BUF\[1\]/X VGND VGND
+ VPWR VPWR Do0[12] sky130_fd_sc_hd__mux4_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[15\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[16\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_32_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[0\].Do_FF\[7\] BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X
+ BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[0\].MUX\[7\]/A2
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_128_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_128_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_113_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_61_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_106_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_54_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_47_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND2/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[28\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_3_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_57_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_57_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_57_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[11\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[29\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_73_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_73_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_73_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[25\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[12\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_132_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_80_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[24\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[8\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_125_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF BLOCK\[0\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[13\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_98_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[2\].Do_FF\[4\] BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X
+ BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[2\].MUX\[4\]/A1
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[22\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_124_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_98_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_98_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_117_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XDo0MUX.M\[0\].MUX\[6\] Do0MUX.M\[0\].MUX\[6\]/A0 Do0MUX.M\[0\].MUX\[6\]/A1 Do0MUX.M\[0\].MUX\[6\]/A2
+ Do0MUX.M\[0\].MUX\[6\]/A3 Do0MUX.SEL0BUF\[0\]/X Do0MUX.SEL1BUF\[0\]/X VGND VGND
+ VPWR VPWR Do0[6] sky130_fd_sc_hd__mux4_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[8\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[17\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[31\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[5\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell BLOCK\[3\].RAM32.WEBUF\[1\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[14\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_94_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XDo0MUX.M\[2\].DIODE_A1MUX\[23\] Do0MUX.M\[2\].MUX\[7\]/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDo0MUX.M\[1\].DIODE_A0MUX\[9\] Do0MUX.M\[1\].MUX\[1\]/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_87_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[26\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell BLOCK\[1\].RAM32.TIE0\[0\].cell/LO
+ BLOCK\[1\].RAM32.FBUFENBUF0\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[15\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[31\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_27_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[0\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[9\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[27\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND5 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND5/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[14\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_130_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_43_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_43_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[10\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[28\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_111_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[11\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_104_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_52_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_68_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_68_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_68_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_45_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_38_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[0\].DIODE\[2\] BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[23\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_84_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_84_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[24\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_84_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[3\].DIODE_A1MUX\[27\] Do0MUX.M\[3\].MUX\[3\]/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_120_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[6\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell BLOCK\[0\].RAM32.TIE0\[2\].cell/LO
+ BLOCK\[0\].RAM32.FBUFENBUF0\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[7\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[19\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[28\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.DIBUF\[5\].cell DIBUF\[5\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DIBUF\[5\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[2\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell BLOCK\[2\].RAM32.WEBUF\[2\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND0/Y
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xfill_66_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[29\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_59_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[16\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[25\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[3\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[30\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[12\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_7_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[1\].DIODE\[4\] BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[24\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND5/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_13_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[13\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[25\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_125_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[8\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_31_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_38_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_38_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.ABUF\[2\] BLOCK\[2\].RAM32.A0BUF\[2\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C sky130_fd_sc_hd__clkbuf_2
Xtap_24_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_17_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_141_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_141_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_54_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_54_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[22\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_9_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_70_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_70_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.DIBUF\[23\].cell DIBUF\[23\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DIBUF\[23\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[5\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[23\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_79_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[17\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_102_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_79_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_79_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_50_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[0\].DIODE_A3MUX\[6\] Do0MUX.M\[0\].MUX\[6\]/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[22\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_139_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_139_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[6\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[31\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_43_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_101_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xtap_95_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_95_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_95_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[0\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_115_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[18\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[5\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[1\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[19\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[28\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xfill_104_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_104_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_104_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_104_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_104_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_104_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[2\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XDo0MUX.M\[3\].DIODE_A3MUX\[31\] Do0MUX.M\[3\].MUX\[7\]/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[14\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[23\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[1\].Do_FF\[0\] BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X
+ BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[1\].MUX\[0\]/A2
+ sky130_fd_sc_hd__dfxtp_1
Xfill_71_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[24\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_57_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[0\].Do_FF\[5\] BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X
+ BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[0\].MUX\[5\]/A0
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_24_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[7\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_5_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[10\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_79_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell BLOCK\[1\].RAM32.TIE0\[1\].cell/LO
+ BLOCK\[1\].RAM32.FBUFENBUF0\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_40_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_40_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[19\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_136_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_136_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_49_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_49_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[20\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_22_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[16\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_65_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_65_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_65_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_15_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[21\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[3\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_8_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_101_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_101_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_81_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_81_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_81_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[4\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_101_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_98_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_0_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[16\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[30\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[13\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDIBUF\[27\].cell Di0[27] VGND VGND VPWR VPWR DIBUF\[27\].cell/X sky130_fd_sc_hd__clkbuf_16
Xfill_36_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[25\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[14\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[23\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[8\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[13\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[22\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[9\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[18\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_19_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_62_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[19\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_35_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_35_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[2\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_91_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_51_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_51_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_136_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[31\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_84_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_129_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.DEC0.AND1 BLOCK\[2\].RAM32.DEC0.AND3/A BLOCK\[2\].RAM32.DEC0.AND3/B
+ BLOCK\[2\].RAM32.DEC0.AND3/C VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DEC0.AND1/X sky130_fd_sc_hd__and3b_2
Xtap_77_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[0\].DIODE\[0\] BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_6_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[5\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[14\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_76_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_76_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[15\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_76_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_20_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_13_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_92_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_112_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_112_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_92_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_92_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[27\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell BLOCK\[2\].RAM32.TIE0\[0\].cell/LO
+ BLOCK\[2\].RAM32.FBUFENBUF0\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_6_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.TIE0\[2\].cell VGND VGND VPWR VPWR BLOCK\[2\].RAM32.TIE0\[2\].cell/HI
+ BLOCK\[2\].RAM32.TIE0\[2\].cell/LO sky130_fd_sc_hd__conb_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[10\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[28\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF BLOCK\[3\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[24\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.DIBUF\[27\].cell DIBUF\[27\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DIBUF\[27\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[11\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[12\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[21\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.WEBUF\[0\].cell WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.WEBUF\[0\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[24\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_34_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_142_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_142_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_142_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND2 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND2/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[30\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND1/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_133_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[4\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[13\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_46_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[31\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_46_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[16\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[25\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XDIBUF\[10\].cell Di0[10] VGND VGND VPWR VPWR DIBUF\[10\].cell/X sky130_fd_sc_hd__clkbuf_16
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND6/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[14\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_62_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_62_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[30\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_141_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_134_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[26\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_82_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_34_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_140_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_127_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[13\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_34_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_75_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[0\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_68_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[9\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[27\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_107_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_87_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_87_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_87_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell BLOCK\[0\].RAM32.TIE0\[3\].cell/LO
+ BLOCK\[0\].RAM32.FBUFENBUF0\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_107_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.DIBUF\[8\].cell DIBUF\[8\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DIBUF\[8\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[10\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_123_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF BLOCK\[0\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[22\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[5\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[23\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[6\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[18\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[7\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_16_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_32_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[1\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[19\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_25_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[28\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_32_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[24\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[2\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[29\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_128_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_61_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.DIBUF\[10\].cell DIBUF\[10\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DIBUF\[10\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_106_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_54_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell BLOCK\[1\].RAM32.WEBUF\[0\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[3\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_47_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_3_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[12\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_57_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_57_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[24\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell BLOCK\[2\].RAM32.TIE0\[3\].cell/LO
+ BLOCK\[2\].RAM32.FBUFENBUF0\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.DIBUF\[15\].cell DIBUF\[15\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DIBUF\[15\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xtap_73_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_73_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_73_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XDo0MUX.M\[1\].DIODE_A1MUX\[12\] Do0MUX.M\[1\].MUX\[4\]/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_132_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_80_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_125_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_73_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_118_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_98_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[21\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_118_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_98_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_98_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[0\] BLOCK\[2\].RAM32.Do0_REG.Root_CLKBUF/X VGND
+ VGND VPWR VPWR BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[4\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[22\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[16\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[21\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[5\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[17\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND4/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[4\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF BLOCK\[1\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[0\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[18\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[27\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_94_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_87_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[1\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XDo0MUX.M\[2\].DIODE_A1MUX\[16\] Do0MUX.M\[2\].MUX\[0\]/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[30\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell BLOCK\[0\].RAM32.WEBUF\[1\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X sky130_fd_sc_hd__clkbuf_2
Xtap_27_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.ABUF\[1\] BLOCK\[3\].RAM32.A0BUF\[1\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B sky130_fd_sc_hd__clkbuf_2
Xtap_27_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND6 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND6/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[13\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_43_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_43_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[1\].DIODE\[6\] BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[14\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[23\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_111_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_104_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_52_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_68_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_68_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_45_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[9\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_38_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[18\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_84_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[7\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_84_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_84_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[19\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_120_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_120_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[20\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[2\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[3\].DIODE\[3\] BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[3\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_122_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.DIBUF\[1\].cell DIBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DIBUF\[1\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[29\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[12\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[1\].DIODE_A2MUX\[8\] Do0MUX.M\[1\].MUX\[0\]/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell BLOCK\[3\].RAM32.TIE0\[0\].cell/LO
+ BLOCK\[3\].RAM32.FBUFENBUF0\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[24\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_92_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[13\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[22\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[25\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_38_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_38_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[12\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_24_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[21\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_17_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_141_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[0\].Do_FF\[7\] BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X
+ BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[0\].MUX\[7\]/A3
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[8\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_54_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_54_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_9_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell BLOCK\[3\].RAM32.WEBUF\[1\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X sky130_fd_sc_hd__clkbuf_2
Xtap_70_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_70_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[9\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_9_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[18\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XDo0MUX.M\[2\].DIODE_A3MUX\[20\] Do0MUX.M\[2\].MUX\[4\]/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_102_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_79_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_79_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_79_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_50_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_139_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[30\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_43_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_101_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_95_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_95_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_36_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_115_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_115_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_95_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[4\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[13\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[31\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_131_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[2\].Do_FF\[4\] BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X
+ BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[2\].MUX\[4\]/A2
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[14\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.DIBUF\[19\].cell DIBUF\[19\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DIBUF\[19\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xfill_104_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_104_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_104_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_104_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_104_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_104_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[26\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[15\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[0\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[9\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[27\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_71_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XDo0MUX.M\[3\].DIODE_A3MUX\[24\] Do0MUX.M\[3\].MUX\[0\]/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_64_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[28\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[10\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[11\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_24_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_40_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_40_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.ABUF\[0\] BLOCK\[1\].RAM32.A0BUF\[0\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A sky130_fd_sc_hd__clkbuf_2
Xtap_136_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell BLOCK\[2\].RAM32.WEBUF\[2\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_49_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_49_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_22_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_65_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[20\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_65_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[29\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[7\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_8_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF BLOCK\[3\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xtap_101_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_101_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_81_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_81_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_81_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[3\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_101_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_98_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[30\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[24\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[4\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[0\].DIODE_A0MUX\[0\] Do0MUX.M\[0\].MUX\[0\]/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[13\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[29\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_100_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[25\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[3\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_126_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[12\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell BLOCK\[0\].RAM32.CLKBUF.cell/X VGND
+ VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[8\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[26\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_36_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[9\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND0/Y
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[21\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[4\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_19_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[22\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_62_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[1\].DIODE\[4\] BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_55_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell BLOCK\[1\].RAM32.WEBUF\[3\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND5/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[5\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[23\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_35_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_35_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[17\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_91_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_51_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_51_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_136_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_84_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[6\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_129_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.DEC0.AND2 BLOCK\[2\].RAM32.DEC0.AND3/B BLOCK\[2\].RAM32.DEC0.AND3/A
+ BLOCK\[2\].RAM32.DEC0.AND3/C VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DEC0.AND2/X sky130_fd_sc_hd__and3b_2
Xtap_77_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[0\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[18\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_6_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[7\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[27\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[1\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_76_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_76_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[28\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_20_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF BLOCK\[0\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[2\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_112_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_112_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_112_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_92_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_92_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_92_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[11\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[3\].DIODE\[1\] BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_6_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[20\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[7\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[3\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[21\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_34_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_142_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_142_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_142_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_142_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[20\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XWEBUF\[1\].cell WE0[1] VGND VGND VPWR VPWR WEBUF\[1\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[4\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[1\].Do_FF\[0\] BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X
+ BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[1\].MUX\[0\]/A3
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[16\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND3 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND3/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[3\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[0\].Do_FF\[5\] BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X
+ BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[0\].MUX\[5\]/A1
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[17\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_46_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_46_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[0\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[29\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_62_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_62_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_141_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_134_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_34_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_82_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_140_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_127_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[12\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_75_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_68_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_107_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_107_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_87_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_87_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_87_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[13\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_107_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[22\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[2\].Do_FF\[2\] BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X
+ BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[2\].MUX\[2\]/A0
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[25\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_123_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_123_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[23\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[8\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF BLOCK\[1\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND3/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[6\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[9\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[18\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[7\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[19\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[2\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.TIE0\[2\].cell VGND VGND VPWR VPWR BLOCK\[0\].RAM32.TIE0\[2\].cell/HI
+ BLOCK\[0\].RAM32.TIE0\[2\].cell/LO sky130_fd_sc_hd__conb_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_32_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfill_25_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfill_18_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell BLOCK\[0\].RAM32.TIE0\[3\].cell/LO
+ BLOCK\[0\].RAM32.FBUFENBUF0\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[28\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[15\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_54_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[11\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[29\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.A0BUF\[1\].cell A0BUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.A0BUF\[1\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
Xtap_3_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_47_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_57_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_57_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[28\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[12\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_73_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_73_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[24\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.ABUF\[1\] BLOCK\[0\].RAM32.A0BUF\[1\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[0\].DIODE\[0\] BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[11\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_132_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_80_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_125_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_73_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_22_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_118_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_118_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_98_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_98_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_98_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_66_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_118_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[8\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[17\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_134_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[20\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[29\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[3\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[30\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[4\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[13\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_94_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[31\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.DIBUF\[21\].cell DIBUF\[21\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DIBUF\[21\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xfill_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[25\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[14\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_27_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[8\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[26\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/X
+ sky130_fd_sc_hd__and4_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[15\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF BLOCK\[2\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xtap_43_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_43_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[27\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[9\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell BLOCK\[1\].RAM32.TIE0\[1\].cell/LO
+ BLOCK\[1\].RAM32.FBUFENBUF0\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[10\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_111_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_104_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_52_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_68_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_68_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_45_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_38_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND6/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_84_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_84_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_17_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[7\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_120_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_120_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[23\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_120_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[19\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_130_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[28\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[6\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_129_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell BLOCK\[1\].RAM32.TIE0\[2\].cell/LO
+ BLOCK\[1\].RAM32.FBUFENBUF0\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[2\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_122_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_115_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[29\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[7\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[3\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[12\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[28\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[24\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[2\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDIBUF\[2\].cell Di0[2] VGND VGND VPWR VPWR DIBUF\[2\].cell/X sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[11\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.FBUFENBUF0\[2\].cell DEC0.AND0/Y VGND VGND VPWR VPWR BLOCK\[0\].RAM32.FBUFENBUF0\[2\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[25\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[8\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_92_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_85_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_38_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_38_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[20\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_17_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_0_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_54_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_54_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.ABUF\[2\] BLOCK\[3\].RAM32.A0BUF\[2\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[3\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[21\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_9_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND0/Y
+ sky130_fd_sc_hd__nor4b_2
Xtap_70_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_70_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[4\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[22\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[31\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_79_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_79_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_79_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[16\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_102_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_50_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell BLOCK\[0\].RAM32.WEBUF\[1\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[5\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_43_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_115_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_95_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_95_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_36_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_115_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_115_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_95_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[17\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_29_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XDo0MUX.M\[0\].DIODE_A1MUX\[5\] Do0MUX.M\[0\].MUX\[5\]/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[6\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[15\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_131_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[0\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_131_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[27\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[18\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_104_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_104_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_104_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_104_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_104_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[1\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xfill_71_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND4/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[7\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[23\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[10\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[19\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[6\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_40_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[20\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[7\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_49_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_49_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[19\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell BLOCK\[2\].RAM32.TIE0\[1\].cell/LO
+ BLOCK\[2\].RAM32.FBUFENBUF0\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[3\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.DIBUF\[25\].cell DIBUF\[25\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DIBUF\[25\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xtap_65_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_65_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[2\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_15_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_8_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_101_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_81_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_81_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[16\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_101_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_101_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_98_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[28\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_30_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_100_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_126_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_126_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[11\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[29\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[12\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_36_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[3\].DIODE\[3\] BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[24\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[13\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[22\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[23\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[8\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[17\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_62_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[6\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_55_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_48_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[18\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_35_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[1\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_51_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_84_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_51_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_129_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_77_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.WEBUF\[3\].cell WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.WEBUF\[3\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.DEC0.AND3 BLOCK\[2\].RAM32.DEC0.AND3/A BLOCK\[2\].RAM32.DEC0.AND3/B
+ BLOCK\[2\].RAM32.DEC0.AND3/C VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DEC0.AND3/X sky130_fd_sc_hd__and3_2
Xtap_6_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[15\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[31\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_76_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[27\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_76_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[14\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_13_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[10\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_112_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_112_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[28\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_92_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_92_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_112_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND2/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[15\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_25_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_96_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[27\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[11\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[10\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_137_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell BLOCK\[2\].RAM32.TIE0\[1\].cell/LO
+ BLOCK\[2\].RAM32.FBUFENBUF0\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[24\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF BLOCK\[1\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[2\].Do_FF\[4\] BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X
+ BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[2\].MUX\[4\]/A3
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.ENBUF BLOCK\[0\].RAM32.DEC0.AND3/X VGND VGND
+ VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_34_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[7\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_142_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_142_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_1_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_142_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_142_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_142_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[19\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[28\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[0\] BLOCK\[3\].RAM32.Do0_REG.Root_CLKBUF/X VGND
+ VGND VPWR VPWR BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND4 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND4/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[2\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[29\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[3\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[12\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[30\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_46_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_46_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[24\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_62_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_62_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[13\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[31\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_141_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[3\].Do_FF\[6\] BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X
+ BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[3\].MUX\[6\]/A0
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[25\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_34_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_34_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_134_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_82_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_127_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_75_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[14\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_68_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[26\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[8\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_107_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_87_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_87_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_107_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_107_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_87_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell BLOCK\[1\].RAM32.WEBUF\[3\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[9\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_123_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_123_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_123_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell BLOCK\[1\].RAM32.TIE0\[3\].cell/LO
+ BLOCK\[1\].RAM32.FBUFENBUF0\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_11_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.DIBUF\[29\].cell DIBUF\[29\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DIBUF\[29\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[23\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[6\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[31\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[22\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[18\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[5\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[1\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[19\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[28\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF BLOCK\[2\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[15\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[6\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[2\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[18\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_32_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[27\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_25_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_18_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[1\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[1\].DIODE\[4\] BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[24\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND5/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_47_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_57_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_57_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_73_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_73_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[7\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XA0BUF\[2\].cell A0[2] VGND VGND VPWR VPWR A0BUF\[2\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[10\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell BLOCK\[3\].RAM32.TIE0\[3\].cell/LO
+ BLOCK\[3\].RAM32.FBUFENBUF0\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[19\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_132_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_80_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_125_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_22_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_73_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_118_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_118_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_118_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_98_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_98_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_98_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[20\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_66_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_118_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_59_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[3\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[3\].DIODE\[1\] BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[21\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XDo0MUX.M\[2\].MUX\[0\] Do0MUX.M\[2\].MUX\[0\]/A0 Do0MUX.M\[2\].MUX\[0\]/A1 Do0MUX.M\[2\].MUX\[0\]/A2
+ Do0MUX.M\[2\].MUX\[0\]/A3 Do0MUX.SEL0BUF\[2\]/X Do0MUX.SEL1BUF\[2\]/X VGND VGND
+ VPWR VPWR Do0[16] sky130_fd_sc_hd__mux4_1
Xtap_134_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_134_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.SEL0BUF\[0\] DEC0.AND3/B VGND VGND VPWR VPWR Do0MUX.SEL0BUF\[0\]/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[4\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[31\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[22\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[16\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[5\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[26\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[17\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_94_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_87_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[0\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.DIBUF\[12\].cell DIBUF\[12\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DIBUF\[12\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[14\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.DIBUF\[4\].cell DIBUF\[4\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DIBUF\[4\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xfill_30_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[23\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_43_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XDo0MUX.M\[1\].MUX\[2\] Do0MUX.M\[1\].MUX\[2\]/A0 Do0MUX.M\[1\].MUX\[2\]/A1 Do0MUX.M\[1\].MUX\[2\]/A2
+ Do0MUX.M\[1\].MUX\[2\]/A3 Do0MUX.SEL0BUF\[1\]/X Do0MUX.SEL1BUF\[1\]/X VGND VGND
+ VPWR VPWR Do0[10] sky130_fd_sc_hd__mux4_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[13\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[0\].Do_FF\[5\] BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X
+ BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[0\].MUX\[5\]/A2
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[22\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[9\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_111_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[18\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_104_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_52_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[23\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_68_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_68_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_45_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[19\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_38_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[6\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_84_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_84_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF BLOCK\[3\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[18\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_17_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[2\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_120_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_120_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_120_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[1\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_33_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_130_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_129_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_129_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_123_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[2\].Do_FF\[2\] BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X
+ BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[2\].MUX\[2\]/A1
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_122_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xfill_115_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[15\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.ENBUF BLOCK\[1\].RAM32.DEC0.AND2/X VGND VGND
+ VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D sky130_fd_sc_hd__clkbuf_2
XDo0MUX.M\[0\].MUX\[4\] Do0MUX.M\[0\].MUX\[4\]/A0 Do0MUX.M\[0\].MUX\[4\]/A1 Do0MUX.M\[0\].MUX\[4\]/A2
+ Do0MUX.M\[0\].MUX\[4\]/A3 Do0MUX.SEL0BUF\[0\]/X Do0MUX.SEL1BUF\[0\]/X VGND VGND
+ VPWR VPWR Do0[4] sky130_fd_sc_hd__mux4_1
Xfill_108_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell BLOCK\[2\].RAM32.TIE0\[0\].cell/LO
+ BLOCK\[2\].RAM32.FBUFENBUF0\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[27\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND3/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[10\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[28\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[11\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_92_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[12\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[21\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XDo0MUX.M\[2\].DIODE_A1MUX\[21\] Do0MUX.M\[2\].MUX\[5\]/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_85_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfill_78_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[24\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_38_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF BLOCK\[0\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[22\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_0_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_54_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_54_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND1 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND1/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[5\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_70_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[8\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_70_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[17\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_79_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_79_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_102_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_50_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_43_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[31\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_95_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDIBUF\[16\].cell Di0[16] VGND VGND VPWR VPWR DIBUF\[16\].cell/X sky130_fd_sc_hd__clkbuf_16
Xtap_36_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_115_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_115_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_115_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_95_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_95_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[0\].DIODE\[0\] BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_28_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[14\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[30\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_131_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_131_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[3\].DIODE_A1MUX\[25\] Do0MUX.M\[3\].MUX\[1\]/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_131_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[26\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[13\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_104_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_104_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[31\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_104_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_104_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_104_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[0\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[9\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[27\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[14\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[26\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[10\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.FBUFENBUF0\[1\].cell DEC0.AND1/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.FBUFENBUF0\[1\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
Xfill_71_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[9\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[1\].DIODE\[2\] BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[23\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[6\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_49_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_49_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[1\].DIODE_A2MUX\[15\] Do0MUX.M\[1\].MUX\[7\]/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[18\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[7\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.ABUF\[0\] BLOCK\[2\].RAM32.A0BUF\[0\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A sky130_fd_sc_hd__clkbuf_2
Xtap_22_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[1\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[19\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_65_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_65_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[28\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND1/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_101_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_81_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_81_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_8_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.DIBUF\[16\].cell DIBUF\[16\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DIBUF\[16\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_101_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_101_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[2\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_14_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_98_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[29\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_14_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[3\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND6/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[12\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_30_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[30\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_100_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[0\].DIODE_A3MUX\[4\] Do0MUX.M\[0\].MUX\[4\]/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_126_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[24\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_126_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_126_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_41_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[13\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[25\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XDo0MUX.M\[2\].DIODE_A2MUX\[19\] Do0MUX.M\[2\].MUX\[3\]/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[8\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.DIBUF\[31\].cell DIBUF\[31\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DIBUF\[31\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[22\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[5\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[21\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_55_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[17\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[0\].Do_FF\[3\] BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X
+ BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[0\].MUX\[3\]/A0
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_48_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[22\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[4\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[31\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[0\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[18\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_51_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[27\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[5\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_77_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[1\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[17\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_6_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_6_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[26\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[0\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_76_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_76_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_112_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_112_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_92_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_92_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_112_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[14\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[23\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_96_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_89_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_41_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_137_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[9\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_137_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[18\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.ENBUF BLOCK\[2\].RAM32.DEC0.AND1/X VGND VGND
+ VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[7\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF BLOCK\[2\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[19\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[2\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[20\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_34_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_142_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_142_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.DIBUF\[7\].cell DIBUF\[7\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DIBUF\[7\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xfill_1_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_1_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfill_142_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_142_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_142_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_142_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[3\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[30\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[21\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND5 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND5/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[4\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND4/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[16\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_60_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_46_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell BLOCK\[3\].RAM32.TIE0\[0\].cell/LO
+ BLOCK\[3\].RAM32.FBUFENBUF0\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_62_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_62_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_141_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_134_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_82_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[13\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_127_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_75_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[22\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_68_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[25\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_107_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_87_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_87_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[12\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_107_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_107_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[21\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[8\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_123_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_123_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[22\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_123_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_36_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[9\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[18\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_4_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[5\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.A0BUF\[4\].cell A0BUF\[4\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DEC0.AND3/A
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[8\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[17\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_138_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[31\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[14\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_32_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[26\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[15\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_18_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[0\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[9\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[27\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell BLOCK\[1\].RAM32.TIE0\[3\].cell/LO
+ BLOCK\[1\].RAM32.FBUFENBUF0\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[10\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[28\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_57_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF BLOCK\[3\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xtap_57_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[11\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_73_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_73_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[12\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[21\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_132_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_80_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_125_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_73_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.ABUF\[1\] BLOCK\[1\].RAM32.A0BUF\[1\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B sky130_fd_sc_hd__clkbuf_2
Xtap_118_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_118_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_98_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_98_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_66_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_118_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_118_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_59_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[16\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_134_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_134_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_134_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[7\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND2/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[30\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[4\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[13\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[29\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[25\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[12\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[3\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_94_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[30\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[8\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[26\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[13\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[25\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[9\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.DIBUF\[0\].cell DIBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DIBUF\[0\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_30_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[8\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_23_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_104_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_52_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF BLOCK\[0\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[22\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_68_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_68_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_45_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_38_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[5\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[23\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_84_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_84_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[3\].Do_FF\[6\] BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X
+ BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[3\].MUX\[6\]/A1
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_17_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[17\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_120_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[6\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_120_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_120_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[0\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[18\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_33_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[1\].DIODE_A1MUX\[10\] Do0MUX.M\[1\].MUX\[2\]/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_130_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[27\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_129_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_129_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_123_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_71_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[7\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_129_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_116_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.ENBUF BLOCK\[3\].RAM32.DEC0.AND0/Y VGND VGND
+ VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D sky130_fd_sc_hd__clkbuf_2
Xfill_122_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[1\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[28\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_115_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_108_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[2\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell BLOCK\[2\].RAM32.TIE0\[2\].cell/LO
+ BLOCK\[2\].RAM32.FBUFENBUF0\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[11\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[29\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[12\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[24\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.WEBUF\[2\].cell WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.WEBUF\[2\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
Xfill_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_85_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_78_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[7\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[21\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_0_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND0/Y
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_54_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_0_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[4\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND2 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND2/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[20\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_70_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[1\].DIODE\[4\] BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[16\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_70_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND5/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[21\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[3\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell BLOCK\[3\].RAM32.CLKBUF.cell/X VGND
+ VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[30\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_79_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_79_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_102_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[17\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_50_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[4\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_43_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_95_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_36_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF BLOCK\[1\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xtap_115_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_115_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_115_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[0\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_95_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[16\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_28_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_131_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_131_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_131_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_44_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_104_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_104_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_104_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_104_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_104_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[3\].DIODE\[1\] BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[13\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[22\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_120_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[25\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[2\].DIODE\[6\] BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[23\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_71_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[8\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[6\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[9\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[18\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[7\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDIBUF\[22\].cell Di0[22] VGND VGND VPWR VPWR DIBUF\[22\].cell/X sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[19\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_90_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_49_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[2\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[20\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_22_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_65_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_65_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[3\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[0\].Do_FF\[5\] BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X
+ BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[0\].MUX\[5\]/A3
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell BLOCK\[3\].RAM32.TIE0\[1\].cell/LO
+ BLOCK\[3\].RAM32.FBUFENBUF0\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_81_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_101_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_101_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_101_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_81_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_98_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[15\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_30_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[29\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_100_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_126_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_126_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_126_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_41_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[12\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_34_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[28\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[24\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[11\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.FBUFENBUF0\[0\].cell DEC0.AND2/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.FBUFENBUF0\[0\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[2\].Do_FF\[2\] BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X
+ BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[2\].MUX\[2\]/A2
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[21\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[12\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[1\].Do_FF\[7\] BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X
+ BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[1\].MUX\[7\]/A0
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[8\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[17\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND3/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[16\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.DIBUF\[22\].cell DIBUF\[22\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DIBUF\[22\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_48_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[30\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.DIBUF\[27\].cell DIBUF\[27\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DIBUF\[27\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xfill_3_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[4\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[13\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[31\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_6_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[25\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_6_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[14\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[8\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[26\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_76_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_76_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[15\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_20_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_112_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_92_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_92_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[9\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[27\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_112_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_112_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_6_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_96_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[10\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_89_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_41_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_41_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_137_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[11\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_137_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_137_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[20\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[23\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_34_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.DIBUF\[3\].cell DIBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DIBUF\[3\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[6\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_142_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_142_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_142_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_142_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_142_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_142_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[29\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[7\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND6 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND6/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[3\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[12\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XDIBUF\[8\].cell Di0[8] VGND VGND VPWR VPWR DIBUF\[8\].cell/X sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[28\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF BLOCK\[3\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[24\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_60_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[11\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[2\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[1\].DIODE\[2\] BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_53_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[29\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[25\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_62_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[12\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[24\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_34_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_134_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[8\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_82_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_127_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_75_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_68_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_87_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_107_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_107_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_107_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_87_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND1/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_123_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_123_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_11_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_123_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[21\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_36_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell BLOCK\[0\].RAM32.TIE0\[1\].cell/LO
+ BLOCK\[0\].RAM32.FBUFENBUF0\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_4_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.A0BUF\[0\].cell A0BUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.A0BUF\[0\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[4\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell BLOCK\[2\].RAM32.TIE0\[3\].cell/LO
+ BLOCK\[2\].RAM32.FBUFENBUF0\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[22\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[31\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_52_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.DIBUF\[10\].cell DIBUF\[10\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DIBUF\[10\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[16\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_138_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[5\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[17\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[6\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[15\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[0\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[18\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[27\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[1\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_32_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xfill_25_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[28\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF BLOCK\[0\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[2\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[11\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[0\].Do_FF\[3\] BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X
+ BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[0\].MUX\[3\]/A1
+ sky130_fd_sc_hd__dfxtp_1
Xtap_3_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[23\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_57_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_73_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_73_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[6\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[20\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[7\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_132_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_80_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_125_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_73_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[3\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_118_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_118_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_98_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_98_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_66_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[19\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_118_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_118_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_59_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[20\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[2\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_134_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_134_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_134_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[2\].Do_FF\[0\] BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X
+ BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[2\].MUX\[0\]/A0
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_47_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[16\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[3\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[29\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[12\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[24\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[13\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[22\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_30_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_23_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfill_16_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND4/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[23\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[8\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[17\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF BLOCK\[1\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xtap_68_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[6\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_52_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_68_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_45_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[18\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_38_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_84_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_84_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_17_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[1\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[19\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_120_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_120_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_120_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[2\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_33_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_130_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_129_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_129_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_123_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[31\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_71_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_129_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_116_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_64_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_122_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_109_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[14\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_108_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[28\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[15\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.TIE0\[0\].cell VGND VGND VPWR VPWR BLOCK\[3\].RAM32.TIE0\[0\].cell/HI
+ BLOCK\[3\].RAM32.TIE0\[0\].cell/LO sky130_fd_sc_hd__conb_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[11\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[27\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[10\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.DIBUF\[14\].cell DIBUF\[14\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DIBUF\[14\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[24\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[20\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[11\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_78_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_0_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_0_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND3 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND3/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_9_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_70_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[29\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_79_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_79_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_102_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_50_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[3\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_43_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[12\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[30\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_115_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_115_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_95_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_95_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_36_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_115_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[24\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_28_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[13\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_131_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[31\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_131_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_131_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_44_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[25\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_44_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_104_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[14\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_104_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_104_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_104_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_104_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[8\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_60_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[26\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND2/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xfill_120_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_113_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF BLOCK\[2\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[9\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[27\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_71_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[10\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[22\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[31\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[5\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xfill_90_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[19\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_83_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[28\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[6\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[15\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_65_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_15_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[18\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[2\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[27\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.ABUF\[0\] BLOCK\[3\].RAM32.A0BUF\[0\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A sky130_fd_sc_hd__clkbuf_2
Xtap_81_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_101_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_101_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_81_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_14_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[1\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.A0BUF\[3\].cell A0BUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DEC0.AND3/B
+ sky130_fd_sc_hd__clkbuf_2
Xtap_98_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_14_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[28\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_14_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[24\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[2\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[11\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_30_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell BLOCK\[0\].RAM32.TIE0\[2\].cell/LO
+ BLOCK\[0\].RAM32.FBUFENBUF0\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[3\].Do_FF\[6\] BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X
+ BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[3\].MUX\[6\]/A2
+ sky130_fd_sc_hd__dfxtp_1
Xtap_100_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_126_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_126_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_126_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_41_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_34_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_27_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[0\].DIODE_A1MUX\[3\] Do0MUX.M\[0\].MUX\[3\]/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_55_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[3\].DIODE_A1MUX\[30\] Do0MUX.M\[3\].MUX\[6\]/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[20\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[3\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[21\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[4\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[22\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[31\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[16\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_48_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[5\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[17\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[26\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[0\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_6_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_6_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[27\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.DIBUF\[18\].cell DIBUF\[18\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DIBUF\[18\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[1\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND0/Y
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_76_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_76_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[10\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_20_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_112_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_92_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_92_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_112_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_25_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[13\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[22\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_6_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_96_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_89_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_41_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_41_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_41_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[23\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_137_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_137_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_137_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[19\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[6\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[2\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[18\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[7\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[19\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[1\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[3\].DIODE\[1\] BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xfill_34_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_142_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_142_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_142_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_142_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_142_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_142_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[2\].DIODE\[6\] BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[2\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/X
+ sky130_fd_sc_hd__and4_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_60_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[28\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_53_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xfill_46_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[11\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_1_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_82_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_127_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[12\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_75_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[3\].DIODE_A2MUX\[28\] Do0MUX.M\[3\].MUX\[4\]/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[21\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_11_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_68_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[24\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_87_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_107_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_107_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_107_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_87_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[22\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_123_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_123_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_123_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[5\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_11_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_36_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_36_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[8\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[17\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_4_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_94_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_52_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_52_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_139_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[18\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_138_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[1\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[30\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[2\].Do_FF\[2\] BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X
+ BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[2\].MUX\[2\]/A3
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[13\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[31\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[1\].Do_FF\[7\] BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X
+ BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[1\].MUX\[7\]/A1
+ sky130_fd_sc_hd__dfxtp_1
Xfill_32_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_25_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[27\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[14\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND3/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell BLOCK\[0\].RAM32.TIE0\[0\].cell/LO
+ BLOCK\[0\].RAM32.FBUFENBUF0\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[10\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[26\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[15\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[27\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[9\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_3_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND0/Y
+ sky130_fd_sc_hd__nor4b_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell BLOCK\[2\].RAM32.TIE0\[3\].cell/LO
+ BLOCK\[2\].RAM32.FBUFENBUF0\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[10\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_73_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF BLOCK\[1\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[3\].Do_FF\[4\] BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X
+ BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[3\].MUX\[4\]/A0
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_132_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_80_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_125_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell BLOCK\[2\].RAM32.WEBUF\[0\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X sky130_fd_sc_hd__clkbuf_2
Xtap_73_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_118_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_98_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_66_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[7\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_118_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_118_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_118_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_98_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_59_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.ABUF\[1\] BLOCK\[2\].RAM32.A0BUF\[1\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B sky130_fd_sc_hd__clkbuf_2
Xtap_134_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_134_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[19\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[28\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_134_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_47_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_47_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[2\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[29\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_63_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[3\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[12\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[30\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[24\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[13\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[25\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[8\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[26\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_23_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[9\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_16_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[1\].DIODE\[2\] BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[21\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_68_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_45_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell BLOCK\[1\].RAM32.WEBUF\[1\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[0\].DIODE\[7\] BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_38_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[4\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_84_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_84_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[22\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[31\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_17_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[18\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_17_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[27\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[5\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_120_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_120_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_33_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[17\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[1\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_130_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[26\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_129_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_123_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[15\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[6\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_129_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_129_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF BLOCK\[2\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND1/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_71_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_116_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_64_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[0\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_122_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xtap_109_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_57_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[27\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_58_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[1\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[10\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell BLOCK\[3\].RAM32.TIE0\[2\].cell/LO
+ BLOCK\[3\].RAM32.FBUFENBUF0\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[7\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[19\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_85_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_78_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[2\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[20\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[7\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_0_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[3\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[21\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[30\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_9_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND4 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND4/X
+ sky130_fd_sc_hd__and4bb_2
XDo0MUX.M\[1\].MUX\[0\] Do0MUX.M\[1\].MUX\[0\]/A0 Do0MUX.M\[1\].MUX\[0\]/A1 Do0MUX.M\[1\].MUX\[0\]/A2
+ Do0MUX.M\[1\].MUX\[0\]/A3 Do0MUX.SEL0BUF\[1\]/X Do0MUX.SEL1BUF\[1\]/X VGND VGND
+ VPWR VPWR Do0[8] sky130_fd_sc_hd__mux4_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[0\].Do_FF\[3\] BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X
+ BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[0\].MUX\[3\]/A2
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[4\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_79_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_102_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_79_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[16\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_50_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_43_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_115_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_115_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_95_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_95_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_36_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_115_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[26\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_28_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[17\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_131_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_131_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_131_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[0\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_44_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.DIBUF\[20\].cell DIBUF\[20\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DIBUF\[20\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_44_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_44_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_104_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xfill_104_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_104_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_104_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_60_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_60_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_121_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[12\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[21\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[2\].Do_FF\[0\] BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X
+ BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[2\].MUX\[0\]/A1
+ sky130_fd_sc_hd__dfxtp_1
Xfill_120_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_113_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XDo0MUX.M\[0\].MUX\[2\] Do0MUX.M\[0\].MUX\[2\]/A0 Do0MUX.M\[0\].MUX\[2\]/A1 Do0MUX.M\[0\].MUX\[2\]/A2
+ Do0MUX.M\[0\].MUX\[2\]/A3 Do0MUX.SEL0BUF\[0\]/X Do0MUX.SEL1BUF\[0\]/X VGND VGND
+ VPWR VPWR Do0[2] sky130_fd_sc_hd__mux4_1
Xfill_106_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[22\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[9\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[18\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[23\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[5\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[8\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[17\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[6\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XEN0BUF.cell EN0 VGND VGND VPWR VPWR DEC0.AND3/C sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[18\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_90_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_83_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.TIE0\[0\].cell VGND VGND VPWR VPWR BLOCK\[1\].RAM32.TIE0\[0\].cell/HI
+ BLOCK\[1\].RAM32.TIE0\[0\].cell/LO sky130_fd_sc_hd__conb_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[1\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_76_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[15\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_8_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_101_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_101_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_81_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[27\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_98_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell BLOCK\[3\].RAM32.WEBUF\[2\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X sky130_fd_sc_hd__clkbuf_2
Xtap_30_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[10\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[28\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[15\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_30_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_100_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_126_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_126_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_126_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_41_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[11\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell BLOCK\[1\].RAM32.TIE0\[0\].cell/LO
+ BLOCK\[1\].RAM32.FBUFENBUF0\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_34_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_55_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[12\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[21\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_55_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_71_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF BLOCK\[0\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[16\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[7\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[17\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[0\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[29\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell BLOCK\[0\].RAM32.TIE0\[2\].cell/LO
+ BLOCK\[0\].RAM32.FBUFENBUF0\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[1\].DIODE\[0\] BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDo0MUX.M\[3\].MUX\[7\] Do0MUX.M\[3\].MUX\[7\]/A0 Do0MUX.M\[3\].MUX\[7\]/A1 Do0MUX.M\[3\].MUX\[7\]/A2
+ Do0MUX.M\[3\].MUX\[7\]/A3 Do0MUX.SEL0BUF\[3\]/X Do0MUX.SEL1BUF\[3\]/X VGND VGND
+ VPWR VPWR Do0[31] sky130_fd_sc_hd__mux4_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[3\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[12\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[30\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_6_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[26\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[13\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[31\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.DIBUF\[6\].cell DIBUF\[6\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DIBUF\[6\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XDo0MUX.M\[1\].DIODE_A2MUX\[13\] Do0MUX.M\[1\].MUX\[5\]/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[9\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_76_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[25\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell BLOCK\[2\].RAM32.WEBUF\[3\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X sky130_fd_sc_hd__clkbuf_2
Xtap_20_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[14\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_13_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_92_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[26\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[8\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_112_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_112_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_92_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_25_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_96_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[9\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_89_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_41_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_41_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_41_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_137_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_137_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_137_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XDo0MUX.M\[0\].DIODE_A3MUX\[2\] Do0MUX.M\[0\].MUX\[2\]/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[23\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_66_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[6\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[2\].DIODE_A2MUX\[17\] Do0MUX.M\[2\].MUX\[1\]/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[18\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[27\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_142_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[7\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_142_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_142_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_142_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND2/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xfill_1_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.DIBUF\[24\].cell DIBUF\[24\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DIBUF\[24\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xfill_142_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_142_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[1\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[28\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[6\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[15\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[2\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[11\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[29\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_60_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[12\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_53_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[0\].Do_FF\[1\] BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X
+ BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[0\].MUX\[1\]/A0
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[24\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_46_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[25\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_75_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[7\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_68_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[8\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_107_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_107_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_87_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_87_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_107_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_123_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_123_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_123_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[20\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_11_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_36_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_36_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_4_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[3\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_94_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_52_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_52_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_52_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[21\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[30\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[3\].Do_FF\[6\] BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X
+ BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[3\].MUX\[6\]/A3
+ sky130_fd_sc_hd__dfxtp_1
Xtap_139_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[17\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_87_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell BLOCK\[1\].RAM32.TIE0\[1\].cell/LO
+ BLOCK\[1\].RAM32.FBUFENBUF0\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[4\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_138_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[31\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell BLOCK\[3\].RAM32.TIE0\[3\].cell/LO
+ BLOCK\[3\].RAM32.FBUFENBUF0\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[16\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[0\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[14\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[5\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[17\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[26\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[0\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[23\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_3_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND1 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND1/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[6\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[9\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[18\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDIBUF\[28\].cell Di0[28] VGND VGND VPWR VPWR DIBUF\[28\].cell/X sky130_fd_sc_hd__clkbuf_16
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[7\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[23\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[19\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF BLOCK\[2\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[6\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_132_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_80_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_22_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_125_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND0/Y
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_73_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_118_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_98_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[2\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[20\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_66_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_118_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_118_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_98_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_59_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_134_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_134_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[3\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_134_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_47_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_47_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_47_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[15\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_63_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_63_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[25\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[16\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_35_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XDo0MUX.SEL1BUF\[3\] DEC0.AND3/A VGND VGND VPWR VPWR Do0MUX.SEL1BUF\[3\]/X sky130_fd_sc_hd__clkbuf_2
Xfill_136_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[28\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[11\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[2\].DIODE\[6\] BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[12\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell BLOCK\[2\].RAM32.TIE0\[0\].cell/LO
+ BLOCK\[2\].RAM32.FBUFENBUF0\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[21\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.TIE0\[3\].cell VGND VGND VPWR VPWR BLOCK\[2\].RAM32.TIE0\[3\].cell/HI
+ BLOCK\[2\].RAM32.TIE0\[3\].cell/LO sky130_fd_sc_hd__conb_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[8\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_16_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[17\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[22\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.DIBUF\[28\].cell DIBUF\[28\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DIBUF\[28\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[16\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[5\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[17\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_38_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.WEBUF\[1\].cell WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.WEBUF\[1\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
Xtap_84_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[0\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_17_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[31\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_120_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_120_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_33_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_130_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_129_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_129_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_129_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[14\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_123_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_71_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_116_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_64_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[26\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_109_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_57_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[15\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[31\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_58_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_58_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[9\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[27\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[14\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_74_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[10\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell BLOCK\[2\].RAM32.WEBUF\[0\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X sky130_fd_sc_hd__clkbuf_2
XDIBUF\[11\].cell Di0[11] VGND VGND VPWR VPWR DIBUF\[11\].cell/X sky130_fd_sc_hd__clkbuf_16
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF BLOCK\[3\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[11\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[20\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell BLOCK\[0\].RAM32.TIE0\[3\].cell/LO
+ BLOCK\[0\].RAM32.FBUFENBUF0\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[23\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.DIBUF\[9\].cell DIBUF\[9\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DIBUF\[9\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[1\].Do_FF\[7\] BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X
+ BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[1\].MUX\[7\]/A2
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_78_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[6\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_0_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[16\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[7\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_9_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND5 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND5/X
+ sky130_fd_sc_hd__and4b_2
Xtap_9_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[28\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_79_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_102_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[2\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_50_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[11\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[29\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_43_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_115_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_95_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_95_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_36_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_115_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_115_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[25\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[3\].Do_FF\[4\] BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X
+ BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[3\].MUX\[4\]/A1
+ sky130_fd_sc_hd__dfxtp_1
Xtap_28_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[12\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[30\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_131_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_131_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_131_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_44_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[8\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[24\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_44_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_44_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[13\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_104_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_104_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_104_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_60_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_60_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_60_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[25\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_121_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_114_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.DIBUF\[11\].cell DIBUF\[11\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DIBUF\[11\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell BLOCK\[1\].RAM32.WEBUF\[1\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_120_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[8\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_113_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_106_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.DIBUF\[16\].cell DIBUF\[16\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DIBUF\[16\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[22\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF BLOCK\[0\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[31\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[5\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[17\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[6\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[31\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[15\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[0\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[18\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_83_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[27\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_76_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[5\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[14\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_69_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[1\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[28\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_101_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_101_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[2\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_98_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[11\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_14_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[1\].DIODE\[2\] BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_30_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[0\].DIODE\[7\] BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_30_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_100_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_126_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_126_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[23\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[24\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_41_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_34_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell BLOCK\[1\].RAM32.TIE0\[2\].cell/LO
+ BLOCK\[1\].RAM32.FBUFENBUF0\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[6\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell BLOCK\[0\].RAM32.WEBUF\[2\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X sky130_fd_sc_hd__clkbuf_2
Xtap_27_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_55_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_55_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_55_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.SEL_DIODE\[1\] DEC0.AND3/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND1/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[7\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_71_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_71_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[19\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[2\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[20\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[2\].DIODE\[4\] BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[16\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[21\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[3\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[30\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[4\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[16\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF BLOCK\[1\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[25\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_6_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.DIBUF\[2\].cell DIBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DIBUF\[2\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_20_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[13\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[22\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_13_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_92_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[0\].Do_FF\[3\] BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X
+ BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[0\].MUX\[3\]/A3
+ sky130_fd_sc_hd__dfxtp_1
Xtap_112_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_112_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_6_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[23\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[8\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_96_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[17\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_89_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_41_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_41_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell BLOCK\[3\].RAM32.TIE0\[0\].cell/LO
+ BLOCK\[3\].RAM32.FBUFENBUF0\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[6\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[22\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_41_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_137_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_137_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_137_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[18\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[5\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_32_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[1\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_66_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[19\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_66_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_82_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[2\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell BLOCK\[3\].RAM32.WEBUF\[2\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[2\].Do_FF\[0\] BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X
+ BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[2\].MUX\[0\]/A2
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_142_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_142_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_142_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_142_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[31\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xfill_1_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xfill_142_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_142_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[1\].Do_FF\[5\] BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X
+ BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[1\].MUX\[5\]/A0
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[14\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XDo0MUX.M\[3\].DIODE_A0MUX\[29\] Do0MUX.M\[3\].MUX\[5\]/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[15\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[27\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_60_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_46_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_39_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[10\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_1_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[24\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[11\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_11_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[20\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_68_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_107_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_107_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_87_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[21\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.DIBUF\[30\].cell DIBUF\[30\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DIBUF\[30\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xtap_123_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_123_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_123_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF BLOCK\[2\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xtap_11_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[4\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_36_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_36_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[16\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_4_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_52_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_52_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_52_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_94_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_139_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_87_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_138_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[30\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell BLOCK\[2\].RAM32.WEBUF\[3\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_77_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[13\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[31\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.Do0_REG.Root_CLKBUF BLOCK\[2\].RAM32.CLKBUF.cell/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.Do0_REG.Root_CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[25\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[14\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[30\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[8\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[26\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[13\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[9\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[27\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[10\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_3_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND2 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND2/X
+ sky130_fd_sc_hd__and4bb_2
Xtap_3_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[1\].DIODE\[0\] BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_51_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[22\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[31\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell BLOCK\[3\].RAM32.TIE0\[3\].cell/LO
+ BLOCK\[3\].RAM32.FBUFENBUF0\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_132_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[5\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_80_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_125_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_73_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_118_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_66_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_118_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_118_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_98_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_98_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[6\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[15\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_59_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_134_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[18\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[27\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_134_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_47_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_47_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_47_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[1\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.ABUF\[1\] BLOCK\[3\].RAM32.A0BUF\[1\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B sky130_fd_sc_hd__clkbuf_2
Xtap_63_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[28\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_63_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_63_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF BLOCK\[3\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xfill_35_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[24\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[2\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_35_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[11\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[29\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_136_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[12\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_129_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[24\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_23_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_16_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.EN0BUF.cell DEC0.AND0/Y VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DEC0.AND3/C
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[21\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[4\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_99_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[22\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[31\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[0\].Do_FF\[1\] BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X
+ BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[0\].MUX\[1\]/A1
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[16\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[5\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[21\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[30\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.DEC0.AND0 BLOCK\[0\].RAM32.DEC0.AND3/B BLOCK\[0\].RAM32.DEC0.AND3/A
+ BLOCK\[0\].RAM32.DEC0.AND3/C VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DEC0.AND0/Y sky130_fd_sc_hd__nor3b_2
Xtap_17_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[17\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_17_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[26\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[4\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_120_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_120_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XWEBUF\[2\].cell WE0[2] VGND VGND VPWR VPWR WEBUF\[2\].cell/X sky130_fd_sc_hd__clkbuf_2
Xtap_33_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[0\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_130_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[27\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_129_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_129_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_129_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_123_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_71_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_116_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[1\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_64_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_109_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[10\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_57_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_58_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_58_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_58_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF BLOCK\[0\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[13\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[22\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_74_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_74_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_90_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[23\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[6\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[18\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[7\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_78_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[1\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[19\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_0_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[20\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[2\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_9_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[29\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_21_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND6 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND6/X
+ sky130_fd_sc_hd__and4b_2
Xtap_9_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_14_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[3\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_50_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_43_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_115_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_95_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_36_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_115_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.TIE0\[3\].cell VGND VGND VPWR VPWR BLOCK\[0\].RAM32.TIE0\[3\].cell/HI
+ BLOCK\[0\].RAM32.TIE0\[3\].cell/LO sky130_fd_sc_hd__conb_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_131_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_131_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND0/Y
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_44_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_44_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_44_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell BLOCK\[0\].RAM32.TIE0\[3\].cell/LO
+ BLOCK\[0\].RAM32.FBUFENBUF0\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[12\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[21\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_104_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_60_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_60_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[24\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_121_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_60_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XDo0MUX.M\[0\].DIODE_A0MUX\[7\] Do0MUX.M\[0\].MUX\[7\]/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_114_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[22\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_62_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_120_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_107_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.A0BUF\[2\].cell A0BUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.A0BUF\[2\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_106_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[5\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[21\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[8\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_85_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[17\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[4\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF BLOCK\[1\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[18\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[1\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[30\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[2\].DIODE\[6\] BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XDo0MUX.M\[1\].DIODE_A3MUX\[9\] Do0MUX.M\[1\].MUX\[1\]/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[13\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[31\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_76_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_69_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[14\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_101_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_101_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_98_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[26\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_14_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[15\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_30_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[9\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[27\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_30_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.DIBUF\[22\].cell DIBUF\[22\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DIBUF\[22\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xtap_100_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_126_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_126_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_41_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[10\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_39_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_55_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_55_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_55_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[20\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[11\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_71_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_71_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_111_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[29\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XDo0MUX.M\[1\].DIODE_A0MUX\[14\] Do0MUX.M\[1\].MUX\[6\]/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[3\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[12\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[30\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[24\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[13\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[29\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell BLOCK\[1\].RAM32.TIE0\[2\].cell/LO
+ BLOCK\[1\].RAM32.FBUFENBUF0\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[1\].Do_FF\[7\] BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X
+ BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[1\].MUX\[7\]/A3
+ sky130_fd_sc_hd__dfxtp_1
Xtap_6_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[25\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[12\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_81_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[8\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[26\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_13_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDIBUF\[3\].cell Di0[3] VGND VGND VPWR VPWR DIBUF\[3\].cell/X sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_112_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_112_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[9\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_6_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.FBUFENBUF0\[3\].cell DEC0.AND0/Y VGND VGND VPWR VPWR BLOCK\[0\].RAM32.FBUFENBUF0\[3\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_96_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_89_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_41_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_41_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[2\].DIODE_A0MUX\[18\] Do0MUX.M\[2\].MUX\[2\]/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[21\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_41_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_137_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_137_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_137_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[3\].Do_FF\[4\] BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X
+ BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[3\].MUX\[4\]/A2
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[4\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[22\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[31\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_32_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_66_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_66_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[0\].DIODE_A1MUX\[1\] Do0MUX.M\[0\].MUX\[1\]/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[5\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_66_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_82_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_82_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[17\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[26\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[6\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_142_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_142_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_142_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[15\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_1_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_142_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_142_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[0\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[27\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[1\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell BLOCK\[0\].RAM32.WEBUF\[2\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[10\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[28\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_60_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[11\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_1_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_11_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_11_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_107_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[20\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_107_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[7\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[3\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_123_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_123_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_11_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_36_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[21\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[30\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_36_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_4_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[0\].DIODE\[7\] BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[4\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_52_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_52_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_52_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[20\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[29\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_94_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_139_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[16\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_87_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[3\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_138_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell BLOCK\[2\].RAM32.TIE0\[1\].cell/LO
+ BLOCK\[2\].RAM32.FBUFENBUF0\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[17\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_77_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_77_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.DIBUF\[26\].cell DIBUF\[26\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DIBUF\[26\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[26\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[0\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_93_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[2\].DIODE_A2MUX\[22\] Do0MUX.M\[2\].MUX\[6\]/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.ABUF\[1\] BLOCK\[0\].RAM32.A0BUF\[1\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[12\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[21\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[2\].DIODE\[4\] BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[22\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_3_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND3 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND3/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[5\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[23\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[8\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[17\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_51_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[6\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_44_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[18\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_80_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_22_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[7\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_125_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_73_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[3\].DIODE_A2MUX\[26\] Do0MUX.M\[3\].MUX\[2\]/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_118_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[19\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[1\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_118_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_118_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_98_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_66_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_59_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_134_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[2\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_134_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_47_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_47_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_47_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_63_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_63_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_63_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_2_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_92_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_35_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_137_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[28\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[15\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_136_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_129_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[11\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_88_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[12\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[2\].Do_FF\[0\] BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X
+ BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[2\].MUX\[0\]/A3
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[21\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[11\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[1\].Do_FF\[5\] BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X
+ BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[1\].MUX\[5\]/A1
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[20\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_23_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[16\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_16_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[17\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell BLOCK\[2\].RAM32.TIE0\[1\].cell/LO
+ BLOCK\[2\].RAM32.FBUFENBUF0\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_99_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[0\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[29\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_17_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.DEC0.AND1 BLOCK\[0\].RAM32.DEC0.AND3/A BLOCK\[0\].RAM32.DEC0.AND3/B
+ BLOCK\[0\].RAM32.DEC0.AND3/C VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DEC0.AND1/X sky130_fd_sc_hd__and3b_2
Xtap_17_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_120_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[3\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[12\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[30\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_120_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[3\].Do_FF\[2\] BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X
+ BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[3\].MUX\[2\]/A0
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_33_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_130_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_129_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_129_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_123_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[13\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_71_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[31\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_116_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_64_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_109_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[25\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_57_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[14\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_58_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_58_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_58_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[8\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[26\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_74_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[15\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_74_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_74_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[9\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_90_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_90_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[19\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[10\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_141_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF BLOCK\[1\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell BLOCK\[1\].RAM32.TIE0\[3\].cell/LO
+ BLOCK\[1\].RAM32.FBUFENBUF0\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[7\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[28\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_21_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/X
+ sky130_fd_sc_hd__and4_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[6\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_9_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_14_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[15\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[2\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[11\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[29\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND0/Y
+ sky130_fd_sc_hd__nor4b_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[1\].DIODE\[0\] BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[12\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[28\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_43_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_36_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_115_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_115_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_28_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[0\].DIODE\[5\] BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[24\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[11\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_28_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_131_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_131_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[25\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_44_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_44_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_44_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_104_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_60_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_60_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[8\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_60_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_121_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_114_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_62_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_120_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xtap_107_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_69_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_55_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_113_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[20\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_106_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_85_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_85_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[3\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[21\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XA0BUF\[3\].cell A0[3] VGND VGND VPWR VPWR A0BUF\[3\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[30\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.ENBUF BLOCK\[3\].RAM32.DEC0.AND3/X VGND VGND
+ VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell BLOCK\[3\].RAM32.CLKBUF.cell/X VGND
+ VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[4\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[31\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[16\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[5\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[14\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[17\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[26\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[15\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_69_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF BLOCK\[2\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[0\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[27\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_101_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[1\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_14_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[10\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[0\].Do_FF\[1\] BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X
+ BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[0\].MUX\[1\]/A2
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_30_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_100_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_126_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_126_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_39_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_41_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[23\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[7\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_55_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.DIBUF\[13\].cell DIBUF\[13\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DIBUF\[13\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xtap_55_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_55_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.DIBUF\[5\].cell DIBUF\[5\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DIBUF\[5\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[19\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell BLOCK\[2\].RAM32.TIE0\[2\].cell/LO
+ BLOCK\[2\].RAM32.FBUFENBUF0\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[6\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_71_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_71_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[0\].DIODE_A2MUX\[6\] Do0MUX.M\[0\].MUX\[6\]/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[2\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[20\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[7\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[3\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[19\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_111_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XDo0MUX.M\[0\].MUX\[0\] Do0MUX.M\[0\].MUX\[0\]/A0 Do0MUX.M\[0\].MUX\[0\]/A1 Do0MUX.M\[0\].MUX\[0\]/A2
+ Do0MUX.M\[0\].MUX\[0\]/A3 Do0MUX.SEL0BUF\[0\]/X Do0MUX.SEL1BUF\[0\]/X VGND VGND
+ VPWR VPWR Do0[0] sky130_fd_sc_hd__mux4_1
Xfill_104_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_96_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[2\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[16\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[25\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND0/Y
+ sky130_fd_sc_hd__nor4b_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[28\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_6_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[11\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_81_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_74_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[12\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[21\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_112_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_112_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_6_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[22\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_96_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_89_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[16\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_41_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[5\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[23\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_41_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_41_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_137_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_137_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[17\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[6\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_32_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_66_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[18\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[0\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_66_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_66_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell BLOCK\[3\].RAM32.TIE0\[1\].cell/LO
+ BLOCK\[3\].RAM32.FBUFENBUF0\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_18_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_82_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_82_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_82_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[1\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_142_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_142_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_142_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_1_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_142_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_70_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[31\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[15\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[27\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDIBUF\[17\].cell Di0[17] VGND VGND VPWR VPWR DIBUF\[17\].cell/X sky130_fd_sc_hd__clkbuf_16
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[14\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_60_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[10\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[15\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[11\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[20\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_1_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDo0MUX.M\[3\].MUX\[5\] Do0MUX.M\[3\].MUX\[5\]/A0 Do0MUX.M\[3\].MUX\[5\]/A1 Do0MUX.M\[3\].MUX\[5\]/A2
+ Do0MUX.M\[3\].MUX\[5\]/A3 Do0MUX.SEL0BUF\[3\]/X Do0MUX.SEL1BUF\[3\]/X VGND VGND
+ VPWR VPWR Do0[29] sky130_fd_sc_hd__mux4_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[10\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[19\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_11_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_11_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.FBUFENBUF0\[2\].cell DEC0.AND1/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.FBUFENBUF0\[2\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_107_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[1\].DIODE_A2MUX\[11\] Do0MUX.M\[1\].MUX\[3\]/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_107_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[16\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF BLOCK\[0\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xtap_123_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_123_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_36_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_36_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[7\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_4_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_52_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_52_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[28\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_94_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_52_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_139_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_87_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_138_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[2\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[11\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[29\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XDo0MUX.M\[0\].DIODE_A3MUX\[0\] Do0MUX.M\[0\].MUX\[0\]/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_77_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_77_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[12\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_77_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[30\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[2\].MUX\[7\] Do0MUX.M\[2\].MUX\[7\]/A0 Do0MUX.M\[2\].MUX\[7\]/A1 Do0MUX.M\[2\].MUX\[7\]/A2
+ Do0MUX.M\[2\].MUX\[7\]/A3 Do0MUX.SEL0BUF\[2\]/X Do0MUX.SEL1BUF\[2\]/X VGND VGND
+ VPWR VPWR Do0[23] sky130_fd_sc_hd__mux4_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[24\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_93_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_93_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[13\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.DIBUF\[17\].cell DIBUF\[17\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DIBUF\[17\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[25\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[14\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[23\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[26\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[8\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[9\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND4 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND4/X
+ sky130_fd_sc_hd__and4bb_2
Xfill_51_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_44_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_37_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[6\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_22_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[15\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_22_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[31\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_73_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[18\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[27\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_118_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_118_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_118_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_66_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[5\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_59_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[14\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[1\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_134_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_134_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[28\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_47_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[15\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_47_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_47_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[2\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[11\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[27\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_63_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_63_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_63_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_92_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.WEBUF\[0\].cell WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.WEBUF\[0\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[1\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[10\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_35_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[3\].Do_FF\[4\] BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X
+ BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[3\].MUX\[4\]/A3
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_137_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_85_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[24\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_136_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_129_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_88_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_88_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF BLOCK\[1\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[7\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[19\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_16_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[2\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[20\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_99_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[3\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[21\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[30\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[4\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[31\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[16\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.DEC0.AND2 BLOCK\[0\].RAM32.DEC0.AND3/B BLOCK\[0\].RAM32.DEC0.AND3/A
+ BLOCK\[0\].RAM32.DEC0.AND3/C VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DEC0.AND2/X sky130_fd_sc_hd__and3b_2
Xtap_17_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[25\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_120_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.DIBUF\[8\].cell DIBUF\[8\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DIBUF\[8\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[14\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[5\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_120_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_130_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[26\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_129_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_129_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_123_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_71_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_116_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_64_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[0\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_109_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[9\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_57_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_58_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_58_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_58_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[0\].DIODE\[7\] BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[23\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_74_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_74_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_74_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell BLOCK\[3\].RAM32.TIE0\[0\].cell/LO
+ BLOCK\[3\].RAM32.FBUFENBUF0\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_0_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_90_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_90_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[22\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[6\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_90_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_141_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDo0MUX.SEL1BUF\[1\] DEC0.AND3/A VGND VGND VPWR VPWR Do0MUX.SEL1BUF\[1\]/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[18\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_134_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_99_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[23\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[5\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[1\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[19\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[6\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF BLOCK\[2\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[2\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[18\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[2\].DIODE\[4\] BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell BLOCK\[2\].RAM32.CLKBUF.cell/X VGND
+ VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[1\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_21_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_9_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_14_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[15\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND1 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND1/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[27\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_36_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_115_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_115_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_28_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[10\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_131_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_131_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_44_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_44_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[11\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[20\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_60_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_60_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_60_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_121_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_114_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell BLOCK\[1\].RAM32.TIE0\[3\].cell/LO
+ BLOCK\[1\].RAM32.FBUFENBUF0\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_62_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[21\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_107_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_55_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_48_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_106_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[4\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[22\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_85_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_85_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_85_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[16\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[5\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[17\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[0\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[31\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[1\].Do_FF\[5\] BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X
+ BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[1\].MUX\[5\]/A2
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[30\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[14\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_69_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[26\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XDo0MUX.M\[1\].DIODE_A1MUX\[8\] Do0MUX.M\[1\].MUX\[0\]/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[13\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_14_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[9\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[27\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[14\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[23\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[10\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[26\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_30_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_100_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_126_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_126_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[9\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_39_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_41_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_34_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF BLOCK\[3\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xtap_27_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[3\].Do_FF\[2\] BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X
+ BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[3\].MUX\[2\]/A1
+ sky130_fd_sc_hd__dfxtp_1
Xtap_1_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.DIBUF\[1\].cell DIBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DIBUF\[1\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xtap_55_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_55_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_55_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_71_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_71_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[6\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[15\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[18\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_112_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[27\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_111_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_96_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_104_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_96_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[1\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[28\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[2\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[11\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[29\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[12\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND1 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND1/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[30\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[24\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[13\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell BLOCK\[2\].RAM32.TIE0\[2\].cell/LO
+ BLOCK\[2\].RAM32.FBUFENBUF0\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_74_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[25\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xfill_67_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_112_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[8\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_25_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_96_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[1\].DIODE\[0\] BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_41_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_89_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_41_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[22\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.WEBUF\[3\].cell WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.WEBUF\[3\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_137_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[31\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[0\].DIODE\[5\] BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF BLOCK\[0\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xtap_137_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[5\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[21\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[30\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_66_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[17\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[26\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_66_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_66_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_25_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[4\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[31\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_18_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[0\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_82_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_82_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_82_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_102_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[27\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[5\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_142_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_142_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[14\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_1_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_142_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[1\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[10\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[26\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_70_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_70_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[0\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[9\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[2\].DIODE\[2\] BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[3\] BLOCK\[0\].RAM32.Do0_REG.Root_CLKBUF/X VGND
+ VGND VPWR VPWR BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[23\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[6\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_1_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[18\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_11_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[7\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_107_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[1\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[19\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_123_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_123_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[2\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_11_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[20\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[29\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_36_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_36_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[0\].Do_FF\[1\] BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X
+ BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[0\].MUX\[1\]/A3
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_4_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[3\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_52_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_52_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_94_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[30\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[2\].DIODE_A0MUX\[23\] Do0MUX.M\[2\].MUX\[7\]/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_139_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_87_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDIBUF\[23\].cell Di0[23] VGND VGND VPWR VPWR DIBUF\[23\].cell/X sky130_fd_sc_hd__clkbuf_16
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_7_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[13\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[4\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[16\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_77_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_77_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[25\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_77_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell BLOCK\[3\].RAM32.TIE0\[1\].cell/LO
+ BLOCK\[3\].RAM32.FBUFENBUF0\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_93_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_93_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_93_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[22\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[1\].Do_FF\[3\] BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X
+ BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[1\].MUX\[3\]/A0
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.ABUF\[1\] BLOCK\[1\].RAM32.A0BUF\[1\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[21\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[5\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[8\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[3\].DIODE_A0MUX\[27\] Do0MUX.M\[3\].MUX\[3\]/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[17\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND5 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND5/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[22\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[4\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.FBUFENBUF0\[1\].cell DEC0.AND2/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.FBUFENBUF0\[1\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
Xfill_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[18\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[5\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_44_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfill_37_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[1\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[17\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_22_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_22_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[0\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_118_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_66_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_118_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_59_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[31\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.DIBUF\[23\].cell DIBUF\[23\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DIBUF\[23\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xtap_134_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_134_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_47_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[14\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_47_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_47_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[26\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_63_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_63_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[15\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_63_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.DIBUF\[28\].cell DIBUF\[28\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DIBUF\[28\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_35_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_35_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell BLOCK\[3\].RAM32.WEBUF\[0\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[9\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_92_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[27\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_137_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_85_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_78_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_136_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_88_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_88_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[10\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_88_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[11\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[20\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[21\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[4\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF BLOCK\[2\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[16\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xfill_99_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[30\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.DEC0.AND3 BLOCK\[0\].RAM32.DEC0.AND3/A BLOCK\[0\].RAM32.DEC0.AND3/B
+ BLOCK\[0\].RAM32.DEC0.AND3/C VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DEC0.AND3/X sky130_fd_sc_hd__and3_2
Xtap_17_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.DIBUF\[4\].cell DIBUF\[4\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DIBUF\[4\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[29\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[13\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_120_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_33_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XDo0MUX.M\[3\].DIODE_A2MUX\[31\] Do0MUX.M\[3\].MUX\[7\]/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_130_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[25\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_129_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_129_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_123_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_71_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[30\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[12\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_116_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_64_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDIBUF\[9\].cell Di0[9] VGND VGND VPWR VPWR DIBUF\[9\].cell/X sky130_fd_sc_hd__clkbuf_16
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[8\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_109_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[26\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_57_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[13\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_58_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_4_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_58_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_58_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[9\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[25\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_74_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_74_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_74_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[8\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_0_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_90_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_90_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_142_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_110_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_90_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_141_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.ENBUF BLOCK\[0\].RAM32.DEC0.AND1/X VGND VGND
+ VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[22\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_99_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_99_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_134_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[31\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_127_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[5\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[17\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[26\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[6\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell BLOCK\[0\].RAM32.TIE0\[1\].cell/LO
+ BLOCK\[0\].RAM32.FBUFENBUF0\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[15\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.A0BUF\[1\].cell A0BUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.A0BUF\[1\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[0\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell BLOCK\[2\].RAM32.TIE0\[3\].cell/LO
+ BLOCK\[2\].RAM32.FBUFENBUF0\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[27\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.DIBUF\[11\].cell DIBUF\[11\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DIBUF\[11\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[1\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[10\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[28\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND2 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND2/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_97_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF BLOCK\[3\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[11\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[29\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_115_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[12\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_131_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_131_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[24\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_44_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_44_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_60_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_60_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_121_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_114_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_62_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_107_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[7\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_55_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_48_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[21\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_106_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_85_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[30\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_105_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_85_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_85_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[4\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[20\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[29\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[16\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[3\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[30\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[17\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[26\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[4\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[13\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[16\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[0\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[25\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[3\].DIODE_A3MUX\[29\] Do0MUX.M\[3\].MUX\[5\]/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_69_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.ABUF\[2\] BLOCK\[0\].RAM32.A0BUF\[2\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_14_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_12_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF BLOCK\[0\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[22\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_30_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[5\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[23\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_126_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_126_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_41_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[8\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[17\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_34_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_27_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[6\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_1_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_55_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_55_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_55_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[18\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[7\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_71_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[1\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_71_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[19\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell BLOCK\[3\].RAM32.TIE0\[2\].cell/LO
+ BLOCK\[3\].RAM32.FBUFENBUF0\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XDo0MUX.M\[0\].DIODE_A0MUX\[5\] Do0MUX.M\[0\].MUX\[5\]/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_112_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_60_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[2\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[20\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_105_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[29\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_96_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_104_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_96_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_96_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[3\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[24\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_105_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[15\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND2 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND2/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[12\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[21\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[2\].DIODE\[4\] BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_74_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_67_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[20\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[11\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.TIE0\[1\].cell VGND VGND VPWR VPWR BLOCK\[3\].RAM32.TIE0\[1\].cell/HI
+ BLOCK\[3\].RAM32.TIE0\[1\].cell/LO sky130_fd_sc_hd__conb_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[16\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_25_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[21\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_96_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[17\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_89_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[4\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_41_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_41_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.DIBUF\[15\].cell DIBUF\[15\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DIBUF\[15\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_137_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_137_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[0\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[16\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF BLOCK\[1\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_32_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_66_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_66_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_66_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[30\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_82_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_82_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[3\].DIODE\[6\] BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_102_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_102_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_82_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_142_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_142_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[13\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[31\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_1_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.ENBUF BLOCK\[1\].RAM32.DEC0.AND0/Y VGND VGND
+ VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[25\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_70_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[14\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_70_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[8\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[26\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[15\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[9\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[1\].DIODE_A0MUX\[12\] Do0MUX.M\[1\].MUX\[4\]/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[10\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[19\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_1_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[20\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[1\].Do_FF\[5\] BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X
+ BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[1\].MUX\[5\]/A3
+ sky130_fd_sc_hd__dfxtp_1
Xtap_11_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[3\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_123_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_11_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_36_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_36_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[6\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[15\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_4_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_52_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[29\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_94_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_52_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_139_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_87_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[2\].DIODE_A0MUX\[16\] Do0MUX.M\[2\].MUX\[0\]/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_7_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_7_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[28\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[12\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[3\].Do_FF\[2\] BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X
+ BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[3\].MUX\[2\]/A2
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[24\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_77_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_77_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_77_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[29\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_30_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[11\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[2\].Do_FF\[7\] BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X
+ BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[2\].MUX\[7\]/A0
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_23_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[25\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_93_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_93_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_93_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[12\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_113_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[8\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[24\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.A0BUF\[4\].cell A0BUF\[4\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DEC0.AND3/A
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell BLOCK\[0\].RAM32.TIE0\[2\].cell/LO
+ BLOCK\[0\].RAM32.FBUFENBUF0\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[21\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND6 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND6/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[30\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_51_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_44_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[4\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_37_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[31\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[16\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[5\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[14\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_22_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_118_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[17\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[26\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_59_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[15\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[0\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_134_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_134_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[27\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_47_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_47_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[1\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[10\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_63_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_63_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[28\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_63_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[0\].DIODE\[5\] BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_35_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_35_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_92_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[11\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_137_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_85_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_78_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_136_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_129_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xtap_88_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_88_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.DIBUF\[19\].cell DIBUF\[19\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DIBUF\[19\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xtap_108_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_88_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell BLOCK\[0\].RAM32.WEBUF\[0\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[23\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[6\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XDo0MUX.M\[2\].DIODE_A2MUX\[20\] Do0MUX.M\[2\].MUX\[4\]/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[20\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[7\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[3\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[2\].DIODE\[2\] BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[19\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.FBUFENBUF0\[0\].cell DEC0.AND3/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.FBUFENBUF0\[0\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF BLOCK\[3\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[2\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[29\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[20\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[16\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[25\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[3\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_17_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[24\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_42_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_33_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_129_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_123_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XDo0MUX.M\[3\].DIODE_A2MUX\[24\] Do0MUX.M\[3\].MUX\[0\]/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_129_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_71_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_116_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_64_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_109_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_57_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[12\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_58_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[21\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_58_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[22\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_74_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_74_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_74_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[16\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_0_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_90_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_142_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_110_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_110_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_90_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_90_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_90_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[5\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[23\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_135_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[17\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_141_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_99_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_99_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_99_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[6\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_134_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_127_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[0\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[18\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[1\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[19\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell BLOCK\[3\].RAM32.WEBUF\[0\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[28\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XDo0MUX.M\[1\].DIODE_A3MUX\[14\] Do0MUX.M\[1\].MUX\[6\]/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[1\].Do_FF\[3\] BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X
+ BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[1\].MUX\[3\]/A1
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF BLOCK\[0\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[2\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[31\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[14\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND3 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND3/X
+ sky130_fd_sc_hd__and4b_2
Xfill_97_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[15\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_28_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[11\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[20\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_131_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_44_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_44_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[3\].Do_FF\[0\] BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X
+ BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[3\].MUX\[0\]/A0
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[19\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[10\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_60_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_60_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell BLOCK\[0\].RAM32.TIE0\[0\].cell/LO
+ BLOCK\[0\].RAM32.FBUFENBUF0\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_121_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[2\].DIODE_A3MUX\[18\] Do0MUX.M\[2\].MUX\[2\]/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_114_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_62_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[20\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_107_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_55_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[16\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[3\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_48_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_106_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_105_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell BLOCK\[2\].RAM32.TIE0\[3\].cell/LO
+ BLOCK\[2\].RAM32.FBUFENBUF0\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_85_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_85_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_85_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_105_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_121_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[29\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell BLOCK\[2\].RAM32.WEBUF\[1\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[12\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[30\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[24\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[13\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_69_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[25\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[14\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[23\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_14_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[8\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[26\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_12_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[9\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_30_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_126_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_41_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[3\] BLOCK\[1\].RAM32.Do0_REG.Root_CLKBUF/X VGND
+ VGND VPWR VPWR BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[19\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[10\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_34_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_27_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[0\].DIODE\[3\] BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_1_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_55_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_55_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[31\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_71_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_71_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF BLOCK\[1\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[5\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[14\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_112_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_60_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[28\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_105_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_53_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_96_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[15\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_116_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_104_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_96_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_96_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell BLOCK\[1\].RAM32.WEBUF\[2\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[2\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[27\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[11\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[1\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[28\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[10\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_105_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_105_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[24\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[11\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND3 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND3/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_67_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell BLOCK\[3\].RAM32.TIE0\[2\].cell/LO
+ BLOCK\[3\].RAM32.FBUFENBUF0\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_25_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[20\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_25_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_8_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_89_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_41_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_41_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[3\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[21\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[30\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_137_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_137_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[4\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[31\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_32_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[16\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[25\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_66_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_66_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[5\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_18_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[14\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_102_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_82_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_82_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_102_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_102_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_82_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[26\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_142_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDo0MUX.M\[0\].DIODE_A2MUX\[4\] Do0MUX.M\[0\].MUX\[4\]/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_1_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[0\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[9\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF BLOCK\[2\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[27\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_70_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_70_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[10\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_102_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[22\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.DIBUF\[21\].cell DIBUF\[21\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DIBUF\[21\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[5\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[23\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_1_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XCLKBUF.cell CLK VGND VGND VPWR VPWR CLKBUF.cell/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[19\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[6\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[2\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[18\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_72_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[7\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[1\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[28\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[19\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_36_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_36_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_52_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[2\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_94_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_52_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_139_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_87_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_7_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_77_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.TIE0\[1\].cell VGND VGND VPWR VPWR BLOCK\[1\].RAM32.TIE0\[1\].cell/HI
+ BLOCK\[1\].RAM32.TIE0\[1\].cell/LO sky130_fd_sc_hd__conb_1
Xtap_77_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_77_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_93_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_93_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[11\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_113_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_113_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_93_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[20\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[21\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell BLOCK\[3\].RAM32.WEBUF\[3\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[4\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[22\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell BLOCK\[1\].RAM32.TIE0\[0\].cell/LO
+ BLOCK\[1\].RAM32.FBUFENBUF0\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[16\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.ABUF\[1\] BLOCK\[2\].RAM32.A0BUF\[1\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[5\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/X
+ sky130_fd_sc_hd__and4_2
Xfill_51_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[17\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_44_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND0/Y
+ sky130_fd_sc_hd__nor4b_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[0\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[18\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[3\].MUX\[3\] Do0MUX.M\[3\].MUX\[3\]/A0 Do0MUX.M\[3\].MUX\[3\]/A1 Do0MUX.M\[3\].MUX\[3\]/A2
+ Do0MUX.M\[3\].MUX\[3\]/A3 Do0MUX.SEL0BUF\[3\]/X Do0MUX.SEL1BUF\[3\]/X VGND VGND
+ VPWR VPWR Do0[27] sky130_fd_sc_hd__mux4_1
Xtap_22_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[1\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[30\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_134_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[13\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_47_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_47_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[27\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_63_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell BLOCK\[0\].RAM32.TIE0\[2\].cell/LO
+ BLOCK\[0\].RAM32.FBUFENBUF0\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_63_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[14\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_2_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[23\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_35_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xtap_92_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[26\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_137_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[10\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_85_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_78_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_136_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_129_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_88_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.DIBUF\[7\].cell DIBUF\[7\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DIBUF\[7\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[9\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_108_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_108_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_88_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_88_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[7\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[3\].DIODE\[6\] BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[10\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[2\].MUX\[5\] Do0MUX.M\[2\].MUX\[5\]/A0 Do0MUX.M\[2\].MUX\[5\]/A1 Do0MUX.M\[2\].MUX\[5\]/A2
+ Do0MUX.M\[2\].MUX\[5\]/A3 Do0MUX.SEL0BUF\[2\]/X Do0MUX.SEL1BUF\[2\]/X VGND VGND
+ VPWR VPWR Do0[21] sky130_fd_sc_hd__mux4_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[19\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_124_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[28\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[2\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[11\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[29\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_17_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_42_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_35_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[12\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[30\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.DIBUF\[25\].cell DIBUF\[25\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DIBUF\[25\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xtap_33_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[1\].MUX\[7\] Do0MUX.M\[1\].MUX\[7\]/A0 Do0MUX.M\[1\].MUX\[7\]/A1 Do0MUX.M\[1\].MUX\[7\]/A2
+ Do0MUX.M\[1\].MUX\[7\]/A3 Do0MUX.SEL0BUF\[1\]/X Do0MUX.SEL1BUF\[1\]/X VGND VGND
+ VPWR VPWR Do0[15] sky130_fd_sc_hd__mux4_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[24\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_129_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[13\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_71_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_116_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_64_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_109_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[25\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_57_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_58_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_58_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[8\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_74_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_74_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[18\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[9\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_90_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_142_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_110_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_110_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_110_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_90_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_90_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[3\].Do_FF\[2\] BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X
+ BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[3\].MUX\[2\]/A3
+ sky130_fd_sc_hd__dfxtp_1
Xtap_90_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_135_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_83_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xfill_141_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_128_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_99_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_99_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[21\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xtap_119_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_99_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[30\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[2\].Do_FF\[7\] BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X
+ BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[2\].MUX\[7\]/A1
+ sky130_fd_sc_hd__dfxtp_1
Xfill_127_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[4\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[31\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[27\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND0/Y
+ sky130_fd_sc_hd__nor4b_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[5\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[14\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[1\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[26\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[10\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell BLOCK\[1\].RAM32.TIE0\[1\].cell/LO
+ BLOCK\[1\].RAM32.FBUFENBUF0\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[15\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell BLOCK\[0\].RAM32.WEBUF\[0\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[0\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[27\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[9\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell BLOCK\[3\].RAM32.TIE0\[3\].cell/LO
+ BLOCK\[3\].RAM32.FBUFENBUF0\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND4 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND4/X
+ sky130_fd_sc_hd__and4bb_2
Xfill_97_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[10\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_28_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF BLOCK\[1\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xtap_44_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_44_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[7\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_60_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_60_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_121_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[19\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_114_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_62_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_107_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_55_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.DEC0.AND0 BLOCK\[3\].RAM32.DEC0.AND3/B BLOCK\[3\].RAM32.DEC0.AND3/A
+ BLOCK\[3\].RAM32.DEC0.AND3/C VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DEC0.AND0/Y sky130_fd_sc_hd__nor3b_2
Xtap_48_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[2\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_106_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[20\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_105_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_105_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[29\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_85_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_85_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_85_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[7\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[0\].DIODE\[5\] BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[3\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDIBUF\[29\].cell Di0[29] VGND VGND VPWR VPWR DIBUF\[29\].cell/X sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[30\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_121_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_121_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[4\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[13\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.DIBUF\[0\].cell DIBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DIBUF\[0\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[16\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[25\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_132_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[26\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_69_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[0\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[9\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[2\].DIODE\[2\] BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_12_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[1\].DIODE\[7\] BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[21\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.ABUF\[2\] BLOCK\[1\].RAM32.A0BUF\[2\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_30_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[4\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[22\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_34_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[18\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_1_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[23\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_27_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[5\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_55_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_55_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[1\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell BLOCK\[2\].RAM32.TIE0\[0\].cell/LO
+ BLOCK\[2\].RAM32.FBUFENBUF0\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[17\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[6\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_71_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_71_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[0\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF BLOCK\[2\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[0\].RAM32.DIBUF\[29\].cell DIBUF\[29\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DIBUF\[29\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[18\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_112_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_60_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[1\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_105_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_53_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_20_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_46_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_116_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_116_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_104_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_96_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_96_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_96_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.WEBUF\[2\].cell WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.WEBUF\[2\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[15\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_132_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[27\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_105_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_105_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[10\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND4 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND4/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[11\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[20\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[7\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[1\].Do_FF\[3\] BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X
+ BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[1\].MUX\[3\]/A2
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[21\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDIBUF\[12\].cell Di0[12] VGND VGND VPWR VPWR DIBUF\[12\].cell/X sky130_fd_sc_hd__clkbuf_16
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell BLOCK\[2\].RAM32.WEBUF\[1\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X sky130_fd_sc_hd__clkbuf_2
Xtap_25_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[4\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_8_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[16\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_41_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_41_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_137_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[17\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell BLOCK\[0\].RAM32.TIE0\[3\].cell/LO
+ BLOCK\[0\].RAM32.FBUFENBUF0\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_32_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_66_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_66_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[0\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[3\].Do_FF\[0\] BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X
+ BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[3\].MUX\[0\]/A1
+ sky130_fd_sc_hd__dfxtp_1
Xtap_18_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[29\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_82_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_102_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_102_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_102_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_82_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[12\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[30\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_15_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[26\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_70_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_70_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[13\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_110_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[9\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_127_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[25\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[14\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_102_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[23\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[8\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[9\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[18\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_1_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF BLOCK\[3\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.DIBUF\[12\].cell DIBUF\[12\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DIBUF\[12\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell BLOCK\[1\].RAM32.WEBUF\[2\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[6\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[15\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_72_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.DIBUF\[17\].cell DIBUF\[17\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DIBUF\[17\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xfill_65_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_36_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_36_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[27\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[1\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[10\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_94_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[28\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_52_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_52_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_139_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[15\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_87_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_7_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_7_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[11\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[0\].DIODE\[3\] BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[29\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_77_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_77_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_77_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[12\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_30_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_113_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_93_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_93_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[24\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_16_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_113_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_113_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_93_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_9_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[25\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[7\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[8\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[2\].DIODE\[0\] BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell BLOCK\[1\].RAM32.TIE0\[2\].cell/LO
+ BLOCK\[1\].RAM32.FBUFENBUF0\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[20\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell BLOCK\[0\].RAM32.WEBUF\[3\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[29\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[1\] BLOCK\[0\].RAM32.Do0_REG.Root_CLKBUF/X VGND
+ VGND VPWR VPWR BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF BLOCK\[0\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xfill_44_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[3\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND1 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND1/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[30\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[17\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[26\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[4\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[31\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[13\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[0\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[25\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[16\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[14\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[26\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_47_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_47_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[9\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[0\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_63_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_63_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_92_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XDo0MUX.M\[2\].DIODE_A0MUX\[21\] Do0MUX.M\[2\].MUX\[5\]/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_137_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_85_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_78_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[23\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.DIBUF\[3\].cell DIBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DIBUF\[3\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_88_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_108_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_108_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_108_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_88_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_88_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[6\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_124_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[18\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_124_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[23\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[7\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_140_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[1\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[19\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[6\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[2\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell BLOCK\[3\].RAM32.TIE0\[0\].cell/LO
+ BLOCK\[3\].RAM32.FBUFENBUF0\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[20\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[29\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[1\].Do_FF\[1\] BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X
+ BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[1\].MUX\[1\]/A0
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[3\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[3\].DIODE_A0MUX\[25\] Do0MUX.M\[3\].MUX\[1\]/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[24\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[15\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_42_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[25\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_35_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell BLOCK\[3\].RAM32.WEBUF\[3\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_28_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[8\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.A0BUF\[0\].cell A0BUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.A0BUF\[0\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
Xtap_64_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_109_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_57_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[11\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_4_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[20\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_58_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_58_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_4_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_74_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_74_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[21\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[17\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_0_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_110_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_110_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_90_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_90_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[22\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[4\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_142_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_110_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_90_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[1\].DIODE_A1MUX\[15\] Do0MUX.M\[1\].MUX\[7\]/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_135_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[0\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_83_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[16\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_141_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_128_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_99_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_99_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_76_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[5\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_134_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_119_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_119_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_99_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[3\] BLOCK\[2\].RAM32.Do0_REG.Root_CLKBUF/X VGND
+ VGND VPWR VPWR BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[17\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_135_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[0\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.DIBUF\[31\].cell DIBUF\[31\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DIBUF\[31\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND1 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND1/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[31\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[14\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_140_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[26\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND5 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND5/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[15\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[9\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XDo0MUX.M\[2\].DIODE_A1MUX\[19\] Do0MUX.M\[2\].MUX\[3\]/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[14\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[23\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_28_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[10\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[19\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_44_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_44_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[20\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_60_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_60_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_121_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_114_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[3\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_62_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_107_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_55_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.DEC0.AND1 BLOCK\[3\].RAM32.DEC0.AND3/A BLOCK\[3\].RAM32.DEC0.AND3/B
+ BLOCK\[3\].RAM32.DEC0.AND3/C VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DEC0.AND1/X sky130_fd_sc_hd__and3b_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_48_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_106_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[6\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_105_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_85_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_85_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[15\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_105_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF BLOCK\[2\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xtap_85_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[16\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_18_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell BLOCK\[3\].RAM32.TIE0\[3\].cell/LO
+ BLOCK\[3\].RAM32.FBUFENBUF0\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_121_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_121_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_121_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_140_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[28\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[3\].DIODE\[6\] BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_132_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[11\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[29\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_125_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[25\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[12\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_69_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[8\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[24\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[13\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[22\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.CLKBUF.cell CLKBUF.cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.CLKBUF.cell/X
+ sky130_fd_sc_hd__clkbuf_4
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[25\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[8\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_95_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_1_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[31\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_55_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_55_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell BLOCK\[3\].RAM32.CLKBUF.cell/X VGND
+ VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[5\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[14\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_71_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_71_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[17\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[26\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[2\].DIODE_A3MUX\[23\] Do0MUX.M\[2\].MUX\[7\]/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[15\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[31\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_112_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_60_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[0\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_105_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[27\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_53_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[14\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_116_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_116_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_96_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_96_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_96_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.EN0BUF.cell DEC0.AND1/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DEC0.AND3/C
+ sky130_fd_sc_hd__clkbuf_2
Xtap_46_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_116_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_104_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[1\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_39_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[10\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[28\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_132_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_132_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[11\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF BLOCK\[3\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xfill_105_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_105_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[2\].Do_FF\[7\] BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X
+ BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[2\].MUX\[7\]/A2
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XWEBUF\[3\].cell WE0[3] VGND VGND VPWR VPWR WEBUF\[3\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND5 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND5/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[23\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[24\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[6\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XDo0MUX.M\[3\].DIODE_A3MUX\[27\] Do0MUX.M\[3\].MUX\[3\]/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_67_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[7\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[19\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.ABUF\[0\] BLOCK\[0\].RAM32.A0BUF\[0\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_10_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_8_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_41_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[2\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[20\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[29\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[16\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[25\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[3\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[30\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_32_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_66_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_66_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[24\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[4\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_18_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[13\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_82_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_102_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_102_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_102_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_82_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[25\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_15_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[8\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_70_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_70_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_31_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[0\].DIODE_A0MUX\[3\] Do0MUX.M\[0\].MUX\[3\]/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_110_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_127_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_127_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_103_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_102_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[22\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF BLOCK\[0\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[5\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[23\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[17\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[22\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_1_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[6\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[0\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[18\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[5\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.A0BUF\[3\].cell A0BUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DEC0.AND3/B
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[1\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[19\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[2\].DIODE\[2\] BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[28\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_72_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_65_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[1\].DIODE\[7\] BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[2\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_58_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_36_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[31\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_52_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_52_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_94_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_139_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[14\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_87_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_7_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[24\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[15\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_77_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_77_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_30_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_93_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_113_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_113_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_113_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_93_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_93_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[10\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[19\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_26_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[3\].DIODE\[4\] BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_9_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[20\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_138_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[16\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.DIBUF\[23\].cell DIBUF\[23\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DIBUF\[23\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[21\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[3\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[4\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XDo0MUX.M\[1\].DIODE_A0MUX\[10\] Do0MUX.M\[1\].MUX\[2\]/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[16\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF BLOCK\[1\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.ABUF\[1\] BLOCK\[3\].RAM32.A0BUF\[1\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND2 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND2/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[30\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[1\].Do_FF\[3\] BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X
+ BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[1\].MUX\[3\]/A3
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[13\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[25\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_47_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_47_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[14\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[23\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[8\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[26\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_63_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_63_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[13\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_2_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[22\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_35_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[9\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_92_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_137_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_85_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell BLOCK\[1\].RAM32.TIE0\[2\].cell/LO
+ BLOCK\[1\].RAM32.FBUFENBUF0\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_12_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_78_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_12_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[10\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_108_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_108_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_108_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[3\].Do_FF\[0\] BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X
+ BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[3\].MUX\[0\]/A2
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_88_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_88_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[19\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_124_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[2\].Do_FF\[5\] BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X
+ BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[2\].MUX\[5\]/A0
+ sky130_fd_sc_hd__dfxtp_1
Xtap_124_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_124_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDIBUF\[4\].cell Di0[4] VGND VGND VPWR VPWR DIBUF\[4\].cell/X sky130_fd_sc_hd__clkbuf_16
Xtap_21_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[31\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_140_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[5\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[14\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[15\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[27\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[1\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[10\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[28\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND6/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xfill_42_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[24\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_35_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[29\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[11\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_28_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[12\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell BLOCK\[0\].RAM32.WEBUF\[3\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X sky130_fd_sc_hd__clkbuf_2
Xtap_57_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[24\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_4_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_58_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_58_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_74_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_74_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_0_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[21\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_110_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_110_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[0\].DIODE\[3\] BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_90_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_90_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_142_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[30\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_110_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_90_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_135_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_83_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_141_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_128_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_99_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_76_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[4\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_119_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_119_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_119_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_99_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_99_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_69_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[31\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[16\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_135_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[25\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[5\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_135_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[14\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[30\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[26\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[4\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND2 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND2/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[13\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[0\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[9\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[27\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[2\].DIODE\[0\] BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_140_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_140_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[10\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND6 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND6/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell BLOCK\[2\].RAM32.TIE0\[1\].cell/LO
+ BLOCK\[2\].RAM32.FBUFENBUF0\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.DIBUF\[27\].cell DIBUF\[27\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DIBUF\[27\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[22\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[5\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_40_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[23\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_44_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[6\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_60_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_60_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_121_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[18\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_114_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_62_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_107_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[7\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_55_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.DEC0.AND2 BLOCK\[3\].RAM32.DEC0.AND3/B BLOCK\[3\].RAM32.DEC0.AND3/A
+ BLOCK\[3\].RAM32.DEC0.AND3/C VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DEC0.AND2/X sky130_fd_sc_hd__and3b_2
Xtap_48_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_106_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[1\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[19\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_105_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_85_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_85_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[28\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_105_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell BLOCK\[2\].RAM32.CLKBUF.cell/X VGND
+ VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_18_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF BLOCK\[3\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[2\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_18_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[29\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_121_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_121_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_121_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_140_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[3\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[12\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_133_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[24\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xfill_132_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_125_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_118_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_69_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XDo0MUX.M\[1\].DIODE_A3MUX\[12\] Do0MUX.M\[1\].MUX\[4\]/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[21\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[1\].Do_FF\[1\] BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X
+ BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[1\].MUX\[1\]/A1
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[4\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[22\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[16\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_95_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[21\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[5\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.ABUF\[2\] BLOCK\[2\].RAM32.A0BUF\[2\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C sky130_fd_sc_hd__clkbuf_2
Xfill_88_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_39_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[17\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[4\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_55_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[0\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[18\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_55_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_71_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_71_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[1\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[30\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[2\].DIODE_A3MUX\[16\] Do0MUX.M\[2\].MUX\[0\]/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_112_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_60_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_105_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_53_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF BLOCK\[0\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xtap_116_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_116_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[13\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_96_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_96_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_46_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_116_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_104_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.DIBUF\[10\].cell DIBUF\[10\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DIBUF\[10\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xtap_29_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[14\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_132_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_132_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_132_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[23\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[26\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_105_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_105_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND6 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND6/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[9\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[7\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[10\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[19\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_67_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[20\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[3\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_8_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[29\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[1\] BLOCK\[1\].RAM32.Do0_REG.Root_CLKBUF/X VGND
+ VGND VPWR VPWR BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X sky130_fd_sc_hd__clkbuf_4
Xtap_32_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell BLOCK\[1\].RAM32.TIE0\[3\].cell/LO
+ BLOCK\[1\].RAM32.FBUFENBUF0\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_66_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_66_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[0\].DIODE\[1\] BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_25_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[12\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[30\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_18_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[24\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_102_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_102_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_82_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_82_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_102_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[29\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_15_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[13\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[25\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_31_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_70_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_70_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[12\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_31_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_110_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_127_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_127_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_103_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[8\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_51_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_127_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_102_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[9\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[18\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[3\].DIODE\[6\] BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[21\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[30\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[4\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[31\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF BLOCK\[1\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[5\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[14\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_65_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_58_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[26\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XA0BUF\[4\].cell A0[4] VGND VGND VPWR VPWR A0BUF\[4\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[15\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[0\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[9\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_52_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[27\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.ABUF\[1\] BLOCK\[0\].RAM32.A0BUF\[1\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B sky130_fd_sc_hd__clkbuf_2
Xfill_6_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_87_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_7_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[28\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[10\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_77_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_77_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[11\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_30_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_23_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_93_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_113_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_113_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_113_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_93_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_26_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_9_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XDo0MUX.M\[0\].DIODE_A2MUX\[2\] Do0MUX.M\[0\].MUX\[2\]/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_99_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_42_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_138_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_138_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[20\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[29\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[7\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_100_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND5/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[3\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[30\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[2\].Do_FF\[7\] BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X
+ BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[2\].MUX\[7\]/A3
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[1\].RAM32.DIBUF\[14\].cell DIBUF\[14\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DIBUF\[14\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.DIBUF\[6\].cell DIBUF\[6\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DIBUF\[6\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell BLOCK\[2\].RAM32.TIE0\[2\].cell/LO
+ BLOCK\[2\].RAM32.FBUFENBUF0\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[4\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[13\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[29\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND3 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND3/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[16\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[25\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[3\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[12\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[26\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[3\] BLOCK\[3\].RAM32.Do0_REG.Root_CLKBUF/X VGND
+ VGND VPWR VPWR BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_70_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[0\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[9\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_47_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF BLOCK\[2\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_63_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_63_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[21\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_92_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_137_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[4\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_85_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_12_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[22\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_78_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_108_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_108_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_88_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_88_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_108_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[5\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[23\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_124_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[17\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_124_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_124_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_21_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[6\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_14_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_37_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_140_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_140_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[0\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[18\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[7\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[19\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[1\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[28\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[2\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell BLOCK\[3\].RAM32.TIE0\[1\].cell/LO
+ BLOCK\[3\].RAM32.FBUFENBUF0\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_42_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_35_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_28_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XDo0MUX.M\[3\].MUX\[1\] Do0MUX.M\[3\].MUX\[1\]/A0 Do0MUX.M\[3\].MUX\[1\]/A1 Do0MUX.M\[3\].MUX\[1\]/A2
+ Do0MUX.M\[3\].MUX\[1\]/A3 Do0MUX.SEL0BUF\[3\]/X Do0MUX.SEL1BUF\[3\]/X VGND VGND
+ VPWR VPWR Do0[25] sky130_fd_sc_hd__mux4_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[11\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[20\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[7\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[1\].DIODE\[7\] BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_4_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDIBUF\[18\].cell Di0[18] VGND VGND VPWR VPWR DIBUF\[18\].cell/X sky130_fd_sc_hd__clkbuf_16
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[21\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_58_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_58_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_74_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[20\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[4\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_74_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[16\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_0_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_110_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_90_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_90_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[3\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_142_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_110_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_110_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_90_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_23_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_135_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_83_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[17\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_23_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_141_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_128_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_99_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_76_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_119_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_119_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_119_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_99_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_99_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_69_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.FBUFENBUF0\[3\].cell DEC0.AND1/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.FBUFENBUF0\[3\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF BLOCK\[3\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[0\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell BLOCK\[0\].RAM32.TIE0\[0\].cell/LO
+ BLOCK\[0\].RAM32.FBUFENBUF0\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_135_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell BLOCK\[1\].RAM32.CLKBUF.cell/X VGND
+ VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_135_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_135_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[29\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[3\].DIODE\[4\] BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDo0MUX.M\[2\].MUX\[3\] Do0MUX.M\[2\].MUX\[3\]/A0 Do0MUX.M\[2\].MUX\[3\]/A1 Do0MUX.M\[2\].MUX\[3\]/A2
+ Do0MUX.M\[2\].MUX\[3\]/A3 Do0MUX.SEL0BUF\[2\]/X Do0MUX.SEL1BUF\[2\]/X VGND VGND
+ VPWR VPWR Do0[19] sky130_fd_sc_hd__mux4_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND3 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND3/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XDo0MUX.SEL0BUF\[3\] DEC0.AND3/B VGND VGND VPWR VPWR Do0MUX.SEL0BUF\[3\]/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[12\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[30\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[13\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_140_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_140_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[25\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[14\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[23\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/X
+ sky130_fd_sc_hd__and4_2
XDo0MUX.M\[3\].DIODE_A0MUX\[30\] Do0MUX.M\[3\].MUX\[6\]/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[8\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[9\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[18\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.DIBUF\[18\].cell DIBUF\[18\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DIBUF\[18\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[7\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_40_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[19\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[1\].MUX\[5\] Do0MUX.M\[1\].MUX\[5\]/A0 Do0MUX.M\[1\].MUX\[5\]/A1 Do0MUX.M\[1\].MUX\[5\]/A2
+ Do0MUX.M\[1\].MUX\[5\]/A3 Do0MUX.SEL0BUF\[1\]/X Do0MUX.SEL1BUF\[1\]/X VGND VGND
+ VPWR VPWR Do0[13] sky130_fd_sc_hd__mux4_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_60_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[2\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_114_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_62_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_107_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_55_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.DEC0.AND3 BLOCK\[3\].RAM32.DEC0.AND3/A BLOCK\[3\].RAM32.DEC0.AND3/B
+ BLOCK\[3\].RAM32.DEC0.AND3/C VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DEC0.AND3/X sky130_fd_sc_hd__and3_2
Xtap_48_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_85_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_105_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_105_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_85_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[28\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_121_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_121_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[15\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_121_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_140_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[11\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[29\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[3\].Do_FF\[0\] BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X
+ BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[3\].MUX\[0\]/A3
+ sky130_fd_sc_hd__dfxtp_1
Xtap_133_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_81_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_126_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_50_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[2\].Do_FF\[5\] BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X
+ BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[2\].MUX\[5\]/A1
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[28\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_125_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[12\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_118_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[24\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[0\].MUX\[7\] Do0MUX.M\[0\].MUX\[7\]/A0 Do0MUX.M\[0\].MUX\[7\]/A1 Do0MUX.M\[0\].MUX\[7\]/A2
+ Do0MUX.M\[0\].MUX\[7\]/A3 Do0MUX.SEL0BUF\[0\]/X Do0MUX.SEL1BUF\[0\]/X VGND VGND
+ VPWR VPWR Do0[7] sky130_fd_sc_hd__mux4_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[11\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_69_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[25\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[8\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.WEBUF\[1\].cell WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.WEBUF\[1\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND6/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[20\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[29\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_95_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_88_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[3\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[30\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_1_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_55_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[4\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[13\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[31\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_71_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_71_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[16\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[25\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[14\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_112_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_20_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_60_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[26\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_20_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_105_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_53_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_116_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_96_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_96_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[15\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_46_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_116_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_116_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_104_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[0\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_29_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[27\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_29_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[9\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[0\].DIODE\[3\] BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_132_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_132_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_132_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[10\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_45_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[3\].DIODE_A1MUX\[28\] Do0MUX.M\[3\].MUX\[4\]/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.DIBUF\[9\].cell DIBUF\[9\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DIBUF\[9\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xfill_105_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_105_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/X
+ sky130_fd_sc_hd__and4_2
Xfill_130_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF BLOCK\[1\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND0/Y
+ sky130_fd_sc_hd__nor4b_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[7\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[23\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[19\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[6\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[2\].DIODE\[0\] BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[2\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[20\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[29\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_8_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[7\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[1\].DIODE\[5\] BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[3\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.ABUF\[0\] BLOCK\[1\].RAM32.A0BUF\[0\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[19\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[28\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[24\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[2\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_32_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_66_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_66_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[25\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_25_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_18_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_102_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_102_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_82_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_82_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[8\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_15_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_31_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[11\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_70_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_31_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_110_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[20\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_127_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_127_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_103_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_51_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[0\].DIODE_A3MUX\[7\] Do0MUX.M\[0\].MUX\[7\]/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_127_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[21\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND4/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_44_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_102_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[4\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[22\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[16\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[5\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[23\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[17\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[6\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND0/Y
+ sky130_fd_sc_hd__nor4b_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[18\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[0\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[27\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[1\].Do_FF\[1\] BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X
+ BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[1\].MUX\[1\]/A2
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF BLOCK\[2\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_58_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[1\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[0\].Do_FF\[6\] BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X
+ BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[0\].MUX\[6\]/A0
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_6_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[15\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_7_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[14\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[23\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_77_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_77_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[10\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[19\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_30_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_23_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_16_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_113_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_113_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_113_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_93_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_93_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[20\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_26_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[7\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_9_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_99_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[19\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_42_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[3\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_42_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_138_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_138_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_138_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[2\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[16\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_100_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.DIBUF\[2\].cell DIBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DIBUF\[2\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.ENBUF BLOCK\[1\].RAM32.DEC0.AND3/X VGND VGND
+ VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[28\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND4 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND4/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[11\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[29\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[12\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[24\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_70_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_63_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[13\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[22\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[25\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_63_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[23\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[8\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_35_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_92_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_137_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_85_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[6\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_78_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[0\].DIODE\[1\] BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[9\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.DIBUF\[20\].cell DIBUF\[20\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DIBUF\[20\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xtap_108_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_108_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_88_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_88_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[18\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_108_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell BLOCK\[2\].RAM32.TIE0\[2\].cell/LO
+ BLOCK\[2\].RAM32.FBUFENBUF0\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_124_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_124_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_124_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_37_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_37_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_140_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_140_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_53_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[15\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[31\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[27\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[14\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[1\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[10\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[28\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[15\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[27\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[11\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_42_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[10\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_35_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[24\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_4_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_58_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[7\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[19\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_74_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_74_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_110_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[2\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_90_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_90_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[20\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_142_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_110_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_90_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[29\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_23_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_135_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_83_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_141_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_128_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_119_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_119_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_99_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_99_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[3\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_76_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[30\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_119_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_69_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_135_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[24\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[4\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_135_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_135_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[13\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[31\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_48_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[25\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND4 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND4/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[14\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[26\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[8\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDIBUF\[24\].cell Di0[24] VGND VGND VPWR VPWR DIBUF\[24\].cell/X sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_140_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_140_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[9\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND5/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[23\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell BLOCK\[3\].RAM32.TIE0\[1\].cell/LO
+ BLOCK\[3\].RAM32.FBUFENBUF0\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_40_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[6\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_33_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[22\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[18\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xfill_26_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[23\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[5\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[1\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[19\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[28\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_62_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_107_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_55_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[6\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_48_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[2\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[18\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_85_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[27\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_105_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_105_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_85_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_18_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.FBUFENBUF0\[2\].cell DEC0.AND2/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.FBUFENBUF0\[2\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[1\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_18_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_121_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_121_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_121_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[24\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_140_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[1\].DIODE_A1MUX\[13\] Do0MUX.M\[1\].MUX\[5\]/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_133_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[15\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_81_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_126_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_74_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_50_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_50_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_119_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.DIBUF\[24\].cell DIBUF\[24\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DIBUF\[24\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xfill_118_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[1\] BLOCK\[2\].RAM32.Do0_REG.Root_CLKBUF/X VGND
+ VGND VPWR VPWR BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[10\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[19\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.ENBUF BLOCK\[2\].RAM32.DEC0.AND2/X VGND VGND
+ VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[20\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.DIBUF\[29\].cell DIBUF\[29\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DIBUF\[29\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell BLOCK\[3\].RAM32.WEBUF\[1\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[3\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[21\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[4\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[31\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[22\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_88_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XDo0MUX.M\[2\].DIODE_A1MUX\[17\] Do0MUX.M\[2\].MUX\[1\]/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[16\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[5\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_1_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.ABUF\[2\] BLOCK\[3\].RAM32.A0BUF\[2\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[17\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_71_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[0\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[1\].DIODE\[7\] BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_112_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_60_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_105_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_53_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[14\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_116_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_96_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_96_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND3/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_46_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[23\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_116_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_116_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_104_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_29_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[26\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_29_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[13\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_132_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_132_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[22\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_132_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.DIBUF\[5\].cell DIBUF\[5\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DIBUF\[5\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_45_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_45_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[9\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_105_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_105_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[23\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[10\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_61_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[19\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[3\].DIODE\[4\] BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[6\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_130_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[9\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_123_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[18\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND1 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND1/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[15\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF BLOCK\[2\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XDo0MUX.M\[1\].DIODE_A2MUX\[9\] Do0MUX.M\[1\].MUX\[1\]/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[27\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_93_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[1\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[10\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[28\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_66_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_25_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[11\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[29\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_18_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell BLOCK\[0\].RAM32.TIE0\[1\].cell/LO
+ BLOCK\[0\].RAM32.FBUFENBUF0\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.A0BUF\[2\].cell A0BUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.A0BUF\[2\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
Xtap_102_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_82_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_82_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell BLOCK\[2\].RAM32.TIE0\[3\].cell/LO
+ BLOCK\[2\].RAM32.FBUFENBUF0\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_102_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.DIBUF\[12\].cell DIBUF\[12\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DIBUF\[12\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[12\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_15_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[24\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_31_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[2\].DIODE_A3MUX\[21\] Do0MUX.M\[2\].MUX\[5\]/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_70_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_31_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[13\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_110_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[22\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_127_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_103_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_127_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_127_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_51_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_44_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xfill_102_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xtap_37_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[8\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_56_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[17\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[2\].Do_FF\[5\] BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X
+ BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[2\].MUX\[5\]/A2
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[31\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[5\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[14\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND1 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND1/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[30\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[26\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[31\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[13\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[4\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[3\].DIODE_A3MUX\[25\] Do0MUX.M\[3\].MUX\[1\]/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[0\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_58_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[9\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[27\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[14\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[26\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND6/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[10\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_6_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_7_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[9\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.ABUF\[1\] BLOCK\[1\].RAM32.A0BUF\[1\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF BLOCK\[3\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xtap_77_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_77_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_23_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[23\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_113_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_113_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_93_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_93_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_113_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[6\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_9_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_99_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_42_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_42_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[18\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_42_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[7\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_138_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_138_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XDo0MUX.M\[0\].DIODE_A0MUX\[1\] Do0MUX.M\[0\].MUX\[1\]/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_138_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[1\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[19\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_101_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[28\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.ENBUF BLOCK\[3\].RAM32.DEC0.AND1/X VGND VGND
+ VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D sky130_fd_sc_hd__clkbuf_2
Xfill_100_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[2\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[29\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[3\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[12\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[30\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND5 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND5/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[24\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell BLOCK\[3\].RAM32.TIE0\[2\].cell/LO
+ BLOCK\[3\].RAM32.FBUFENBUF0\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[13\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[25\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[2\].DIODE\[0\] BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[8\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_70_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_63_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[1\].DIODE\[5\] BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_56_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[22\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_92_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF BLOCK\[0\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xtap_137_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_85_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[21\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[5\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_78_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_12_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[17\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_108_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_88_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_88_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_108_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[22\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[4\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[31\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.TIE0\[2\].cell VGND VGND VPWR VPWR BLOCK\[3\].RAM32.TIE0\[2\].cell/HI
+ BLOCK\[3\].RAM32.TIE0\[2\].cell/LO sky130_fd_sc_hd__conb_1
Xtap_124_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_124_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_124_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[0\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[18\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_21_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_37_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[5\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_37_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_37_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_140_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[1\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[17\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[3\].DIODE\[2\] BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_140_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_53_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_53_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[0\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.DIBUF\[16\].cell DIBUF\[16\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DIBUF\[16\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND4/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[14\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[23\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[26\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[9\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_35_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[7\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[10\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[19\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[1\].Do_FF\[1\] BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X
+ BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[1\].MUX\[1\]/A3
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[0\].Do_FF\[6\] BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X
+ BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[0\].MUX\[6\]/A1
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[20\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_4_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_74_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[3\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[21\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_0_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_90_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[4\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_110_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_110_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_90_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_90_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_135_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[16\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_23_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_83_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_141_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_128_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_119_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_119_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_99_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_99_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_76_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_119_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_69_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF BLOCK\[1\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_135_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_135_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_135_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[30\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_48_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_48_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[2\].Do_FF\[3\] BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X
+ BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[2\].MUX\[3\]/A0
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND5 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND5/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[13\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_64_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[29\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[25\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[12\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_140_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_140_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[8\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[22\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[13\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[9\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[18\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[8\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[17\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_40_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell BLOCK\[1\].RAM32.WEBUF\[0\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_26_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_19_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[31\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell BLOCK\[0\].RAM32.TIE0\[2\].cell/LO
+ BLOCK\[0\].RAM32.FBUFENBUF0\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[5\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_55_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND2/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[14\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_48_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[26\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_105_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_105_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[15\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_85_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_85_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDIBUF\[30\].cell Di0[30] VGND VGND VPWR VPWR DIBUF\[30\].cell/X sky130_fd_sc_hd__clkbuf_16
Xtap_18_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[0\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[9\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_121_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[27\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_121_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_121_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.ABUF\[2\] BLOCK\[0\].RAM32.A0BUF\[2\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[0\].DIODE\[1\] BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_140_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[10\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[28\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_133_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_81_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_50_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_126_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_74_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_50_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_50_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_119_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_67_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[11\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xfill_118_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_59_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[12\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[21\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[24\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF BLOCK\[2\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[7\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell BLOCK\[0\].RAM32.WEBUF\[1\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X sky130_fd_sc_hd__clkbuf_2
Xfill_95_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[30\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[4\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[13\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_1_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[29\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[16\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[25\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[30\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[12\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[3\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.FBUFENBUF0\[1\].cell DEC0.AND3/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.FBUFENBUF0\[1\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[26\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.DIBUF\[30\].cell DIBUF\[30\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DIBUF\[30\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[13\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_112_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[0\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_60_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[25\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_20_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_105_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[9\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_53_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_96_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_46_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_116_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_116_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xfill_104_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_96_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_29_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[8\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_29_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_132_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_132_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_132_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_45_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_45_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_45_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_105_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfill_105_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[22\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_61_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_61_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_131_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[5\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[23\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_130_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_123_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_116_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[17\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND2 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND2/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[6\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[0\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[18\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[7\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XDo0MUX.M\[1\].DIODE_A3MUX\[10\] Do0MUX.M\[1\].MUX\[2\]/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[1\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[19\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[28\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND5/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[2\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF BLOCK\[3\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[29\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_93_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[3\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.ABUF\[0\] BLOCK\[2\].RAM32.A0BUF\[0\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A sky130_fd_sc_hd__clkbuf_2
Xfill_86_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[12\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[24\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell BLOCK\[3\].RAM32.WEBUF\[1\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_18_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_102_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_82_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_102_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[7\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_70_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[21\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_110_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_127_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_127_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_127_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_103_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_51_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[20\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_44_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[4\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_102_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_37_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[0\].DIODE_A1MUX\[6\] Do0MUX.M\[0\].MUX\[6\]/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[16\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_56_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_56_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[21\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[3\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[17\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_72_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[4\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell BLOCK\[0\].RAM32.TIE0\[0\].cell/LO
+ BLOCK\[0\].RAM32.FBUFENBUF0\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[0\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[16\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND2 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND2/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[30\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_69_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_58_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[13\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF BLOCK\[0\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[25\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell BLOCK\[2\].RAM32.WEBUF\[2\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[14\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[23\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_7_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[8\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_77_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[9\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[18\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_30_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[7\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_23_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_113_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_113_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_93_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_93_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_16_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[19\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_26_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_9_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_99_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_42_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[2\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[20\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_42_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_42_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND3/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_138_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_138_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_138_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[3\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_101_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xtap_67_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[15\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND6 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND6/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[3\].DIODE\[4\] BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[29\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[12\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[28\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[24\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[11\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell BLOCK\[1\].RAM32.WEBUF\[3\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[25\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_70_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_63_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[21\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[12\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_56_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[8\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_49_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[24\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_4_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_85_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_78_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_108_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_88_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_88_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_108_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[30\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_124_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_124_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_21_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[4\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_14_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_37_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_37_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_37_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell BLOCK\[3\].RAM32.TIE0\[2\].cell/LO
+ BLOCK\[3\].RAM32.FBUFENBUF0\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[13\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[31\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_140_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[16\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_140_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[25\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_53_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_53_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[14\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF BLOCK\[1\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xtap_53_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_97_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[0\].DIODE_A2MUX\[0\] Do0MUX.M\[0\].MUX\[0\]/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[26\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[15\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[0\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[9\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[27\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[2\].Do_FF\[5\] BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X
+ BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[2\].MUX\[5\]/A3
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[10\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[28\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[11\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_35_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[23\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND1/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[1\] BLOCK\[3\].RAM32.Do0_REG.Root_CLKBUF/X VGND
+ VGND VPWR VPWR BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_4_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[6\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[20\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND6/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[29\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.DIBUF\[22\].cell DIBUF\[22\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DIBUF\[22\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[7\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_0_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_90_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[19\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[3\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_110_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_110_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[3\].Do_FF\[7\] BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X
+ BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[3\].MUX\[7\]/A0
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[28\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_90_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_135_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_83_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_128_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[24\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_119_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_99_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_99_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_76_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[29\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[2\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_119_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_119_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_69_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[25\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[3\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_135_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_135_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_135_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[12\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_48_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_48_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_48_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[24\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND6 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND6/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[8\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_12_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_64_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_64_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xfill_36_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_80_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_140_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_140_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[21\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.TIE0\[2\].cell VGND VGND VPWR VPWR BLOCK\[1\].RAM32.TIE0\[2\].cell/HI
+ BLOCK\[1\].RAM32.TIE0\[2\].cell/LO sky130_fd_sc_hd__conb_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[4\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[22\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[16\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[5\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[23\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[17\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_26_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[6\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_19_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[0\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[18\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[27\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.WEBUF\[0\].cell WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.WEBUF\[0\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[1\].DIODE\[5\] BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell BLOCK\[1\].RAM32.TIE0\[0\].cell/LO
+ BLOCK\[1\].RAM32.FBUFENBUF0\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[1\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_48_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[28\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_105_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_105_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_85_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_18_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[2\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_121_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[11\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_121_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_140_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_133_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_81_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[14\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_126_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_74_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[23\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_50_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_50_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_50_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_119_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_67_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_59_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_59_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[3\].DIODE\[2\] BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDo0MUX.M\[2\].MUX\[1\] Do0MUX.M\[2\].MUX\[1\]/A0 Do0MUX.M\[2\].MUX\[1\]/A1 Do0MUX.M\[2\].MUX\[1\]/A2
+ Do0MUX.M\[2\].MUX\[1\]/A3 Do0MUX.SEL0BUF\[2\]/X Do0MUX.SEL1BUF\[2\]/X VGND VGND
+ VPWR VPWR Do0[17] sky130_fd_sc_hd__mux4_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[20\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_75_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[7\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.SEL0BUF\[1\] DEC0.AND3/B VGND VGND VPWR VPWR Do0MUX.SEL0BUF\[1\]/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[19\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[3\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND4/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[20\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[2\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.DIBUF\[8\].cell DIBUF\[8\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DIBUF\[8\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[16\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_95_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[3\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_1_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF BLOCK\[3\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xfill_31_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[29\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XDo0MUX.M\[1\].MUX\[3\] Do0MUX.M\[1\].MUX\[3\]/A0 Do0MUX.M\[1\].MUX\[3\]/A1 Do0MUX.M\[1\].MUX\[3\]/A2
+ Do0MUX.M\[1\].MUX\[3\]/A3 Do0MUX.SEL0BUF\[1\]/X Do0MUX.SEL1BUF\[1\]/X VGND VGND
+ VPWR VPWR Do0[11] sky130_fd_sc_hd__mux4_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[12\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[0\].Do_FF\[6\] BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X
+ BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[0\].MUX\[6\]/A2
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_112_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_60_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_20_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[24\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_105_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_53_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_96_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[13\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_46_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_116_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_116_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_96_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[22\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_29_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[25\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_29_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_132_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[23\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell BLOCK\[1\].RAM32.WEBUF\[0\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X sky130_fd_sc_hd__clkbuf_2
Xtap_132_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_45_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_45_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[8\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_45_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_105_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.DIBUF\[26\].cell DIBUF\[26\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DIBUF\[26\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xtap_61_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[6\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_61_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_61_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[9\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_131_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[18\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_124_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_130_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[2\].Do_FF\[3\] BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X
+ BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[2\].MUX\[3\]/A1
+ sky130_fd_sc_hd__dfxtp_1
Xfill_123_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_116_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND3 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND3/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[19\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[0\].MUX\[5\] Do0MUX.M\[0\].MUX\[5\]/A0 Do0MUX.M\[0\].MUX\[5\]/A1 Do0MUX.M\[0\].MUX\[5\]/A2
+ Do0MUX.M\[0\].MUX\[5\]/A3 Do0MUX.SEL0BUF\[0\]/X Do0MUX.SEL1BUF\[0\]/X VGND VGND
+ VPWR VPWR Do0[5] sky130_fd_sc_hd__mux4_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_109_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[2\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell BLOCK\[3\].RAM32.CLKBUF.cell/X VGND
+ VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[31\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[14\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDEC0.AND0 DEC0.AND3/B DEC0.AND3/A DEC0.AND3/C VGND VGND VPWR VPWR DEC0.AND0/Y sky130_fd_sc_hd__nor3b_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[28\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.Do0_REG.Root_CLKBUF BLOCK\[1\].RAM32.CLKBUF.cell/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.Do0_REG.Root_CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[15\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_93_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[2\].DIODE_A1MUX\[22\] Do0MUX.M\[2\].MUX\[6\]/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDo0MUX.M\[1\].DIODE_A0MUX\[8\] Do0MUX.M\[1\].MUX\[0\]/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[11\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_86_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[27\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_79_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[28\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[10\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_102_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[24\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_102_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_15_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[11\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_15_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell BLOCK\[1\].RAM32.TIE0\[1\].cell/LO
+ BLOCK\[1\].RAM32.FBUFENBUF0\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell BLOCK\[0\].RAM32.WEBUF\[1\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND2/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell BLOCK\[3\].RAM32.TIE0\[3\].cell/LO
+ BLOCK\[3\].RAM32.FBUFENBUF0\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_31_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_70_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_110_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_127_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_127_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_127_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_103_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_51_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_44_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_37_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[0\].DIODE\[1\] BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_56_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_56_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_56_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[20\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[29\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XDo0MUX.M\[3\].DIODE_A1MUX\[26\] Do0MUX.M\[3\].MUX\[2\]/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_72_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_72_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[3\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[30\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[24\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[4\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[13\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[31\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND3 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND3/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[25\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_69_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[14\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xfill_69_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[8\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_58_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[26\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[9\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.DIBUF\[1\].cell DIBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DIBUF\[1\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[27\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[1\].DIODE\[3\] BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_7_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[10\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_30_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[22\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.ABUF\[1\] BLOCK\[2\].RAM32.A0BUF\[1\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B sky130_fd_sc_hd__clkbuf_2
Xtap_23_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_113_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_93_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_16_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_113_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF BLOCK\[1\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xtap_26_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[5\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[23\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_26_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_9_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_42_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[19\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_99_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_42_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_42_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[28\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[6\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_138_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_138_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_138_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[18\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[2\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_101_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[7\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[27\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[0\].DIODE_A3MUX\[5\] Do0MUX.M\[0\].MUX\[5\]/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_42_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_67_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_67_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[28\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[1\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell BLOCK\[2\].RAM32.TIE0\[0\].cell/LO
+ BLOCK\[2\].RAM32.FBUFENBUF0\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[24\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[2\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_83_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[11\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/X
+ sky130_fd_sc_hd__and4_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND0/Y
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XDo0MUX.M\[3\].DIODE_A3MUX\[30\] Do0MUX.M\[3\].MUX\[6\]/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.WEBUF\[3\].cell WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.WEBUF\[3\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
Xfill_70_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND5/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[20\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_56_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[0\].Do_FF\[4\] BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X
+ BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[0\].MUX\[4\]/A0
+ sky130_fd_sc_hd__dfxtp_1
Xfill_49_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[3\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[21\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_4_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[4\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_78_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[22\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_12_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[31\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_88_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[16\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_108_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_108_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[5\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_124_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_124_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[17\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_21_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_37_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_37_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_37_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell BLOCK\[2\].RAM32.WEBUF\[2\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X sky130_fd_sc_hd__clkbuf_2
XDIBUF\[13\].cell Di0[13] VGND VGND VPWR VPWR DIBUF\[13\].cell/X sky130_fd_sc_hd__clkbuf_16
Xtap_14_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[0\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[18\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_140_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_140_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_53_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[27\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_53_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_53_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_97_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF BLOCK\[2\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[1\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell BLOCK\[0\].RAM32.TIE0\[3\].cell/LO
+ BLOCK\[0\].RAM32.FBUFENBUF0\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_78_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[13\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[22\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[23\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_35_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[10\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[19\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[6\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[18\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[9\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[7\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_4_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[19\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_61_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[2\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_110_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_110_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_90_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_23_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_135_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_83_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell BLOCK\[1\].RAM32.WEBUF\[3\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.DIBUF\[13\].cell DIBUF\[13\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DIBUF\[13\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xtap_128_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_119_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_99_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_99_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_76_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[28\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_119_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_69_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_135_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_135_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_135_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[11\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[29\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_48_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_48_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_48_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.DIBUF\[18\].cell DIBUF\[18\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DIBUF\[18\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/B BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/X
+ sky130_fd_sc_hd__and4_2
Xtap_12_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[12\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_64_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_64_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND3/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_64_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[24\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_5_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_36_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_36_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND0/Y
+ sky130_fd_sc_hd__nor4b_2
Xtap_80_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_80_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[13\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[22\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_140_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_140_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_139_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[8\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[17\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[18\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_33_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[1\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[30\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[4\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[13\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[31\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell BLOCK\[1\].RAM32.TIE0\[2\].cell/LO
+ BLOCK\[1\].RAM32.FBUFENBUF0\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[27\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_105_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_105_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[14\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_18_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[10\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[26\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_121_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_121_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[15\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_140_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[27\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[9\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_133_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_81_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_126_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_50_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_50_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_50_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_74_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.ABUF\[2\] BLOCK\[1\].RAM32.A0BUF\[2\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C sky130_fd_sc_hd__clkbuf_2
Xtap_119_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_67_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[10\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_59_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_59_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_59_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_75_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_75_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND0/Y
+ sky130_fd_sc_hd__nor4b_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[7\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_91_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[19\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[28\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.DIBUF\[4\].cell DIBUF\[4\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DIBUF\[4\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[2\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[29\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[7\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell BLOCK\[2\].RAM32.CLKBUF.cell/X VGND
+ VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[3\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[12\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[30\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_1_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[24\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_31_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[13\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND1/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_24_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell BLOCK\[3\].RAM32.TIE0\[0\].cell/LO
+ BLOCK\[3\].RAM32.FBUFENBUF0\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[25\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_60_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_105_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[8\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_53_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[26\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_116_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_116_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_96_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_46_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[9\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_29_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_132_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[3\].Do_FF\[7\] BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X
+ BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[3\].MUX\[7\]/A1
+ sky130_fd_sc_hd__dfxtp_1
Xtap_132_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_45_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_45_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_45_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_105_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[21\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_61_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_61_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_61_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[1\].DIODE_A1MUX\[11\] Do0MUX.M\[1\].MUX\[3\]/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_131_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.A0BUF\[1\].cell A0BUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.A0BUF\[1\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
Xtap_124_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[4\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_72_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[22\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_130_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_117_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[31\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[18\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_116_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND4 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND4/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[5\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xfill_109_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_86_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[17\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[1\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[6\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[15\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[27\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[18\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[0\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDEC0.AND1 DEC0.AND3/A DEC0.AND3/B DEC0.AND3/C VGND VGND VPWR VPWR DEC0.AND1/X sky130_fd_sc_hd__and3b_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[1\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_86_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_79_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF BLOCK\[1\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.ABUF\[0\] BLOCK\[3\].RAM32.A0BUF\[0\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[7\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_102_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_102_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_15_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[10\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_15_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[19\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[1\].DIODE\[5\] BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_31_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[20\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_110_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[7\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_127_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_127_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_103_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_51_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_44_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[3\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[21\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_37_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_56_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_56_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_56_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[4\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_72_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_72_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_72_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[16\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[17\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[3\].DIODE\[2\] BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[26\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND4 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND4/X
+ sky130_fd_sc_hd__and4bb_2
Xfill_121_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[0\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[2\].DIODE\[7\] BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND4/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[29\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_69_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_69_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_69_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_58_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[12\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[13\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_7_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[22\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_7_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[9\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[18\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[23\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_91_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[17\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[8\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[6\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_23_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_113_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_113_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[18\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_26_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[0\].Do_FF\[6\] BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X
+ BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[0\].MUX\[6\]/A3
+ sky130_fd_sc_hd__dfxtp_1
Xtap_9_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_99_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[1\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_42_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_42_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_42_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_138_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_138_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_101_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.CLKBUF.cell CLKBUF.cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.CLKBUF.cell/X
+ sky130_fd_sc_hd__clkbuf_4
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[15\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_42_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_67_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_67_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_67_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_35_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[27\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF BLOCK\[2\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_83_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[10\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_83_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[28\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[15\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[2\].Do_FF\[3\] BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X
+ BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[2\].MUX\[3\]/A2
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[11\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[12\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[21\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_70_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[24\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_49_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.EN0BUF.cell DEC0.AND2/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DEC0.AND3/C
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[7\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_4_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[8\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[17\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_12_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_108_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_108_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[29\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_124_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_124_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[3\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_21_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_37_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_37_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[12\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[30\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_14_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_37_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND2/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_140_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_140_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_53_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[26\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_53_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_53_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[31\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[13\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_97_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[0\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[9\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[25\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[14\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[26\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[8\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_78_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_78_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_94_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[9\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF BLOCK\[3\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xfill_35_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[23\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[6\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_4_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[18\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[7\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xfill_61_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[1\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[19\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[1\].DIODE\[3\] BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_54_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[28\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[6\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[15\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_110_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_110_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[2\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[29\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_90_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_135_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_83_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_128_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_99_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_76_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[3\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_119_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_119_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_69_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[12\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.A0BUF\[4\].cell A0BUF\[4\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DEC0.AND3/A
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[24\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_135_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_135_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_48_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_48_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_48_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_12_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[25\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_64_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_64_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_64_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[3\].DIODE\[0\] BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[7\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_5_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[8\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_36_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_36_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND1 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND1/X
+ sky130_fd_sc_hd__and4bb_2
Xtap_80_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_80_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_80_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_140_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_139_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_89_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[20\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[3\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[21\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF BLOCK\[0\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[17\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[22\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[4\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[31\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_33_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND0/Y
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[16\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[0\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[5\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.DIBUF\[24\].cell DIBUF\[24\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DIBUF\[24\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[26\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[17\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell BLOCK\[1\].RAM32.CLKBUF.cell/X VGND
+ VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[0\].Do_FF\[4\] BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X
+ BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[0\].MUX\[4\]/A1
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[0\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_105_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_105_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[14\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_121_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_121_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[23\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_140_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_133_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_81_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_50_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_50_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_126_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_74_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_50_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[9\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_119_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_67_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[18\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_59_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[7\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_59_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_59_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[23\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[19\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[2\].Do_FF\[1\] BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X
+ BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[2\].MUX\[1\]/A0
+ sky130_fd_sc_hd__dfxtp_1
Xtap_75_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_75_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[6\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_75_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[2\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[20\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_91_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_91_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND1 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND1/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[3\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.DIBUF\[0\].cell DIBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DIBUF\[0\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[15\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[16\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDIBUF\[5\].cell Di0[5] VGND VGND VPWR VPWR DIBUF\[5\].cell/X sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[28\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_31_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_24_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_17_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[11\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_20_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[25\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_20_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_53_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[12\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_116_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_116_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[21\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_46_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[24\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[8\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[22\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_132_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_132_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_45_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_45_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_45_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_105_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.ABUF\[0\] BLOCK\[0\].RAM32.A0BUF\[0\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[5\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_61_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_61_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_61_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[8\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell BLOCK\[0\].RAM32.TIE0\[1\].cell/LO
+ BLOCK\[0\].RAM32.FBUFENBUF0\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_131_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[17\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_124_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_72_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_130_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xtap_117_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_65_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND5 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND5/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND3/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[31\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_86_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_86_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[14\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[26\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[15\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[31\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XDEC0.AND2 DEC0.AND3/B DEC0.AND3/A DEC0.AND3/C VGND VGND VPWR VPWR DEC0.AND2/X sky130_fd_sc_hd__and3b_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[0\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[9\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[27\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[14\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_93_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[10\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_86_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[28\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_79_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[11\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_102_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_15_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[23\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_31_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_110_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell BLOCK\[2\].RAM32.TIE0\[1\].cell/LO
+ BLOCK\[2\].RAM32.FBUFENBUF0\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_127_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_127_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[6\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_103_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.DIBUF\[28\].cell DIBUF\[28\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DIBUF\[28\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xtap_51_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[16\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_44_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF BLOCK\[2\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xtap_37_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[7\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_56_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_56_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_56_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[19\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[28\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_72_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_72_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_72_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[2\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[29\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[25\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[3\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[30\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND5 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND5/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[12\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_121_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_114_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_97_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[8\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[24\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_69_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_69_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[13\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_69_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_69_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[25\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[8\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_7_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[22\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_91_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_84_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[5\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[23\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND1/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_16_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_113_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_113_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[17\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[22\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_26_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.ABUF\[1\] BLOCK\[3\].RAM32.A0BUF\[1\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[6\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_9_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[31\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.DEC0.AND0 BLOCK\[1\].RAM32.DEC0.AND3/B BLOCK\[1\].RAM32.DEC0.AND3/A
+ BLOCK\[1\].RAM32.DEC0.AND3/C VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DEC0.AND0/Y sky130_fd_sc_hd__nor3b_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[0\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_99_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[18\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_42_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_42_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[27\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[5\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND6/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_138_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_138_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[1\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[28\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[3\].Do_FF\[7\] BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X
+ BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[3\].MUX\[7\]/A2
+ sky130_fd_sc_hd__dfxtp_1
Xtap_101_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_42_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_67_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_67_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_67_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[2\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_35_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[11\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_28_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[0\].DIODE_A1MUX\[4\] Do0MUX.M\[0\].MUX\[4\]/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF BLOCK\[3\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_83_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[3\].DIODE_A1MUX\[31\] Do0MUX.M\[3\].MUX\[7\]/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_83_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_83_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[14\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[23\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[24\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xfill_71_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[7\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.DIBUF\[11\].cell DIBUF\[11\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DIBUF\[11\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_70_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[19\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_56_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[2\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[20\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[16\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_12_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[21\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[3\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[30\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_108_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_108_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[4\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_124_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[16\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_124_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_37_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_37_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_14_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_37_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_140_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_140_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_53_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_53_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_53_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_97_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[13\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[22\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[25\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_78_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_78_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_78_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF BLOCK\[0\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[23\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell BLOCK\[1\].RAM32.TIE0\[3\].cell/LO
+ BLOCK\[1\].RAM32.FBUFENBUF0\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[8\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_94_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_94_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[6\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[22\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_35_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[3\].DIODE\[2\] BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[9\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[18\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[5\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[2\].DIODE\[7\] BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[19\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[2\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[31\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_61_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_54_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[14\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_47_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_110_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_2_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[15\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_83_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell BLOCK\[0\].RAM32.CLKBUF.cell/X VGND
+ VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X sky130_fd_sc_hd__clkbuf_2
Xtap_128_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_76_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[3\].DIODE_A2MUX\[29\] Do0MUX.M\[3\].MUX\[5\]/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_119_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_119_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.A0BUF\[0\].cell A0BUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.A0BUF\[0\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[27\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_69_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_135_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_135_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[10\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[28\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_48_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_48_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_48_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[24\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_12_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XA0BUF\[5\].cell A0[5] VGND VGND VPWR VPWR DEC0.AND3/B sky130_fd_sc_hd__clkbuf_2
Xtap_64_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[11\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_64_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_64_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_5_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_36_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_36_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND2 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND2/X
+ sky130_fd_sc_hd__and4bb_2
Xtap_95_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_80_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_80_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_80_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[21\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[12\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_100_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_140_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_139_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_89_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_89_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[16\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[2\].Do_FF\[3\] BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X
+ BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[2\].MUX\[3\]/A3
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[30\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[4\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[13\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[31\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[25\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[14\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[30\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF BLOCK\[1\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[8\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_105_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[26\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[13\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.DIBUF\[15\].cell DIBUF\[15\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DIBUF\[15\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.DIBUF\[7\].cell DIBUF\[7\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DIBUF\[7\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xtap_18_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell BLOCK\[2\].RAM32.TIE0\[2\].cell/LO
+ BLOCK\[2\].RAM32.FBUFENBUF0\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[9\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[27\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_121_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_121_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_140_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[3\].Do_FF\[5\] BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X
+ BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[3\].MUX\[5\]/A0
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[10\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_133_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_81_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_50_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_50_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_126_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_74_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_119_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_67_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_5_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[22\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_59_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_59_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_59_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND2/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.ABUF\[2\] BLOCK\[2\].RAM32.A0BUF\[2\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_75_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_75_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[5\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[23\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_75_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.DIBUF\[30\].cell DIBUF\[30\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DIBUF\[30\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_91_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_91_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_91_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[6\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND2 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND2/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[18\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[27\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[7\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[1\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[28\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[24\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[2\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[29\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[11\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[12\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_24_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[24\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_17_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_20_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_20_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[1\].DIODE\[3\] BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_116_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_46_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_116_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_132_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_132_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[21\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_45_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_45_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_45_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[4\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[22\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[31\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_61_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_61_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_61_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_131_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_124_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[16\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[21\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[5\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_72_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[30\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_130_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xtap_117_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_65_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDIBUF\[19\].cell Di0[19] VGND VGND VPWR VPWR DIBUF\[19\].cell/X sky130_fd_sc_hd__clkbuf_16
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[17\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_58_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND6 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND6/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[4\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_86_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_86_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_86_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[3\].DIODE\[0\] BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[0\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[18\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[27\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[1\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XDEC0.AND3 DEC0.AND3/A DEC0.AND3/B DEC0.AND3/C VGND VGND VPWR VPWR DEC0.AND3/X sky130_fd_sc_hd__and3_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[13\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[22\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_93_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell BLOCK\[0\].RAM32.TIE0\[0\].cell/LO
+ BLOCK\[0\].RAM32.FBUFENBUF0\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_86_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[23\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND0/Y
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[6\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[9\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_15_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[18\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[1\].MUX\[1\] Do0MUX.M\[1\].MUX\[1\]/A0 Do0MUX.M\[1\].MUX\[1\]/A1 Do0MUX.M\[1\].MUX\[1\]/A2
+ Do0MUX.M\[1\].MUX\[1\]/A3 Do0MUX.SEL0BUF\[1\]/X Do0MUX.SEL1BUF\[1\]/X VGND VGND
+ VPWR VPWR Do0[9] sky130_fd_sc_hd__mux4_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[7\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND5/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[0\].Do_FF\[4\] BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X
+ BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[0\].MUX\[4\]/A2
+ sky130_fd_sc_hd__dfxtp_1
Xtap_31_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[19\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_110_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_127_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_127_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_103_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_51_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_44_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[20\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[2\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_37_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_56_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_56_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_56_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.DIBUF\[19\].cell DIBUF\[19\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DIBUF\[19\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[3\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_72_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_72_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_72_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_122_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[2\].Do_FF\[1\] BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X
+ BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[2\].MUX\[1\]/A1
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF BLOCK\[3\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[29\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_121_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND6 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND6/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_97_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_97_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_114_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XDo0MUX.M\[0\].MUX\[3\] Do0MUX.M\[0\].MUX\[3\]/A0 Do0MUX.M\[0\].MUX\[3\]/A1 Do0MUX.M\[0\].MUX\[3\]/A2
+ Do0MUX.M\[0\].MUX\[3\]/A3 Do0MUX.SEL0BUF\[0\]/X Do0MUX.SEL1BUF\[0\]/X VGND VGND
+ VPWR VPWR Do0[3] sky130_fd_sc_hd__mux4_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[12\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_107_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_69_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_69_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_69_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xfill_69_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_69_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[24\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[13\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[22\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[12\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[21\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[8\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[17\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_91_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDo0MUX.M\[2\].DIODE_A1MUX\[20\] Do0MUX.M\[2\].MUX\[4\]/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_84_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_77_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[18\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_113_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[1\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_26_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_26_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.WEBUF\[2\].cell WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.WEBUF\[2\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
Xtap_9_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[30\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.DEC0.AND1 BLOCK\[1\].RAM32.DEC0.AND3/A BLOCK\[1\].RAM32.DEC0.AND3/B
+ BLOCK\[1\].RAM32.DEC0.AND3/C VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DEC0.AND1/X sky130_fd_sc_hd__and3b_2
Xtap_99_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_42_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_42_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[4\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[13\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[31\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_138_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_138_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF BLOCK\[0\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xtap_101_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[14\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_42_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_67_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_67_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_35_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[26\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_67_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[15\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_83_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_103_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_83_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_83_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[9\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[3\].DIODE_A1MUX\[24\] Do0MUX.M\[3\].MUX\[0\]/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[27\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[10\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_71_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_71_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[20\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[11\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xfill_70_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[1\].DIODE\[1\] BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_12_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[29\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_12_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[7\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_108_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[3\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XDo0MUX.M\[1\].DIODE_A2MUX\[14\] Do0MUX.M\[1\].MUX\[6\]/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[12\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[30\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_124_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_124_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[24\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_21_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_37_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[13\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[29\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_14_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_37_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_37_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_140_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_140_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[25\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_53_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_53_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_53_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[12\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_97_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[8\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[26\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_8_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XDo0MUX.M\[0\].DIODE_A3MUX\[3\] Do0MUX.M\[0\].MUX\[3\]/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_78_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_78_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_78_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[9\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_40_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_94_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_94_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_94_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[21\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XDo0MUX.M\[2\].DIODE_A2MUX\[18\] Do0MUX.M\[2\].MUX\[2\]/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[4\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[22\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[31\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[5\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF BLOCK\[1\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[17\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[6\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[15\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[0\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[18\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_54_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[0\].Do_FF\[2\] BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X
+ BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[0\].MUX\[2\]/A0
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[27\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_47_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[1\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[28\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_2_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_76_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[2\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_119_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_119_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[11\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_69_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_135_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND1/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_135_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_48_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_48_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell BLOCK\[1\].RAM32.TIE0\[0\].cell/LO
+ BLOCK\[1\].RAM32.FBUFENBUF0\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_64_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_64_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_64_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND6/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_5_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xfill_36_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND3 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND3/X
+ sky130_fd_sc_hd__and4b_2
Xtap_95_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_80_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_80_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[3\].Do_FF\[7\] BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X
+ BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[3\].MUX\[7\]/A3
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[20\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_100_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_100_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_80_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[7\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_140_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_88_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_89_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_139_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[3\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[21\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_89_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_89_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[20\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[4\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[16\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[3\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[17\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[26\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[0\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[29\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF BLOCK\[2\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xfill_139_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.DIBUF\[3\].cell DIBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DIBUF\[3\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[12\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_18_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_121_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell BLOCK\[2\].RAM32.WEBUF\[0\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[13\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[22\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_140_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_133_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_81_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_50_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_126_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_74_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[23\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_50_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_119_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[8\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_67_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[17\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_5_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_59_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_59_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_59_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[6\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_5_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[18\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_75_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_75_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_75_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[7\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[19\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[1\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_91_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_91_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_91_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND3 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND3/X
+ sky130_fd_sc_hd__and4b_2
Xtap_3_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_111_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[2\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_137_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.DIBUF\[21\].cell DIBUF\[21\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DIBUF\[21\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[28\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[15\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[2\].DIODE\[7\] BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[11\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_31_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_24_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_17_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND4/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[12\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[21\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[24\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_20_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[11\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_116_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[20\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_29_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_132_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_132_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[8\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_45_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_45_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_45_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[17\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_61_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_61_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_131_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_61_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_124_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_72_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.ABUF\[0\] BLOCK\[1\].RAM32.A0BUF\[0\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A sky130_fd_sc_hd__clkbuf_2
Xtap_117_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[29\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell BLOCK\[1\].RAM32.TIE0\[1\].cell/LO
+ BLOCK\[1\].RAM32.FBUFENBUF0\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_65_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_58_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[3\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/X
+ sky130_fd_sc_hd__and4_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[12\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_86_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_86_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[30\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_106_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_86_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[13\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[31\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[25\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[14\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[8\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[26\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[15\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[27\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[9\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_86_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_79_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[10\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_15_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XDIBUF\[25\].cell Di0[25] VGND VGND VPWR VPWR DIBUF\[25\].cell/X sky130_fd_sc_hd__clkbuf_16
Xfill_22_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_31_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_31_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[7\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_127_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_127_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_103_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_51_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_44_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[19\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[28\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_37_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[6\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell BLOCK\[3\].RAM32.TIE0\[1\].cell/LO
+ BLOCK\[3\].RAM32.FBUFENBUF0\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_56_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[15\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[3\].Do_FF\[5\] BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X
+ BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[3\].MUX\[5\]/A1
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_56_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[2\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[29\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_72_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_72_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_72_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[3\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[12\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[28\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_122_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_70_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_115_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[24\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[2\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[11\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/X
+ sky130_fd_sc_hd__and4_2
Xfill_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_97_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_97_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_97_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xfill_114_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[25\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xfill_107_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_69_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_69_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_69_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.FBUFENBUF0\[3\].cell DEC0.AND2/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.FBUFENBUF0\[3\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_69_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_69_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_69_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND0/Y
+ sky130_fd_sc_hd__nor4b_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[8\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_106_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[20\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.TIE0\[0\].cell VGND VGND VPWR VPWR BLOCK\[2\].RAM32.TIE0\[0\].cell/HI
+ BLOCK\[2\].RAM32.TIE0\[0\].cell/LO sky130_fd_sc_hd__conb_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[3\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_91_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[21\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.DIBUF\[25\].cell DIBUF\[25\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DIBUF\[25\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xfill_84_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_77_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[4\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[22\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[31\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[16\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_26_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell BLOCK\[3\].RAM32.WEBUF\[2\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[5\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_99_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[17\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_42_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_42_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.DEC0.AND2 BLOCK\[1\].RAM32.DEC0.AND3/B BLOCK\[1\].RAM32.DEC0.AND3/A
+ BLOCK\[1\].RAM32.DEC0.AND3/C VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DEC0.AND2/X sky130_fd_sc_hd__and3b_2
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[1\].DIODE\[3\] BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[6\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[26\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[15\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_138_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_138_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[0\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[27\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_101_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_42_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_67_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_67_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[1\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_35_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_67_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[10\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_28_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_103_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_103_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_83_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_83_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_83_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF BLOCK\[1\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xfill_71_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_71_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[7\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[3\].DIODE\[0\] BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[23\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[19\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[2\].DIODE\[5\] BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[6\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_70_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[2\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[20\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[7\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.DIBUF\[6\].cell DIBUF\[6\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DIBUF\[6\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[19\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[3\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[2\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_12_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND0/Y
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[16\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_124_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_37_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[28\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_14_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_37_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND5/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_140_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_140_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[0\].Do_FF\[4\] BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X
+ BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[0\].MUX\[4\]/A3
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_53_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_53_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_53_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[11\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_97_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_8_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[12\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[21\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[24\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_78_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_78_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_78_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND0/Y
+ sky130_fd_sc_hd__nor4b_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_40_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[22\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_33_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_94_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_114_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_94_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_94_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.A0BUF\[3\].cell A0BUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DEC0.AND3/B
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[5\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[23\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell BLOCK\[2\].RAM32.TIE0\[3\].cell/LO
+ BLOCK\[2\].RAM32.FBUFENBUF0\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.DIBUF\[13\].cell DIBUF\[13\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DIBUF\[13\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[8\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[17\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[2\].Do_FF\[1\] BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X
+ BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[2\].MUX\[1\]/A2
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[6\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[18\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[1\].Do_FF\[6\] BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X
+ BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[1\].MUX\[6\]/A0
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[1\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[31\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[15\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[27\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_2_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xtap_23_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[14\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF BLOCK\[2\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[10\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_119_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[28\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_69_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[15\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_135_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_135_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[11\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_48_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[27\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_48_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_12_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[10\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_64_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_64_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_36_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND4 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND4/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_100_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_80_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_80_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_100_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_100_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_95_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_80_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_140_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_88_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[16\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_139_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_89_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_89_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_89_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_109_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[7\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[19\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[28\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[2\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[29\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND3/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[3\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[12\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[30\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[24\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[13\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[31\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_139_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_139_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[25\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_18_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[14\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[1\].DIODE\[1\] BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_52_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[26\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[8\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell BLOCK\[3\].RAM32.TIE0\[2\].cell/LO
+ BLOCK\[3\].RAM32.FBUFENBUF0\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[9\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_133_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_81_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_50_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_126_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_74_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_50_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_119_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_67_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_5_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF BLOCK\[3\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xtap_59_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_59_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[23\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_59_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_75_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[6\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_75_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_75_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[31\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[22\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.ABUF\[2\] BLOCK\[3\].RAM32.A0BUF\[2\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/C sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[18\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[27\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_111_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_91_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_91_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_91_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND4 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND4/X
+ sky130_fd_sc_hd__and4bb_2
Xtap_3_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[5\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_111_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[1\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[28\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[15\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[6\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_137_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[2\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[11\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[27\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.TIE0\[3\].cell VGND VGND VPWR VPWR BLOCK\[3\].RAM32.TIE0\[3\].cell/HI
+ BLOCK\[3\].RAM32.TIE0\[3\].cell/LO sky130_fd_sc_hd__conb_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[1\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[10\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[24\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_31_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_24_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.DIBUF\[17\].cell DIBUF\[17\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DIBUF\[17\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[7\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_20_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[19\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[0\].Do_FF\[2\] BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X
+ BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[0\].MUX\[2\]/A1
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_29_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_132_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[2\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[20\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_45_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_45_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[3\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[21\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_61_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_61_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[30\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF BLOCK\[0\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xtap_131_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_124_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_72_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[4\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_117_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_65_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[31\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_58_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[16\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_10_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[5\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_86_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_86_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[14\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_106_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND6/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_86_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell BLOCK\[2\].RAM32.WEBUF\[0\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[26\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[17\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_122_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[0\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[23\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_86_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[6\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[22\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[9\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[18\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[5\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[23\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell BLOCK\[0\].RAM32.TIE0\[1\].cell/LO
+ BLOCK\[0\].RAM32.FBUFENBUF0\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_15_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[19\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_22_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[6\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_15_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_31_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[18\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_31_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[2\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_127_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_51_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[1\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_44_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_37_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_56_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_2_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_56_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[15\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_72_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_72_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell BLOCK\[1\].RAM32.WEBUF\[1\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[27\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell BLOCK\[0\].RAM32.TIE0\[2\].cell/LO
+ BLOCK\[0\].RAM32.FBUFENBUF0\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_122_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_70_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_115_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[10\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[28\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_63_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_121_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xtap_108_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_97_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_97_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_117_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_114_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_97_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_107_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[11\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_69_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_69_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_69_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_69_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_69_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND1 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND1/X
+ sky130_fd_sc_hd__and4bb_2
XDIBUF\[31\].cell Di0[31] VGND VGND VPWR VPWR DIBUF\[31\].cell/X sky130_fd_sc_hd__clkbuf_16
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[12\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xfill_106_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_106_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[21\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[22\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[16\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[5\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[2\].DIODE\[7\] BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_77_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[17\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND4/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[0\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_26_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[31\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_99_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_42_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.DEC0.AND3 BLOCK\[1\].RAM32.DEC0.AND3/A BLOCK\[1\].RAM32.DEC0.AND3/B
+ BLOCK\[1\].RAM32.DEC0.AND3/C VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DEC0.AND3/X sky130_fd_sc_hd__and3_2
Xtap_42_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[30\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_138_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_138_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[14\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell BLOCK\[0\].RAM32.WEBUF\[2\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[26\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_101_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[31\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[13\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_42_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_67_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[9\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_67_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_67_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_35_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[27\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[14\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_28_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_103_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_103_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_83_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_83_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_83_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_103_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[10\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[26\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.DIBUF\[31\].cell DIBUF\[31\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DIBUF\[31\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[3\].RAM32.FBUFENBUF0\[2\].cell DEC0.AND3/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.FBUFENBUF0\[2\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[9\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_71_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_71_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_112_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.ENBUF BLOCK\[0\].RAM32.DEC0.AND2/X VGND VGND
+ VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/D sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[23\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_70_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XDo0MUX.M\[1\].DIODE_A0MUX\[15\] Do0MUX.M\[1\].MUX\[7\]/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[6\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[18\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[27\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[7\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF BLOCK\[2\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[1\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[28\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[2\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_82_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[11\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[29\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[12\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_14_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[30\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_37_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_37_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_140_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.TIE0\[0\].cell VGND VGND VPWR VPWR BLOCK\[0\].RAM32.TIE0\[0\].cell/HI
+ BLOCK\[0\].RAM32.TIE0\[0\].cell/LO sky130_fd_sc_hd__conb_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_53_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_53_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[24\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_7_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[13\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_97_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_8_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[25\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[2\].DIODE_A0MUX\[19\] Do0MUX.M\[2\].MUX\[3\]/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[3\].Do_FF\[5\] BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X
+ BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[3\].MUX\[5\]/A2
+ sky130_fd_sc_hd__dfxtp_1
Xtap_78_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_78_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[8\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND1 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND1/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_78_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_40_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_33_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell BLOCK\[3\].RAM32.WEBUF\[2\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X sky130_fd_sc_hd__clkbuf_2
Xtap_94_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[0\].DIODE_A1MUX\[2\] Do0MUX.M\[0\].MUX\[2\]/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_114_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_114_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_94_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_94_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[22\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[31\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND2/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_130_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[5\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[30\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[21\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[17\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[4\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[31\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[0\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[18\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[27\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[14\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[5\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[17\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[1\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[26\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[0\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell BLOCK\[0\].RAM32.TIE0\[0\].cell/LO
+ BLOCK\[0\].RAM32.FBUFENBUF0\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_23_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF BLOCK\[3\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[23\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_135_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_48_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_48_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[6\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_12_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[9\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[18\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_64_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_64_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[7\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_5_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_36_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND5 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND5/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell BLOCK\[2\].RAM32.WEBUF\[3\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X sky130_fd_sc_hd__clkbuf_2
Xtap_80_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_100_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_100_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_100_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_95_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[19\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_80_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_88_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xfill_139_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_109_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_89_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_89_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_89_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[2\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[20\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_109_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_125_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[3\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[21\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[30\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[4\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[2\].DIODE_A2MUX\[23\] Do0MUX.M\[2\].MUX\[7\]/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[3\].DIODE\[0\] BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.ABUF\[2\] BLOCK\[0\].RAM32.A0BUF\[2\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[25\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[16\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[2\].DIODE\[5\] BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_139_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_139_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_139_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[13\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[22\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_52_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[12\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_45_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDIBUF\[0\].cell Di0[0] VGND VGND VPWR VPWR DIBUF\[0\].cell/X sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF BLOCK\[0\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[21\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[8\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_0_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[17\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_81_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_126_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_74_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_50_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_50_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.FBUFENBUF0\[0\].cell DEC0.AND0/Y VGND VGND VPWR VPWR BLOCK\[0\].RAM32.FBUFENBUF0\[0\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[22\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[3\].DIODE_A2MUX\[27\] Do0MUX.M\[3\].MUX\[3\]/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_119_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[18\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_67_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_5_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_59_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_59_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[5\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_5_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND5/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[17\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[1\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_75_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_75_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_75_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_10_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[0\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_111_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_91_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_91_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND5 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND5/X
+ sky130_fd_sc_hd__and4b_2
Xtap_3_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_111_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_111_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_91_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[31\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_93_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_138_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[14\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xfill_137_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.ENBUF BLOCK\[1\].RAM32.DEC0.AND1/X VGND VGND
+ VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[26\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[15\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[2\].Do_FF\[1\] BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X
+ BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[2\].MUX\[1\]/A3
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[9\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[27\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[10\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[1\].Do_FF\[6\] BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X
+ BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[1\].MUX\[6\]/A1
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xfill_24_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xfill_17_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[11\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[20\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[21\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_29_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_29_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[4\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_45_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_45_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[16\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_61_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[3\].Do_FF\[3\] BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X
+ BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[3\].MUX\[3\]/A0
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[7\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_61_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_131_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_124_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_72_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[30\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_117_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_65_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell BLOCK\[2\].RAM32.CLKBUF.cell/X VGND
+ VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X sky130_fd_sc_hd__clkbuf_2
Xtap_58_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.ABUF\[0\] BLOCK\[2\].RAM32.A0BUF\[0\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A sky130_fd_sc_hd__clkbuf_2
Xtap_86_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[29\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[13\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_106_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_106_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_86_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_86_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell BLOCK\[2\].RAM32.TIE0\[1\].cell/LO
+ BLOCK\[2\].RAM32.FBUFENBUF0\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[25\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.DIBUF\[23\].cell DIBUF\[23\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DIBUF\[23\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xtap_122_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[30\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[12\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_122_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[8\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[26\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[13\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_142_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[9\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[25\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[8\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND3/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[22\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[31\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_22_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_15_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[5\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_31_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[17\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[6\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.TIE0\[3\].cell VGND VGND VPWR VPWR BLOCK\[1\].RAM32.TIE0\[3\].cell/HI
+ BLOCK\[1\].RAM32.TIE0\[3\].cell/LO sky130_fd_sc_hd__conb_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[1\].DIODE\[1\] BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[15\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[0\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_44_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[18\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[27\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_37_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_2_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[0\].DIODE\[6\] BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_56_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_56_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[1\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[28\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_72_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_72_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[2\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[11\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[29\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_122_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_70_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_115_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell BLOCK\[1\].RAM32.TIE0\[0\].cell/LO
+ BLOCK\[1\].RAM32.FBUFENBUF0\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_63_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.WEBUF\[1\].cell WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.WEBUF\[1\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[12\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_121_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_108_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_97_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_97_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_56_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_117_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_117_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_114_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_97_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[24\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_69_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_69_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xfill_69_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_69_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_69_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_133_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND2 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND2/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_106_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_106_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[7\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[21\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[4\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[20\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[16\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[21\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[3\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[30\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[17\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_26_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[26\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[4\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[16\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_42_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[0\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[25\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_42_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[0\].Do_FF\[2\] BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X
+ BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[0\].MUX\[2\]/A2
+ sky130_fd_sc_hd__dfxtp_1
Xtap_138_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.DIBUF\[9\].cell DIBUF\[9\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DIBUF\[9\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_101_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_67_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_42_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_67_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_35_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_28_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[13\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[22\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_103_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_103_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_83_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_83_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_83_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_103_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_16_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND1/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[23\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XDo0MUX.M\[0\].DIODE_A2MUX\[7\] Do0MUX.M\[0\].MUX\[7\]/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[8\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[17\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_71_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_120_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[6\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.ENBUF BLOCK\[2\].RAM32.DEC0.AND0/Y VGND VGND
+ VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND6/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_128_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[18\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_112_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[7\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[0\].MUX\[1\] Do0MUX.M\[0\].MUX\[1\]/A0 Do0MUX.M\[0\].MUX\[1\]/A1 Do0MUX.M\[0\].MUX\[1\]/A2
+ Do0MUX.M\[0\].MUX\[1\]/A3 Do0MUX.SEL0BUF\[0\]/X Do0MUX.SEL1BUF\[0\]/X VGND VGND
+ VPWR VPWR Do0[1] sky130_fd_sc_hd__mux4_1
Xfill_105_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[1\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[19\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell BLOCK\[1\].RAM32.WEBUF\[1\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.DIBUF\[27\].cell DIBUF\[27\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DIBUF\[27\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[2\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[20\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[29\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[3\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_82_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[15\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_75_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_37_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_37_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF BLOCK\[3\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_53_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_53_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[12\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[21\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_97_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_8_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[24\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_8_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[11\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[20\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_78_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_78_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_40_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND2 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND2/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[21\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_33_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_114_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_114_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[8\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[17\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_94_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_94_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_94_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_114_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[4\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_19_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[16\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_130_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_130_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XA0BUF\[0\].cell A0[0] VGND VGND VPWR VPWR A0BUF\[0\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell BLOCK\[0\].RAM32.WEBUF\[2\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell BLOCK\[3\].RAM32.TIE0\[3\].cell/LO
+ BLOCK\[3\].RAM32.FBUFENBUF0\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[30\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[13\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[31\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[25\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF BLOCK\[0\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[14\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[8\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[26\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[3\].MUX\[6\] Do0MUX.M\[3\].MUX\[6\]/A0 Do0MUX.M\[3\].MUX\[6\]/A1 Do0MUX.M\[3\].MUX\[6\]/A2
+ Do0MUX.M\[3\].MUX\[6\]/A3 Do0MUX.SEL0BUF\[3\]/X Do0MUX.SEL1BUF\[3\]/X VGND VGND
+ VPWR VPWR Do0[30] sky130_fd_sc_hd__mux4_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[15\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[9\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[27\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND4/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XDo0MUX.M\[1\].DIODE_A2MUX\[12\] Do0MUX.M\[1\].MUX\[4\]/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[10\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_48_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_48_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_12_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_64_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_64_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[20\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[11\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_5_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.DIBUF\[10\].cell DIBUF\[10\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DIBUF\[10\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xfill_36_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_80_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.DIBUF\[2\].cell DIBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DIBUF\[2\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND6 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND6/X
+ sky130_fd_sc_hd__and4b_2
Xtap_100_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_100_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_100_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_95_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_80_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_88_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_139_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_109_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_89_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_89_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_109_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_109_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_89_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[6\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[15\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[0\].DIODE_A3MUX\[1\] Do0MUX.M\[0\].MUX\[1\]/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_125_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_125_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[29\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_141_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[3\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[28\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[2\].DIODE_A2MUX\[16\] Do0MUX.M\[2\].MUX\[0\]/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[12\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[24\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[2\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[29\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[11\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[25\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[12\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_139_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_139_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_139_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[8\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[24\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_139_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell BLOCK\[2\].RAM32.TIE0\[0\].cell/LO
+ BLOCK\[2\].RAM32.FBUFENBUF0\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xfill_52_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[0\].Do_FF\[0\] BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X
+ BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[0\].MUX\[0\]/A0
+ sky130_fd_sc_hd__dfxtp_1
Xfill_45_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfill_38_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_0_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[21\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_50_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_50_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_74_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_119_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_67_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_59_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[4\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[22\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[31\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_59_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[16\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[5\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_75_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_75_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF BLOCK\[1\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xtap_10_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_111_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_91_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_91_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[17\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[26\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND6 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND6/X
+ sky130_fd_sc_hd__and4b_2
Xtap_3_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_111_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_111_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_91_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[6\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[15\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_93_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[3\].Do_FF\[5\] BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X
+ BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[3\].MUX\[5\]/A3
+ sky130_fd_sc_hd__dfxtp_1
Xtap_138_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[0\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_86_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[27\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell BLOCK\[1\].RAM32.CLKBUF.cell/X VGND
+ VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X sky130_fd_sc_hd__clkbuf_2
Xfill_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[1\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[10\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[28\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_136_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND2/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XDIBUF\[14\].cell Di0[14] VGND VGND VPWR VPWR DIBUF\[14\].cell/X sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[11\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell BLOCK\[2\].RAM32.WEBUF\[3\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[23\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_24_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_0_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell BLOCK\[0\].RAM32.TIE0\[3\].cell/LO
+ BLOCK\[0\].RAM32.FBUFENBUF0\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[6\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[20\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[7\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_29_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[3\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[19\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_45_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_45_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[20\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[2\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_61_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[29\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_61_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_131_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[16\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_124_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_72_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[3\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_117_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_65_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_10_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_58_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_86_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_106_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_106_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_86_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_19_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_122_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_122_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_122_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_1_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF BLOCK\[2\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[12\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[21\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.DIBUF\[14\].cell DIBUF\[14\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DIBUF\[14\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xfill_142_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDo0MUX.SEL1BUF\[2\] DEC0.AND3/A VGND VGND VPWR VPWR Do0MUX.SEL1BUF\[2\]/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[24\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_135_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[22\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.DIBUF\[19\].cell DIBUF\[19\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DIBUF\[19\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[5\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[23\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[8\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[17\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[2\].DIODE\[5\] BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[6\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[18\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_15_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[1\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[19\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[2\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_37_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[31\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_56_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_56_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF BLOCK\[0\].RAM32.SLICE\[2\].RAM8.DEC0.AND0/Y
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[14\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_72_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_72_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[28\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND5/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[15\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_122_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_70_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[11\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_115_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_63_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[27\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_108_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_97_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell BLOCK\[1\].RAM32.TIE0\[2\].cell/LO
+ BLOCK\[1\].RAM32.FBUFENBUF0\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_56_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_117_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_117_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_117_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_114_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_97_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_97_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_49_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_69_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_69_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[10\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_69_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_69_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_69_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_133_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND3 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND3/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_133_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[11\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xfill_106_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfill_106_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[20\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[16\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_34_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[1\].Do_FF\[6\] BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X
+ BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[1\].MUX\[6\]/A2
+ sky130_fd_sc_hd__dfxtp_1
Xfill_77_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF BLOCK\[3\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[29\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XDo0MUX.M\[1\].DIODE_A1MUX\[9\] Do0MUX.M\[1\].MUX\[1\]/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[3\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[12\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[30\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_20_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[24\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_42_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.DIBUF\[5\].cell DIBUF\[5\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DIBUF\[5\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[13\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[31\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_101_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[25\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[14\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_42_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[8\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_67_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_67_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_35_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[26\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_28_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[3\].Do_FF\[3\] BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X
+ BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[3\].MUX\[3\]/A1
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_103_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_83_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_83_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_103_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_103_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[9\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_16_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell BLOCK\[3\].RAM32.TIE0\[0\].cell/LO
+ BLOCK\[3\].RAM32.FBUFENBUF0\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_71_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[19\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[10\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_32_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_120_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_113_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_128_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_128_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_112_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[22\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_105_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[31\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[5\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[28\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[6\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[15\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.A0BUF\[2\].cell A0BUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.A0BUF\[2\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[2\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[27\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[11\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND3/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF BLOCK\[0\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[1\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_82_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[28\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[10\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_75_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[24\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_68_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[11\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_37_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_53_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_53_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_97_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[1\].DIODE\[1\] BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_8_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[0\].DIODE\[6\] BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_78_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_78_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_40_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[20\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND3 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND3/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_33_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_114_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_114_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_94_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_94_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_114_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_19_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[3\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[21\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[30\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XDo0MUX.SEL_DIODE\[0\] DEC0.AND3/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_130_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_130_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_130_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[4\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[31\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[16\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[5\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[14\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[17\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[2\].DIODE\[3\] BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[26\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[0\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[27\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[1\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[10\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[22\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_48_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_48_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[5\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF BLOCK\[1\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[23\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_12_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_64_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_64_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[0\].Do_FF\[2\] BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X
+ BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[0\].MUX\[2\]/A3
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[19\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[6\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_5_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_36_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[2\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/B BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/C
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.DEC0.AND7/X
+ sky130_fd_sc_hd__and4_2
Xtap_100_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_100_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_100_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_95_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_80_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_80_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[18\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_88_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_13_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[7\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_139_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_109_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_89_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_89_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[19\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[1\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_109_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_109_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_89_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_125_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_125_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_125_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND1/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[2\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_31_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_141_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_141_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell BLOCK\[0\].RAM32.CLKBUF.cell/X VGND
+ VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[28\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[1\].Do_FF\[4\] BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X
+ BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[1\].MUX\[4\]/A0
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.ABUF\[2\] BLOCK\[1\].RAM32.A0BUF\[2\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[11\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_139_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XDo0MUX.M\[3\].DIODE_A0MUX\[28\] Do0MUX.M\[3\].MUX\[4\]/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_139_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_139_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_139_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_139_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[12\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[21\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.CLKBUF.cell CLKBUF.cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.CLKBUF.cell/X
+ sky130_fd_sc_hd__clkbuf_4
Xfill_52_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_45_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_38_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[22\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xfill_0_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[16\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[5\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_50_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_67_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[17\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.WEBUF\[0\].cell WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.WEBUF\[0\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_59_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_5_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_59_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[0\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[18\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_75_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_75_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_10_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[1\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_91_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_111_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_111_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_111_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_91_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/X
+ sky130_fd_sc_hd__and4_2
Xtap_3_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[30\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_24_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_93_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_138_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_86_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_79_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[13\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[31\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_40_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND0/Y
+ sky130_fd_sc_hd__nor4b_2
Xfill_137_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[3\].RAM32.EN0BUF.cell DEC0.AND3/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DEC0.AND3/C
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[27\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_136_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_136_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[14\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[10\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF BLOCK\[2\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[26\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[15\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[9\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_141_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_0_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[10\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[19\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_50_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_45_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[7\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[28\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_61_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_61_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_131_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND4/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_124_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[2\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_72_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_117_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[11\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[29\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_65_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDIBUF\[20\].cell Di0[20] VGND VGND VPWR VPWR DIBUF\[20\].cell/X sky130_fd_sc_hd__clkbuf_16
Xtap_58_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_106_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_106_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[12\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_86_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_86_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[30\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_19_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[24\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_122_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[13\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.ABUF\[0\] BLOCK\[3\].RAM32.A0BUF\[0\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND7/A sky130_fd_sc_hd__clkbuf_2
Xtap_122_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_122_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_1_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_35_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell BLOCK\[3\].RAM32.TIE0\[1\].cell/LO
+ BLOCK\[3\].RAM32.FBUFENBUF0\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[25\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xfill_142_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[8\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[26\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_135_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_128_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[9\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[21\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[30\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[4\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[31\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[18\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[27\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[5\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_98_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[14\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[0\].Do_FF\[0\] BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X
+ BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[0\].MUX\[0\]/A1
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[1\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[26\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[17\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_2_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[15\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_56_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_56_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.DIBUF\[20\].cell DIBUF\[20\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DIBUF\[20\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[0\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[27\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_72_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_72_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[10\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[1\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND0/Y
+ sky130_fd_sc_hd__nor4b_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.DIBUF\[25\].cell DIBUF\[25\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DIBUF\[25\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_122_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_70_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_115_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_63_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_108_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_97_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_56_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_117_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_117_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_117_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_97_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_97_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_49_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_69_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_69_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_69_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_69_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_69_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_133_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_133_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND4 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND4/X
+ sky130_fd_sc_hd__and4bb_2
Xtap_133_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[7\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[19\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_106_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[2\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[20\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[7\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_34_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_34_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND2/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[3\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[21\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[30\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[4\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[16\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[25\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_20_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.DIBUF\[1\].cell DIBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DIBUF\[1\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xfill_13_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[26\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[0\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[9\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_42_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_67_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_67_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDIBUF\[6\].cell Di0[6] VGND VGND VPWR VPWR DIBUF\[6\].cell/X sky130_fd_sc_hd__clkbuf_16
Xtap_35_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_28_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[12\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[21\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_103_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_83_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_83_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_103_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_103_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[22\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_32_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[18\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_120_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_71_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[5\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_128_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[23\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[0\].DIODE_A0MUX\[6\] Do0MUX.M\[0\].MUX\[6\]/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_128_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_128_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_113_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_61_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[1\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_106_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[17\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_112_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[6\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_105_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[18\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[0\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[1\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell BLOCK\[0\].RAM32.TIE0\[1\].cell/LO
+ BLOCK\[0\].RAM32.FBUFENBUF0\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[15\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[27\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[2\].DIODE\[5\] BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDo0MUX.M\[1\].DIODE_A3MUX\[8\] Do0MUX.M\[1\].MUX\[0\]/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_75_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_68_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[10\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[15\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_53_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[11\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_97_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[20\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_8_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[21\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_78_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_78_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF BLOCK\[1\].RAM32.SLICE\[2\].RAM8.DEC0.AND0/Y
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND4 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND4/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[4\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_40_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_114_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_94_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_94_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[16\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_26_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_114_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_114_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[7\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[3\].DIODE\[7\] BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_130_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_130_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_130_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[17\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_43_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[0\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[29\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.DIBUF\[29\].cell DIBUF\[29\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DIBUF\[29\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xfill_110_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[12\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[30\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XDo0MUX.M\[1\].DIODE_A0MUX\[13\] Do0MUX.M\[1\].MUX\[5\]/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[26\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[13\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[9\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[25\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[14\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[23\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[8\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[1\].Do_FF\[6\] BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X
+ BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[1\].MUX\[6\]/A3
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[26\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xfill_80_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[9\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_48_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_12_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_64_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_64_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_5_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_36_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_100_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_100_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_95_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_80_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_80_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_88_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[2\].DIODE_A0MUX\[17\] Do0MUX.M\[2\].MUX\[1\]/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[6\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[15\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_139_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_89_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[18\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_109_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_109_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_109_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_89_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[27\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[3\].Do_FF\[3\] BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X
+ BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[3\].MUX\[3\]/A2
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF BLOCK\[2\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_125_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_125_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[1\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_31_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_125_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[28\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_24_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_38_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[0\].DIODE_A1MUX\[0\] Do0MUX.M\[0\].MUX\[0\]/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[15\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_141_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_141_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_141_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[2\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[11\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[29\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[12\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[24\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_139_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_139_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_139_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_139_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[25\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_139_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_139_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[7\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_52_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[8\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_38_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_0_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND3/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[20\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.DIBUF\[12\].cell DIBUF\[12\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DIBUF\[12\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xtap_5_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[3\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_59_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_59_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[21\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[30\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[17\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[26\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_75_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_75_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[4\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_10_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[31\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[0\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_91_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[25\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[16\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_111_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_111_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_111_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_91_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[14\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_24_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[5\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[0\].DIODE\[6\] BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_24_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_93_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_138_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_86_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[26\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_79_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_40_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND1 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND1/X
+ sky130_fd_sc_hd__and4bb_2
Xfill_137_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_40_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[9\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[0\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_136_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_136_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_136_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF BLOCK\[3\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[23\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[2\].DIODE_A2MUX\[21\] Do0MUX.M\[2\].MUX\[5\]/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.ABUF\[0\] BLOCK\[0\].RAM32.A0BUF\[0\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[6\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_141_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[2\].DIODE\[3\] BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_0_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[18\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[7\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[23\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[1\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[19\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell BLOCK\[1\].RAM32.TIE0\[3\].cell/LO
+ BLOCK\[1\].RAM32.FBUFENBUF0\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[6\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[2\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[20\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[29\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_50_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[3\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_61_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_124_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_72_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[3\].DIODE_A2MUX\[25\] Do0MUX.M\[3\].MUX\[1\]/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_117_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[15\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_65_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_10_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_58_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[25\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[16\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_106_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_106_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_86_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_86_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_19_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_122_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_122_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_122_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_1_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_35_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_35_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_91_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[11\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[20\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_136_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_51_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.A0BUF\[1\].cell A0BUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.A0BUF\[1\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_142_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND1/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xfill_135_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[21\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_128_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF BLOCK\[0\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[8\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[17\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[4\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[22\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XA0BUF\[6\].cell A0[6] VGND VGND VPWR VPWR DEC0.AND3/A sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND6/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[16\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[5\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[1\].DIODE_A3MUX\[15\] Do0MUX.M\[1\].MUX\[7\]/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[1\].Do_FF\[4\] BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X
+ BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[1\].MUX\[4\]/A1
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[17\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_15_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[0\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_98_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[31\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_2_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[14\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_56_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[26\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[15\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_72_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_72_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[3\].Do_FF\[1\] BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X
+ BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[3\].MUX\[1\]/A0
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND1 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND1/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[9\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[27\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[14\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[23\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_122_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_70_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_21_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[2\].DIODE_A3MUX\[19\] Do0MUX.M\[2\].MUX\[3\]/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_115_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[10\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_63_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_108_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_56_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_117_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_117_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_117_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_97_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_97_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xfill_69_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_49_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_69_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_69_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_69_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[11\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.DIBUF\[8\].cell DIBUF\[8\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DIBUF\[8\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.DIBUF\[16\].cell DIBUF\[16\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DIBUF\[16\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xtap_133_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_69_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[20\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND5 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND5/X
+ sky130_fd_sc_hd__and4b_2
Xtap_133_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_133_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell BLOCK\[2\].RAM32.TIE0\[2\].cell/LO
+ BLOCK\[2\].RAM32.FBUFENBUF0\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_46_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_106_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_34_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_140_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[6\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_34_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[15\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[16\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[28\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.DIBUF\[31\].cell DIBUF\[31\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DIBUF\[31\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[2\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[11\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[29\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_20_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_13_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[25\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[30\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[12\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[8\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[24\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[13\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[14\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_42_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_67_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_67_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_35_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[25\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_28_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[0\].DIODE\[4\] BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_83_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_103_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_103_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_103_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_83_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[8\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_16_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_32_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_71_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[22\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_120_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_128_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_128_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_128_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[31\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_113_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_61_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_106_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_54_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_112_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[5\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_105_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[17\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[26\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[6\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[31\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[15\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[0\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[27\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[5\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[14\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[1\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[10\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[28\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[11\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_68_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[23\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[24\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xfill_9_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[6\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_8_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[0\].Do_FF\[0\] BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X
+ BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[0\].MUX\[0\]/A2
+ sky130_fd_sc_hd__dfxtp_1
Xtap_8_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF BLOCK\[2\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell BLOCK\[0\].RAM32.TIE0\[0\].cell/LO
+ BLOCK\[0\].RAM32.FBUFENBUF0\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[7\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_78_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_78_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND5 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND5/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[19\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_40_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_33_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_114_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_94_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_94_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_114_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_114_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_19_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[2\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[20\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_27_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[29\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_130_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_130_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_130_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[16\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[3\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_43_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_43_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[0\].DIODE_A2MUX\[5\] Do0MUX.M\[0\].MUX\[5\]/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[30\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_139_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[13\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[4\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[16\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_110_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[25\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_103_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND2/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[22\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[5\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[23\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xfill_80_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[8\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[17\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_73_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[6\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[22\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_64_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[18\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[5\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_5_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_36_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_100_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_100_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_95_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[1\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_80_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_80_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[19\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_88_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_89_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_139_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_109_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_109_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_109_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_89_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[2\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[31\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_125_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_125_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_31_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_125_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_38_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_38_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[14\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_24_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[24\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_141_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_141_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.WEBUF\[3\].cell WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.WEBUF\[3\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
Xtap_54_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[15\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[27\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF BLOCK\[3\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[10\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_139_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_139_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_139_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_139_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_139_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_139_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.ABUF\[2\] BLOCK\[2\].RAM32.A0BUF\[2\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[11\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[20\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_52_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[16\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[21\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_0_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDo0MUX.M\[3\].MUX\[4\] Do0MUX.M\[3\].MUX\[4\]/A0 Do0MUX.M\[3\].MUX\[4\]/A1 Do0MUX.M\[3\].MUX\[4\]/A2
+ Do0MUX.M\[3\].MUX\[4\]/A3 Do0MUX.SEL0BUF\[3\]/X Do0MUX.SEL1BUF\[3\]/X VGND VGND
+ VPWR VPWR Do0[28] sky130_fd_sc_hd__mux4_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[4\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[16\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_5_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_59_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0MUX.M\[1\].DIODE_A2MUX\[10\] Do0MUX.M\[1\].MUX\[2\]/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_75_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_75_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[30\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_111_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_111_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_91_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_91_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[13\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_111_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[31\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_24_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_93_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_138_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[25\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_86_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF BLOCK\[2\].RAM32.SLICE\[2\].RAM8.DEC0.AND0/Y
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_79_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[30\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF BLOCK\[0\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xtap_40_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_40_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND2 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND2/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[14\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_40_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_136_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_136_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[8\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[26\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_136_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_49_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[13\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[3\].DIODE\[7\] BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDo0MUX.M\[2\].MUX\[6\] Do0MUX.M\[2\].MUX\[6\]/A0 Do0MUX.M\[2\].MUX\[6\]/A1 Do0MUX.M\[2\].MUX\[6\]/A2
+ Do0MUX.M\[2\].MUX\[6\]/A3 Do0MUX.SEL0BUF\[2\]/X Do0MUX.SEL1BUF\[2\]/X VGND VGND
+ VPWR VPWR Do0[22] sky130_fd_sc_hd__mux4_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[9\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND5/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[10\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[19\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_141_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_0_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[22\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[31\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[5\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_50_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[6\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[15\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_43_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfill_36_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[27\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[1\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[10\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_72_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[28\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_117_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_65_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_10_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_58_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[24\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_106_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_86_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_86_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[29\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[11\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_106_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_19_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[12\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_122_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_122_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_122_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_35_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_35_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[24\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[3\].Do_FF\[3\] BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X
+ BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[3\].MUX\[3\]/A3
+ sky130_fd_sc_hd__dfxtp_1
Xtap_91_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_51_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_51_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_136_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_84_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_142_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_129_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_128_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell BLOCK\[3\].RAM32.WEBUF\[0\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[21\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[30\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell BLOCK\[1\].RAM32.TIE0\[0\].cell/LO
+ BLOCK\[1\].RAM32.FBUFENBUF0\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[4\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[31\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[16\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[5\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[30\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[14\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[17\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[26\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF BLOCK\[1\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[4\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_98_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[13\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[0\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[27\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_2_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_2_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[1\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[10\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_72_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND2 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND2/X
+ sky130_fd_sc_hd__and4bb_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell BLOCK\[0\].RAM32.TIE0\[2\].cell/LO
+ BLOCK\[0\].RAM32.FBUFENBUF0\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_122_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[22\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_70_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_115_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_63_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_108_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_117_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_117_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[5\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_97_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_97_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[23\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_56_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_117_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_49_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xfill_69_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_69_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_69_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_69_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.DIBUF\[4\].cell DIBUF\[4\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DIBUF\[4\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xtap_133_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND6 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND6/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[0\].DIODE\[6\] BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_133_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_133_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[6\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_46_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell BLOCK\[2\].RAM32.WEBUF\[1\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_46_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_106_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[18\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[7\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_62_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[1\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[19\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_34_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDo0MUX.SEL1BUF\[0\] DEC0.AND3/A VGND VGND VPWR VPWR Do0MUX.SEL1BUF\[0\]/X sky130_fd_sc_hd__clkbuf_2
Xfill_140_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_34_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_34_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_133_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[20\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[2\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[29\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[3\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[2\].DIODE\[3\] BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[24\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.DIBUF\[22\].cell DIBUF\[22\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DIBUF\[22\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[12\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[21\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_67_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_35_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_28_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[22\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_83_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_103_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_103_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_83_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_16_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[16\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_16_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[5\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[21\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_32_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[17\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_71_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[4\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_32_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_120_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_128_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_128_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_128_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_113_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_61_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_106_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[0\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[18\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_54_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_112_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_47_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_105_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[1\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_57_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[30\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND1/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[13\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[31\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[14\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell BLOCK\[1\].RAM32.TIE0\[1\].cell/LO
+ BLOCK\[1\].RAM32.FBUFENBUF0\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND6/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[26\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[1\].Do_FF\[4\] BLOCK\[2\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X
+ BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[1\].MUX\[4\]/A2
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[15\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_68_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[9\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[10\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[19\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_9_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xtap_8_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[20\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_78_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_78_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND6 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND6/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[3\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_40_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_33_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_94_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_26_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_114_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_114_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_94_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[3\].Do_FF\[1\] BLOCK\[1\].RAM32.Do0_REG.Do_CLKBUF\[3\]/X
+ BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[25\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[3\].MUX\[1\]/A1
+ sky130_fd_sc_hd__dfxtp_1
Xtap_19_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_130_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_130_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDIBUF\[26\].cell Di0[26] VGND VGND VPWR VPWR DIBUF\[26\].cell/X sky130_fd_sc_hd__clkbuf_16
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_130_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_43_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_43_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_43_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[29\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF BLOCK\[3\].RAM32.SLICE\[2\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[12\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_111_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[30\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[24\].cell/X BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_110_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_103_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[29\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[13\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[25\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[12\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[8\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[26\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[9\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_80_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_73_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[21\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[30\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_66_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[4\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[31\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell BLOCK\[2\].RAM32.TIE0\[0\].cell/LO
+ BLOCK\[2\].RAM32.FBUFENBUF0\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_100_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_95_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_80_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.TIE0\[1\].cell VGND VGND VPWR VPWR BLOCK\[2\].RAM32.TIE0\[1\].cell/HI
+ BLOCK\[2\].RAM32.TIE0\[1\].cell/LO sky130_fd_sc_hd__conb_1
Xtap_100_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_88_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[5\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[14\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_13_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_109_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_109_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_109_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_89_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_89_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[17\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.Do0_REG.OUTREG_BYTE\[0\].DIODE\[4\] BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.DIBUF\[26\].cell DIBUF\[26\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.DIBUF\[26\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[26\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[15\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_125_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[0\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND4/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_125_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_125_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[27\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_31_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_38_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_38_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_38_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_141_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_141_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[1\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell BLOCK\[3\].RAM32.WEBUF\[3\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X sky130_fd_sc_hd__clkbuf_2
Xtap_54_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_54_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[28\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF BLOCK\[0\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[10\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[11\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_70_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[2\].DIODE\[1\] BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_139_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_139_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_139_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_139_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_139_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[2\] BLOCK\[0\].RAM32.Do0_REG.Root_CLKBUF/X VGND
+ VGND VPWR VPWR BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[2\]/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[20\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[7\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_0_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[3\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[21\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[30\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_5_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[4\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[20\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[29\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[16\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[25\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_75_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[3\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.DIBUF\[7\].cell DIBUF\[7\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DIBUF\[7\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xtap_10_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[0\].Do_FF\[0\] BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[0\]/X
+ BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[0\].MUX\[0\]/A3
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_111_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_111_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_91_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_91_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[26\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_3_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_93_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XDo0MUX.M\[2\].DIODE_A0MUX\[22\] Do0MUX.M\[2\].MUX\[6\]/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_138_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_86_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[0\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[9\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_79_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND3 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND3/X
+ sky130_fd_sc_hd__and4b_2
Xtap_40_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_40_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_40_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_136_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_136_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_136_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[12\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_49_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_49_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[21\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[22\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_65_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[5\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[23\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xfill_141_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF BLOCK\[1\].RAM32.SLICE\[1\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
Xfill_0_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[17\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[1\].Do_FF\[2\] BLOCK\[0\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X
+ BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[10\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[1\].MUX\[2\]/A0
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[6\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.ABUF\[0\] BLOCK\[1\].RAM32.A0BUF\[0\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[0\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[18\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XDo0MUX.M\[3\].DIODE_A0MUX\[26\] Do0MUX.M\[3\].MUX\[2\]/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[7\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[19\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.A0BUF\[4\].cell A0BUF\[4\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.DEC0.AND3/A
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[1\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_50_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[28\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell BLOCK\[2\].RAM32.TIE0\[3\].cell/LO
+ BLOCK\[2\].RAM32.FBUFENBUF0\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_43_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.DIBUF\[14\].cell DIBUF\[14\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.DIBUF\[14\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xfill_36_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[2\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_29_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_65_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_58_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_10_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_106_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_86_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_86_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_106_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[15\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_19_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[11\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[20\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_122_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_122_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_35_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_35_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[21\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_91_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_51_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_51_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_136_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_84_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_51_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_142_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_129_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_77_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[4\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[20\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_128_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[16\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[3\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[17\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell BLOCK\[0\].RAM32.WEBUF\[0\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[0\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[29\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[12\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[30\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[13\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_2_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[25\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[14\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[23\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND3 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.DEC0.AND3/X
+ sky130_fd_sc_hd__and4b_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[8\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[26\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF BLOCK\[2\].RAM32.SLICE\[3\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XDo0MUX.M\[3\].DIODE_A2MUX\[30\] Do0MUX.M\[3\].MUX\[6\]/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_122_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_70_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_115_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[9\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_21_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[3\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_63_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_117_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_117_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_108_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_97_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_97_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_56_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[7\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_117_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.DIBUF\[0\].cell DIBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DIBUF\[0\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xtap_49_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_69_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_69_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_69_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[10\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[17\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/X
+ sky130_fd_sc_hd__and4_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[19\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_133_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_133_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_133_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xtap_46_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xtap_46_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_46_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF BLOCK\[3\].RAM32.SLICE\[2\].RAM8.DEC0.AND0/Y
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xfill_106_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_62_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_62_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_141_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell BLOCK\[3\].RAM32.TIE0\[2\].cell/LO
+ BLOCK\[3\].RAM32.FBUFENBUF0\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_34_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_34_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_34_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_34_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_140_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.Do0_REG.OUTREG_BYTE\[3\].DIODE\[7\] BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_133_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF BLOCK\[1\].RAM32.SLICE\[1\].RAM8.DEC0.AND5/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xfill_126_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[28\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[15\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[2\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[11\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[29\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[28\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[12\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell BLOCK\[3\].RAM32.WEBUF\[0\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[0\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[24\].cell/X BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[11\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[25\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_96_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[8\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_28_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_103_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_103_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_83_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_16_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[20\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.DIBUF\[18\].cell DIBUF\[18\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.DIBUF\[18\].cell/X
+ sky130_fd_sc_hd__clkbuf_16
Xtap_32_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
Xfill_71_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_120_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[3\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[6\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[21\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_128_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_128_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_113_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[30\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_61_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_128_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_106_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_54_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[4\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[31\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_47_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_105_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_57_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WEBUF\[2\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[16\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_57_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[25\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[5\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[14\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_73_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[26\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[15\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[0\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[27\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[9\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[10\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell BLOCK\[2\].RAM32.WEBUF\[1\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XDo0MUX.M\[3\].DIODE_A3MUX\[28\] Do0MUX.M\[3\].MUX\[4\]/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
Xfill_68_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.ABUF\[1\] BLOCK\[0\].RAM32.A0BUF\[1\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xfill_11_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_9_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[23\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[7\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_8_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[19\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[6\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_78_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/B BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/C
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/X
+ sky130_fd_sc_hd__and4_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF BLOCK\[0\].RAM32.SLICE\[1\].RAM8.DEC0.AND3/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[18\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_40_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[2\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[20\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[29\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[7\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_33_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_94_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_114_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_114_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_94_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[3\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[5\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[19\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[28\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_27_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/B BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND0/Y
+ sky130_fd_sc_hd__nor4b_2
XBLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell BLOCK\[0\].RAM32.TIE0\[1\].cell/LO
+ BLOCK\[0\].RAM32.FBUFENBUF0\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_130_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_130_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[2\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_43_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_43_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_43_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[16\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[25\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[0\].DIODE_A0MUX\[4\] Do0MUX.M\[0\].MUX\[4\]/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_111_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_104_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[8\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_110_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_68_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_103_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[23\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[11\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WEBUF\[1\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[20\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.ENBUF BLOCK\[2\].RAM32.DEC0.AND3/X VGND VGND
+ VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.DEC0.AND7/D sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell BLOCK\[1\].RAM32.WEBUF\[2\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WEBUF\[2\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[20\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[21\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[4\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[22\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[26\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[2\].DIODE\[3\] BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[16\].cell/X BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[5\].cell/X BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0 BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[13\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_66_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[23\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[11\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[28\].cell/Z sky130_fd_sc_hd__ebufn_2
Xfill_59_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[17\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[6\].cell/X BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_100_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[18\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[0\].FLOATBUF0\[7\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[0\].cell/X BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_100_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_95_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_88_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_109_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_109_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_89_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_89_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[1\].cell/X BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[0\].FLOATBUF0\[4\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WEBUF\[3\].cell/X VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[2\].FLOATBUF0\[21\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_125_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_125_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_125_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_38_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_38_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[0\].FLOATBUF0\[1\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[16\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_24_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_38_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[15\].cell/X BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_17_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_141_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_141_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[1\].RAM32.SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[27\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CLKINV BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
Xtap_54_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_54_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_54_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[0\].RAM32.Do0_REG.OUTREG_BYTE\[3\].DIODE\[5\] BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[29\].cell/Z
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y
+ sky130_fd_sc_hd__inv_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[14\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF BLOCK\[1\].RAM32.SLICE\[0\].RAM8.CLKBUF.cell/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XBLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0 BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[3\].FLOATBUF0\[31\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[23\].cell/X BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_70_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[10\].cell/X BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.DIODE_CLK BLOCK\[2\].RAM32.SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XWEBUF\[0\].cell WE0[0] VGND VGND VPWR VPWR WEBUF\[0\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell BLOCK\[0\].RAM32.WEBUF\[3\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WEBUF\[3\].cell/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0 BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[2\].FLOATBUF0\[22\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[11\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[20\].cell/X BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_139_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_139_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_139_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[7\].cell/X BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_139_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_139_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[10\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0 BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[2\].FLOATBUF0\[19\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0 BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[0\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[0\].RAM32.DIBUF\[19\].cell/X BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XDo0MUX.M\[1\].DIODE_A0MUX\[11\] Do0MUX.M\[1\].MUX\[3\]/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.DIODE_CLK BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK sky130_fd_sc_hd__dlclkp_1
XBLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.ABUF\[2\] BLOCK\[3\].RAM32.A0BUF\[2\].cell/X
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[1\].RAM8.DEC0.AND7/C sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0 BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[3\].FLOATBUF0\[30\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0 BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[1\].FLOATBUF0\[15\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.FBUFENBUF0\[3\].cell DEC0.AND3/X VGND VGND VPWR VPWR BLOCK\[3\].RAM32.FBUFENBUF0\[3\].cell/X
+ sky130_fd_sc_hd__clkbuf_2
XBLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WEBUF\[0\].cell/X VGND VGND VPWR VPWR BLOCK\[0\].RAM32.SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0 BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ BLOCK\[0\].RAM32.SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[0\].RAM32.BYTE\[0\].FLOATBUF0\[2\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF BLOCK\[2\].RAM32.SLICE\[1\].RAM8.DEC0.AND6/X
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XBLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE
+ BLOCK\[1\].RAM32.DIBUF\[16\].cell/X BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xfill_0_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_104_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CLKINV BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ sky130_fd_sc_hd__inv_1
XBLOCK\[3\].RAM32.Do0_REG.OUTREG_BYTE\[1\].Do_FF\[4\] BLOCK\[3\].RAM32.Do0_REG.Do_CLKBUF\[1\]/X
+ BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z VGND VGND VPWR VPWR Do0MUX.M\[1\].MUX\[4\]/A3
+ sky130_fd_sc_hd__dfxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0 BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[1\].FLOATBUF0\[12\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0 BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0/A
+ BLOCK\[1\].RAM32.SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[1\].RAM32.BYTE\[3\].FLOATBUF0\[27\].cell/Z sky130_fd_sc_hd__ebufn_2
Xtap_5_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[28\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0 BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0/A
+ BLOCK\[3\].RAM32.SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[3\].RAM32.BYTE\[1\].FLOATBUF0\[9\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0 BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0/A
+ BLOCK\[2\].RAM32.SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR
+ VPWR BLOCK\[2\].RAM32.BYTE\[3\].FLOATBUF0\[24\].cell/Z sky130_fd_sc_hd__ebufn_2
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[2\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE
+ BLOCK\[3\].RAM32.DIBUF\[11\].cell/X BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[3\].RAM32.SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
XBLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE
+ BLOCK\[2\].RAM32.DIBUF\[29\].cell/X BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR BLOCK\[2\].RAM32.SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0/A
+ sky130_fd_sc_hd__dlxtp_1
Xtap_10_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

