VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM256
  CLASS BLOCK ;
  FOREIGN RAM256 ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 700.000 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 12.960 500.000 13.560 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 27.920 500.000 28.520 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 42.880 500.000 43.480 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 57.840 500.000 58.440 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 72.800 500.000 73.400 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 87.760 500.000 88.360 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 102.720 500.000 103.320 ;
    END
  END A0[6]
  PIN A0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 117.680 500.000 118.280 ;
    END
  END A0[7]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 446.800 500.000 447.400 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 207.440 500.000 208.040 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 357.040 500.000 357.640 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 372.000 500.000 372.600 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 386.960 500.000 387.560 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 401.920 500.000 402.520 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 416.880 500.000 417.480 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 431.840 500.000 432.440 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 461.760 500.000 462.360 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 476.720 500.000 477.320 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 491.680 500.000 492.280 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 506.640 500.000 507.240 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 222.400 500.000 223.000 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 521.600 500.000 522.200 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 536.560 500.000 537.160 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 551.520 500.000 552.120 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 566.480 500.000 567.080 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 581.440 500.000 582.040 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 596.400 500.000 597.000 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 611.360 500.000 611.960 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 626.320 500.000 626.920 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 641.280 500.000 641.880 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 656.240 500.000 656.840 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 237.360 500.000 237.960 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 671.200 500.000 671.800 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 686.160 500.000 686.760 ;
    END
  END Di0[31]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 252.320 500.000 252.920 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 267.280 500.000 267.880 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 282.240 500.000 282.840 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 297.200 500.000 297.800 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 312.160 500.000 312.760 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 327.120 500.000 327.720 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 342.080 500.000 342.680 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 696.000 14.630 700.000 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 696.000 166.430 700.000 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 696.000 181.610 700.000 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 696.000 196.790 700.000 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 696.000 211.970 700.000 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.870 696.000 227.150 700.000 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 696.000 242.330 700.000 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 696.000 257.510 700.000 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 696.000 272.690 700.000 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 696.000 287.870 700.000 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 696.000 303.050 700.000 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 696.000 29.810 700.000 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 696.000 318.230 700.000 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.130 696.000 333.410 700.000 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.310 696.000 348.590 700.000 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 696.000 363.770 700.000 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.670 696.000 378.950 700.000 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.850 696.000 394.130 700.000 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 696.000 409.310 700.000 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.210 696.000 424.490 700.000 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 696.000 439.670 700.000 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.570 696.000 454.850 700.000 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 696.000 44.990 700.000 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.750 696.000 470.030 700.000 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 696.000 485.210 700.000 ;
    END
  END Do0[31]
  PIN Do0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 696.000 60.170 700.000 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 696.000 75.350 700.000 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 696.000 90.530 700.000 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 696.000 105.710 700.000 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 696.000 120.890 700.000 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 696.000 136.070 700.000 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 696.000 151.250 700.000 ;
    END
  END Do0[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 192.480 500.000 193.080 ;
    END
  END EN0
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -6.300 -0.020 -4.700 699.060 ;
    END
    PORT
      LAYER met5 ;
        RECT -6.300 -0.020 505.860 1.580 ;
    END
    PORT
      LAYER met5 ;
        RECT -6.300 697.460 505.860 699.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 504.260 -0.020 505.860 699.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 96.920 -0.020 98.520 699.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 250.520 -0.020 252.120 699.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.120 -0.020 405.720 699.060 ;
    END
    PORT
      LAYER met5 ;
        RECT -6.300 91.730 505.860 93.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -6.300 221.730 505.860 223.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -6.300 351.730 505.860 353.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -6.300 481.730 505.860 483.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -6.300 611.730 505.860 613.330 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -3.000 3.280 -1.400 695.760 ;
    END
    PORT
      LAYER met5 ;
        RECT -3.000 3.280 502.560 4.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -3.000 694.160 502.560 695.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 500.960 3.280 502.560 695.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 20.120 -0.020 21.720 699.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 173.720 -0.020 175.320 699.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 327.320 -0.020 328.920 699.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 480.920 -0.020 482.520 699.060 ;
    END
    PORT
      LAYER met5 ;
        RECT -6.300 26.730 505.860 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -6.300 156.730 505.860 158.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -6.300 286.730 505.860 288.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -6.300 416.730 505.860 418.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -6.300 546.730 505.860 548.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -6.300 676.730 505.860 678.330 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 132.640 500.000 133.240 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 147.600 500.000 148.200 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 162.560 500.000 163.160 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 177.520 500.000 178.120 ;
    END
  END WE0[3]
  OBS
      LAYER li1 ;
        RECT 4.600 10.795 494.960 688.245 ;
      LAYER met1 ;
        RECT 4.600 8.540 499.950 690.160 ;
      LAYER met2 ;
        RECT 5.150 695.720 14.070 696.730 ;
        RECT 14.910 695.720 29.250 696.730 ;
        RECT 30.090 695.720 44.430 696.730 ;
        RECT 45.270 695.720 59.610 696.730 ;
        RECT 60.450 695.720 74.790 696.730 ;
        RECT 75.630 695.720 89.970 696.730 ;
        RECT 90.810 695.720 105.150 696.730 ;
        RECT 105.990 695.720 120.330 696.730 ;
        RECT 121.170 695.720 135.510 696.730 ;
        RECT 136.350 695.720 150.690 696.730 ;
        RECT 151.530 695.720 165.870 696.730 ;
        RECT 166.710 695.720 181.050 696.730 ;
        RECT 181.890 695.720 196.230 696.730 ;
        RECT 197.070 695.720 211.410 696.730 ;
        RECT 212.250 695.720 226.590 696.730 ;
        RECT 227.430 695.720 241.770 696.730 ;
        RECT 242.610 695.720 256.950 696.730 ;
        RECT 257.790 695.720 272.130 696.730 ;
        RECT 272.970 695.720 287.310 696.730 ;
        RECT 288.150 695.720 302.490 696.730 ;
        RECT 303.330 695.720 317.670 696.730 ;
        RECT 318.510 695.720 332.850 696.730 ;
        RECT 333.690 695.720 348.030 696.730 ;
        RECT 348.870 695.720 363.210 696.730 ;
        RECT 364.050 695.720 378.390 696.730 ;
        RECT 379.230 695.720 393.570 696.730 ;
        RECT 394.410 695.720 408.750 696.730 ;
        RECT 409.590 695.720 423.930 696.730 ;
        RECT 424.770 695.720 439.110 696.730 ;
        RECT 439.950 695.720 454.290 696.730 ;
        RECT 455.130 695.720 469.470 696.730 ;
        RECT 470.310 695.720 484.650 696.730 ;
        RECT 485.490 695.720 499.920 696.730 ;
        RECT 5.150 8.510 499.920 695.720 ;
      LAYER met3 ;
        RECT 5.125 687.160 499.035 688.325 ;
        RECT 5.125 685.760 495.600 687.160 ;
        RECT 5.125 672.200 499.035 685.760 ;
        RECT 5.125 670.800 495.600 672.200 ;
        RECT 5.125 657.240 499.035 670.800 ;
        RECT 5.125 655.840 495.600 657.240 ;
        RECT 5.125 642.280 499.035 655.840 ;
        RECT 5.125 640.880 495.600 642.280 ;
        RECT 5.125 627.320 499.035 640.880 ;
        RECT 5.125 625.920 495.600 627.320 ;
        RECT 5.125 612.360 499.035 625.920 ;
        RECT 5.125 610.960 495.600 612.360 ;
        RECT 5.125 597.400 499.035 610.960 ;
        RECT 5.125 596.000 495.600 597.400 ;
        RECT 5.125 582.440 499.035 596.000 ;
        RECT 5.125 581.040 495.600 582.440 ;
        RECT 5.125 567.480 499.035 581.040 ;
        RECT 5.125 566.080 495.600 567.480 ;
        RECT 5.125 552.520 499.035 566.080 ;
        RECT 5.125 551.120 495.600 552.520 ;
        RECT 5.125 537.560 499.035 551.120 ;
        RECT 5.125 536.160 495.600 537.560 ;
        RECT 5.125 522.600 499.035 536.160 ;
        RECT 5.125 521.200 495.600 522.600 ;
        RECT 5.125 507.640 499.035 521.200 ;
        RECT 5.125 506.240 495.600 507.640 ;
        RECT 5.125 492.680 499.035 506.240 ;
        RECT 5.125 491.280 495.600 492.680 ;
        RECT 5.125 477.720 499.035 491.280 ;
        RECT 5.125 476.320 495.600 477.720 ;
        RECT 5.125 462.760 499.035 476.320 ;
        RECT 5.125 461.360 495.600 462.760 ;
        RECT 5.125 447.800 499.035 461.360 ;
        RECT 5.125 446.400 495.600 447.800 ;
        RECT 5.125 432.840 499.035 446.400 ;
        RECT 5.125 431.440 495.600 432.840 ;
        RECT 5.125 417.880 499.035 431.440 ;
        RECT 5.125 416.480 495.600 417.880 ;
        RECT 5.125 402.920 499.035 416.480 ;
        RECT 5.125 401.520 495.600 402.920 ;
        RECT 5.125 387.960 499.035 401.520 ;
        RECT 5.125 386.560 495.600 387.960 ;
        RECT 5.125 373.000 499.035 386.560 ;
        RECT 5.125 371.600 495.600 373.000 ;
        RECT 5.125 358.040 499.035 371.600 ;
        RECT 5.125 356.640 495.600 358.040 ;
        RECT 5.125 343.080 499.035 356.640 ;
        RECT 5.125 341.680 495.600 343.080 ;
        RECT 5.125 328.120 499.035 341.680 ;
        RECT 5.125 326.720 495.600 328.120 ;
        RECT 5.125 313.160 499.035 326.720 ;
        RECT 5.125 311.760 495.600 313.160 ;
        RECT 5.125 298.200 499.035 311.760 ;
        RECT 5.125 296.800 495.600 298.200 ;
        RECT 5.125 283.240 499.035 296.800 ;
        RECT 5.125 281.840 495.600 283.240 ;
        RECT 5.125 268.280 499.035 281.840 ;
        RECT 5.125 266.880 495.600 268.280 ;
        RECT 5.125 253.320 499.035 266.880 ;
        RECT 5.125 251.920 495.600 253.320 ;
        RECT 5.125 238.360 499.035 251.920 ;
        RECT 5.125 236.960 495.600 238.360 ;
        RECT 5.125 223.400 499.035 236.960 ;
        RECT 5.125 222.000 495.600 223.400 ;
        RECT 5.125 208.440 499.035 222.000 ;
        RECT 5.125 207.040 495.600 208.440 ;
        RECT 5.125 193.480 499.035 207.040 ;
        RECT 5.125 192.080 495.600 193.480 ;
        RECT 5.125 178.520 499.035 192.080 ;
        RECT 5.125 177.120 495.600 178.520 ;
        RECT 5.125 163.560 499.035 177.120 ;
        RECT 5.125 162.160 495.600 163.560 ;
        RECT 5.125 148.600 499.035 162.160 ;
        RECT 5.125 147.200 495.600 148.600 ;
        RECT 5.125 133.640 499.035 147.200 ;
        RECT 5.125 132.240 495.600 133.640 ;
        RECT 5.125 118.680 499.035 132.240 ;
        RECT 5.125 117.280 495.600 118.680 ;
        RECT 5.125 103.720 499.035 117.280 ;
        RECT 5.125 102.320 495.600 103.720 ;
        RECT 5.125 88.760 499.035 102.320 ;
        RECT 5.125 87.360 495.600 88.760 ;
        RECT 5.125 73.800 499.035 87.360 ;
        RECT 5.125 72.400 495.600 73.800 ;
        RECT 5.125 58.840 499.035 72.400 ;
        RECT 5.125 57.440 495.600 58.840 ;
        RECT 5.125 43.880 499.035 57.440 ;
        RECT 5.125 42.480 495.600 43.880 ;
        RECT 5.125 28.920 499.035 42.480 ;
        RECT 5.125 27.520 495.600 28.920 ;
        RECT 5.125 13.960 499.035 27.520 ;
        RECT 5.125 12.560 495.600 13.960 ;
        RECT 5.125 6.980 499.035 12.560 ;
      LAYER met4 ;
        RECT 6.735 6.975 19.720 681.865 ;
        RECT 22.120 6.975 96.520 681.865 ;
        RECT 98.920 6.975 173.320 681.865 ;
        RECT 175.720 6.975 250.120 681.865 ;
        RECT 252.520 6.975 326.920 681.865 ;
        RECT 329.320 6.975 403.720 681.865 ;
        RECT 406.120 6.975 480.520 681.865 ;
        RECT 482.920 6.975 489.145 681.865 ;
  END
END RAM256
END LIBRARY

